

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BXBb5I9xGRSs6sKck5vZDQXRkGljsGXwVGvqGMiKdsV6XfpENxhts93MXuSzN6nwMoqehO0wTaEx
k1DIj/UpXg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MnmM+Vq43VfUtOIhY9KEmYMnTOpr5zGRbR3yK+0dJHKXwwZLH8B0qYakf7wLIspjX3+ovqpgjWJs
eexIlQRGL1OO+SY8TKMpSpPoC27AE5XzJfVNJuTctUe4JhGeFQiByX+5cA58rG1UIyVu4V9mVip8
ZoHCg+AzWCi4RfYkPls=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eUhGO4Zv/WnFxc3Ba+3s+f/DLJpOX9sq8Be4gTyMUz382PTb/f4BzSbBQRui6DY3i5eftyc5tZ/r
9jkyaJJvfnT8O4dD86LmVGY8oX+idQzuT6rIw4oeMAjWU5UjY5v/yaTsmQhBcHwnQgC8DRkf42i0
XEqPpWe8H0ufxTjsCna4pW0lhD9kJOaO1+xySDotb2/KYHQnYNgk39dnpd8h1YlG59y1ow7rFcMy
UWmIcilGbYic3ZbL45pqq3Qc+KgOsRMiUkaRnpDoftYq6Hztbz42lF8rrwZUxldZ6UU735PTIlv7
l6EfQivncRW7xiJFPLrOQ8ajBNaclxJkf5APAg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TNh0egv4UJH4qDDvfs7rXQ/oEKQ1bFPgcWj3XkmFI7ALViHSkmG5TFA/n4HynV9CZVIa6lLn7sVz
2VsjFg4wMgfj/qaRkJPKAmoO8Zq84qzu762YbuzOfvXSTxIp4C5s/tA205oxU6Bij7tlu4cynXfZ
lFBFIXMYrDdJJSGr1PVtShFqGfeO/gOaN8Al/Y+raWaS/oDGb/ciu6GlxhyZoLR1gRfhmyCmS8GM
P68kAzVoPMQn4USscnGiG24w7VaFPNwxt5dQyTyiqFXrzy8YCO/QtdWk+3H4JxyUkdc0AwGH3qCS
tHz+2HVWZ9bzU6mSDu5okJQ6uKpzarA83QoPoA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FItfQ2y6HUxZgqq1+z0f6GElOMCJtzq6hAcJow3VuOey3t/fInfKfPHNfOH41ZYZwQ6bTMfh9UMm
TXbo3fDmT24V9QM5TX4F2RsHpHTe6NXTFElDX4CFzFTQ4nfp9vXo6X1FOz1QsSeQfNUheFN7XO8E
2UuJBJpMAKO3NlSK2A9X7FVt71yCUYCH5AItGCmtXYE8uLTQ8HfJqrPnTjU1th6jBb9Dh2jwhsnB
cM+Sq5N4MHCkgFOy7p437lRlySPo2Z5NRIBrOG/H6oD4T/8NBdsbQayFqVottK0Dh3VfTb1jwtAN
ZyTiNjnG4FJkzHGCyhcqEappQGlGNKwPGrmPOw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
s82pH+ra+n/uhrGCxzeh8pyCj7n05kyecs8hkcYvPeb2OjaTPUGyWjw6P4VgViM0Cp36AVrVKmZx
e2XRK8zinyrzSNWlmzmsfbhUdTgcreMAg1sD4GLrIibiVMk5z+2lk3OaXcx+3+h0+lEyIScEAUGm
JgpYhahET98Duw22gQU=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
f/e0qWgpwoVoit5qAqHiNIT3ektReghM3GOKqZv5m0PybAN0oNXP7+6xTCTySe5DzU06uDk/ZZ9z
SUxaA3ulymUsx/QeMKs53Et46+1ZEM+Mt5JN7uwe6ztqbgJCorX5ko1wXdg8eQ44KJx1WQqYtROE
Q2juHs2Oiu3TOo6Jnj+eAsirCCc95dhuajyl+16nZfO3YcBO3gOOOMP4AKok95MuILn71qEWpNwj
eukGjfxurCMjbVmULTQxLOJyMUyNxSIL56J5miPGfdxf3TdfDsU7oGDM07mla9EmyExnYwBAAPlT
26Ak2A4bYHWiEWl6jtGtmWCwshl7qyszHdXrsA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967904)
`protect data_block
mFpaA1Kpwp+jeZZdKkKltBZW1y7EcxaPxqrE4Jb9gseTOC6Wx+bbrXoCE33hq06cDtBUk14F50Hc
hUkD47rIHT0s7x6Pnc5frufXizOwLS64GE3Sy2sy1dwKCnlbYTIZOI2uazCPsV21w1WXd2ZoaL4g
Bk5AVEwHSKJPMVfuSIxRdH77M+102fZcahFQOIyoD3IbmmfNnhSeU/DkRrz6IZRhD8qvU9d4xGTd
la1V/TiQ1uCql70Y2SLP0X4cVf+MLQ1CmUN4utgbdzpdU0wIt6SRWpkxFfx5zIkQMUQn5o47W4gI
bOYsKUzdNwloW6gTX33OphADujMCdAm90C7X6Wdg9eAvFBmJoIf5TxKhxh1nJhh+qYkDOQe23W5B
pCEsrYJSYT4UuIZAZodPcWbQzM8FgzvfjvJx1cQ7IOrcRqHMBJFJ6NtRdpV3O6BbgwSmV3D1KldC
W/k3UPNJHUWXymiiQtoXNREk9kKvdG/agtymdlOv43yNU0hv1T6cr640YdxnVj5g2cQL+qZrYqRh
nKjS29REdZ4hMSfTwjKxePstNbb/tjT8bKCpi8CwQepfwkL4RYCYOgOvkvppRkNdt/ugfb+4XSeN
WIOpuFv+gD2wYuoD0r3TJibJyUWMG2NRi+XUgcO5WnaB8h+QfTKd3JsWWse7MeePaw7dEtE5esvP
z0+jhb99r+DQkS84/AZJRi83VRkMMx8c7DkYRoug2P68B2Sml/AyztOtQbOrWFYbZX4jgm27C1k4
TEKfdgx5MyyvBvP0Ww+gsFMjGizVZCCbppQSO060wrlk20p/UQI8/TGMC6cwLkrhhbv6RKMxMtq7
lQ1tu0uzbx+OvvU9ir1KSwPgd3lp/kNGK2ou602g8CExYX4S90lbX7VLMWqNs41tpL5DXUsbumhn
HTLb8UipokUQSGTiYkl+PqVIDVIWiQ/mFKsLYzlxq2lGbhmxJP4PA2tiYQ64U2bTqmHPkSjRj6mV
x2vGarSA24lCCf2iA0VJmlIiEYvcQ7feMEOMGxfwJZIjfUwm+ZVTY8+oRnngxZPHDraT2lU71woo
eWxotOygWiIQTohVp78n7k/LGkEi7oNvBZkLGbrR1J28nM2Md7m8OzgzHzIAWaeR2/QSWk7J9ISD
oNs4oLbvNuB0FPDj7lYRhyXi3SeCHTAUPlq5Hi/e+R/uLoy3EiuA5MUvG3sWJxw6mNRKf37ulsW0
VaviGDgq9UjrKMXSG4kN+ZaMT+XReRGuDJdvoC6bMoaRadPNqXep5gwwRChpXeZuauot9iaSJUc7
h0IONF469oaHtfht6HkNottN7gYzrYVRBeSSLw4LtyXkWaN7rWAQ44h/ZPCSBooe4UL/hQVgVUxP
19mkxuR+OCI+LEHpCixfVDPmuwOX/O6xkrUiBo3NN6SL+HAFpjNFQs6amWCIt1HjLnn3GBTTLSwg
wy9Zqr3k6n2IoanS3+taYCa0uH/hU89/DL79WGoYpp9JUmOEh1nk6M6sZ1cBJ069uoBBHmLHI9Ie
g5x9/Thi4gOkxTe9HhbneD/n1YqKcFMy+Q7ERjqCb88bBytm+lCfZdsX0HSgP8cjr2cqAiQPqndx
HJGPga7G3+YEFsn59UWv7JrLRI+MWJJ1GCLCkJn7D0U8c8VyCRgEEl9AdaZJn8tqcqE2RpzQEkMB
RhWouPgM/IljCeN38EXrXP95vW81eE02T6CZmuiBUyVB0kHB1NpX5Vs7LtS8Xf+HC7ublwNEPnU0
DyR7kOHYdpM8cbjNWhd6vQhe4uNhpfkPf+U2NNP0LOOWedY+EZGHfAlpmjyxZnstiiVrrnzIYaSd
K5c6PUTslHxM8DzolK0Hv7afVLr2rr/EbDIWJHIvXZ+MIHypa4AFadkSVEkRnM5mnMIUaq0HqDpr
FZLwlbUeLjSmi8AGI73TkK3NgmMQnI+cTVsu2Jqgz1uxmzdDyI9U7UuhDNwj9QD8hHgZJeizeX6I
/7TAsX/MtdXlHv4IapXORR5bHTWA/wAgp6E57hxd16dWxWiH9aGurxjuc7yr3VMjBNigFhNGZsYd
b24Auhaw4QVU49SVD+Rsp2FrLX0O7xaTgkazM6LbrqzgCt7+kC9vWDwdHeG5LyhVB0x/eg6SwIzz
otyyAnL2ScygiZQD6j9l5RZFh4Rk4cjEX6wr59e1LDa3EQ0382DPm0wV4xVESNPyMNE6s8jIp0Xx
eBo3VZDoaqtGQh3ySsOGYjjpRsZUTco0YBQCXWO2KUDDEDokwUe51rb/5YRdcereKI9x3jl8pWXh
3D+Iq/2in9YYPnaMYCqEXMOst0ZoDoWUSd0M6yEiYWlD3lO/Cbk3Oe3rKxrfxTHBe2IFPH8SlbYW
2o1kQu8H8PRVNpKz7HjSMR7aPW/bbfIZtq+4u9hCmVyfEzsNNZn50FYMdYW5PuL3aMvWQLiaJjfB
yUGDB+wc2XJbNyse97A4D8+XwwZIjEaCxlFA348dnWpwYXiwxGr+tmKy+MotbkWu4kucLLsjNS3o
s0W6SBMEsf+7yfuvMN/orf0G5oP1bZEEu1chmcLD1NeOt92HXH/82Owr4rXRtzBFislR9ewgEa58
9iEZUwRDQclO+f20rHF6sx9Fbena75JWvAMrH2EBNfG/njJaM3BXgHahk6EoHTGz1h5TqIx1DK76
v1q302fU9x1D8Cqmb258qFO0QC/KTnYYtxdJWbymP21bavelvKyjM5Xw5WIkeHu3Lz74WPJz4jyr
wDkrfneVlZXNK1EXJFK5Lrx8atxIPoBZvI76XoXl0TC1iiQeWB0KVbsNOAASTouKGPIw27LVGQFB
5iIry1RCPZ+z3xv/Z2Ih8sYV/hkkyhTKmkjBH29uOwzWZrMzUG6IS5BVbRk27iY+sru0rF4jjqPN
Lqe+kSBLwdm+MM8O4Y1gdu2nU6/t7d7TC/e2qilqqgLCJQvAbrKy3XMfZZR4IeM8a57wj8zo/hSZ
GERRANLFbj0CmgAu6plGZU19GR1orcJLzYNY9spE5iZ/OLviJpXpqh3lCBW3pBGF2sIA0rsl3cNQ
jS9zQMwrWR+qGJeLX7xo9GU5QOfjurB6DcTN+3ClyJ36UtmaDjRoOsvNABlF/e2ygNz23Ow8u19Y
vlhaR2Nzs4Mn8rQHyY7YX1pt7s74hJHMoFZORIpOL18g2+Kh5jRPeUX97lw5NfyK58MFtWK/0/Gx
IhtAhIp1SnchoYU4SXj2fZHKhGq6qS/5FUcz5U3LSVZtOtfqVKtXatUGbxG1V2XygdDqWxqVsMWs
aFP5o5xEU2LyVnFvZMWksypbR/Xo0UFS8JwtJOH89N3Q0mVHv1/cNjulUyRg++SCUM3XNVLqTfVq
nfAFN8N4Dk5U4gR/HyE1Cd1PkDriL6Kj/Nb30i9+YIPdVE7zgWQcTvmNOguuCqFz1OJ+ZHy+z2Yd
RMMUNKvxTfrRNdKlfDvfg56QjTO8fudL6+5KhPA6dZ4UtZDubw8ueAmiVp+pEMK1pZCdZxUh+4Bz
ytVP1uABl2l05OxRIcVmjZocO36qTDmEaHz9KPVUhL1bnxUQv77wNOss9RlERBYtwRORJahkVNXp
iEC870PHnoRbyZvFiePZUmIBP+ua8m9sawqIEAi/HGEoiC5FFPx0kuMCu8XLSfao7cWLMPpjPxi5
yDoavxtPOGLFYF19dlsHcBPfa4rmwnsHS1786RbRjTFmH4Im+520NMEs38hZxTI8LqWpfqtAQYRv
PKnE39mf9V9zhGOWYUWr9Kf5k4Pe8qXtIBcC41hhRhB5NpjEWMiQAewFwEhm6bWD0uF+a6nMLzv4
BO6E2X+o/5H4Mk/pru7Mskqbqf7Z9l7kvB82abeG5lfZLVWlKwHIX7EKhKD3VwPQeR2RePpMMX5X
HRJ8KZerLvLXeDZDXABzdA72r3acByZZZnDBxxbyAE5HmR6lacIf2gYupSZ3nUQ/layPAnfVKW9i
ZBtlvK1OIotNH77wWhxFiYQmW82vzQpJ7dIl6xkNlJEtURjp5SMMny99FpV2LHXKUEYXDmNq/EmZ
VrzQmYS7FHQHUj9rKXUfr9jVyTaZYRKYlG4ojicJgVdojP8NTpmgX+OPG5VYHFWS1u0tiaJx8lKf
lqejOftHMtRokfh7Ay17+OEu7tbCci4aaS4tFhJXsbrD1q3nazplWCQre52qynplt9mYG26hS6nu
QmDV6pnSWxYSwe0WSBae6Y9jxideRGzcyQgXQKEpRRIHUA6NAU0n5RHlKx4NyAyxT/zoUeP9GsEN
cbhJrQeMHw9jpVnRtJrtk07F02Jx1jABsB45iN6Qh+KPTpVAomfTNRj+Es63YgYVvaiV/1ZX/fHB
FDyGpVpeVVeIJjmnRSv6BQZVQRomGgi0O2CiGuQIwdRagStwX2D7RdBx6XjpdS/PdQLSOn9zLEqi
1GcpSgOyhDygYYVotll5jJJS1yGdka9bwTVTantDziU5Tu0uwWikiS1b1JE1XjhlZQOJMhzdVw4D
5g7Fz1su6iOwN6O7bfc94IXqLV6ZYFhYUHUBJ2cBkecqOjzwuzbjR1O1sTCawCF0DqNYvHwyiL/7
SloAEij28QnQTfDTkP7ZK48BFgbFR9G1sytxjxk5qBgtbfmF4ked5FoaAcFRL2KTO/KfcHNQGWSn
qA4TCCDA2j+MhxSVkNknUg0wrKOO1hQepq6TA5OXMZYB1SJxnmMFd/fBTDfmTWVFF/5K8rUwDg9X
GvjmDJnu4IavobBUgMGmT33fpS6F6E5osC3It1fz5QmaoBmfyvF5KbDBnzck2fwIte/qiwhS2JLU
q5khUyFmK9ANLENXCztHGtMIDn0rfVUq4cnpxSQ8Brusj8Q5CS954DO/t3Ql3DJg01RNLyCqTSG+
qvnaHm2LzcZfCmHCtOatDomVmxlhHFTjv2fq3T2Xl5+LpISFjj4dduQlkx4VG1W0ClSWrxS/B/R1
3O3EZFFyHROD7Bzz+8Y5o24GqCfAQY+sk5kQEOjjJ7/08sOD716BNYauZcR6bygMgTJOatQdiPQU
x6BkOf1aXdyeWhHoEeXRlRLf3fdjTx8yAiQToaaW85VfiN24LUV8JJ25o1CNXrONNKCxXI3FKKtz
gyg/oPGfwMjURZR00lkldSc7OfywRdyHOy2zfulIji9+Ume6qRvtdbFOshrdd02GkWTjgsr1Kktc
ZakShyo1B214PoMsXcJgLVITmLkuRFWB+LlxW+Nslp/yZpmoLfhxzywDoN7KhTlZIPMyrLwPuqM4
GpqXbL7jEqW1J+37agG5q9ytKIWB79DARazExk3MMC0MUOdbZzQASBmihJ8aAYzjB21wNQQ0/fj+
rKVYv1teL4/gkbRQ4r2UszYEYL/hIbzzczfNzS/TYR4P5DlVlBUx1Y/I3t6gRGyKF8y1zm9TnSiV
gY2OH4CEsOmo9OCQ7apxcekn5tjoxQux/YdwnX6aeUIZQGf/vTzt8G/HVATRzNT2dsgxDdVtqBni
jytzHLmdQzto6XgdzgQoeGUVR0sWiFmpbAgBCwRavbLFExypLssD3tRBg8vkqANRGzS/lh+lcG7i
PaRWz2UmtcWHPvUmB+lG585/yGhK3dO3ciXkhZu+v4EVq0yoKwXzNeD6+eX5Swmc847b7QoyRc8p
mDcm2ehd5nPxbvt+vW1gLYxTriIQGPoIeaSLLWuvOztGWaItJuTKBYjLhuTx2B0+Lx0yp7mpsi3I
9Aj4KIaklVLuTUdHO19dsnSYHc0HDFxcoUCdVvNf1YHxhsvhwflI8td+dc2gI36apxyzArTvARCV
DkyAHBOzXcpvmMg2U7GBu8Ebq84RdYJFe6bJnCVfIFg6eKr+YJMTFm5U7sSBBkH8RKKHzpeZQGr5
af1n90WH7znIJTurMy2BWZacHbhlI4Jic0XRcwN+g425K7EG3okgJKAgJagdL4ADdgORFrecSmab
WzZ3xjRG6/1U2JAahqi58XjSvr592xki9JMZ3hME2HZ92r5RqmI1pJpC7GIDHemuLB9wgmcwVhcC
A8CLmwbYvy1niVtd9djuj7BtWd7PQp400TeQwQPMp5ivdnIzBwF6uet0W7rZZb2hdgVqHYsskJv1
7Oz7D9hnRPS3xuwL0THwouDmnwROm2R6QXaoYjjXO09rrgSXhjr32BKT5iMV7SRWet5xIQr5FJv4
pv0LztJ8SxbVSu9zD032dBKlxJ4XnogyZ1kcxhYocmj6GRH1vUPh/a+nXUhw43jlmP2GZBdHa90E
IdmJ880ZD+AvAen0lEOd/sKI7gh14IpxTmZNDhSEvD/cZMK5Ug8lvUSH1AjWMCWv6q7Yz8XI/Ygv
DM7JVqzpx8RdmW2ScCFuLJd/BDTu8/W8JoWV2Epev389/e+VJOF9Sm1NHbWAtt2gZTynxnotVrkq
OURFMVew1IFsyDp7+WmIDF7IFi2EZP2rZMejglyOaZPu2hIAk+AFC9O84hm1GsuI3rqbCct5EgCc
R31rwNiit7ka1td58ZndL5k+TkBR/0eLSwSxp5jExVHA8OiHxC08vnl/ndNVuGkuB17vWok0G4Ep
HvNUfiDl1iA8NBOJ3mlrjXI2O1h96Yiw/lYmixyZeFFP6d4FclZEwR/ykU52+tJ6W91s+0RQ/2Zy
gLJ/1kWEuIJXy9U73ZauLGOA6QVwI8n2NPIje0tG2V/6qAStVSDbN5lJdtZoZaE/3amv/k2Ocx7Y
WaRgC7g4NXvqLafFSgVYn/3ejJytepGGYpx+guK/kzgQxRA307AcICIQqfKIhrDUwjrnYP/J6wDG
qKYupwMRCPNCoDTJUv+6Wh3A2o3C0nY3W/+TcCnl3ynM01u5q0ZuU8f9kSDOufeMinwzHxcu/41n
JMIRSI+saWAKX5mH/qBk+VjhlBJO+CDF1mLWez5S4IBgB+OP4hzQrMhSeqpjGozVTRWqkUmoJJLE
Edwwl88SxFE5irmmj8NE+o4rHQBPpO8U5Ce1rfzV1BFUfF1Zatpmie693HKjfhlcDN95SQMbVcLS
dN7vmnZI0A66HGyjgjOQ9n8c/Zd/XOAFndFDUtfavdozQYW9htqWVa8dvqipVtBwJZmoXu5qBSwk
yJ1paC7GzLV5Xj981T5pResZ0EEP9/5N0Pp4j1idNsM9hw26CWSz64Pryn37dKczgxrWFJf8kyyW
/s9HcTpDuMKbRqS0II87ygf1JX2lNQpBo4fUBcWi3Q3ORclv2VaQoVgP41hQfZa0J0+B+IU2MWu+
XYRzwT+ltB7/+wi7LYU+Fqig0gk3OPj+4s0s1AdvYA5cZKh1iE23XH+2lS4JM1iN/7XOwVJsMTD/
ERZo9Pm7JLeETETpQJMXhqt7hXnc1zd7LG977OUg9voI5ukEeid/K+Yy+btVStToDNxetXhOy4Mn
s4mKHhG4uOtWURTZ57UYPG1GH1YorqeS9ZFVZq44HsT1+9eysus5UvGvfShoSDTGjVlnkwkZRmch
ZvAbiD/XS3pvTHTaSUWz+mztWkwQQWl8z28lwYKwV3Pv1/xR6F+EAmf6Ta9KrAwhnTHEkqkb8Lux
0ow9F8FUiv047qa9+O0iwN9tQ4/LPRFSgKLi2uzlF3XQz7iAr7naMe6z3MmIek9N8qKro1bB3OTI
XYdKyj1D0OZSvx/zQeilGg0T2Lz7hEyczSbouWCnBLYoRtdIaoXXg+7R0J7P3v7Zb+2wvMUf0kdw
0z15m73UMv6FqdK7A8opjD5UFEoZqS2kMNisONNhysQPd6pD1925xSYrH5mIhRp7PTCvYDoGrsNE
fVaisI1+9EwPSm+YJQdXimrQmjFpHO89uf/aPbkKRBC4UiNB14UG+EjG0vl12nhAuZKWP0mhC7n5
aDEFY8WaFjEHZ+TcDUuph1v2a7F3sg3j3M7IIOAZlcRTbT6dM1XJBDFLJpdAZXcWl/MUCpNcmlxs
IC/6L6bZiYVDgB0xHiKEWtLaJOiRBoy7VR8CV3Xd6Z+/dGlIisrpf4CDv/8mKJEbMCNg/CjZX3lE
HRW3WfYP+GLAKvGW5zi/MnR+FBB7KYrWi+3QLHYXh9xgxjd6R6JCPGWqjF1ocVecsLvazFnHgbck
LWKI4CtYXxcoynPNrlw3kd6ddOveL/yuPn+1LhBtZEZoL+uSojZQXP2LlnF7hmH+hGF9QHKbuH0O
EaGIYex6c29JMg8XkvNjszGtlWVMmuFKczgvWqi6o53zzjQORkZw1X3SFS3i4o9JFUfsUwQRRkwY
b6pgf8n107TduOAHtoHZ+ifOv1dShies58QpsKd1rJTvbewsJbs/yaWDDSRN78Cw1lI8ATgXbDTF
ydP1/o6tEKX7+9PzXgD+l7+pmzBc0Pi3pRn//SDviUON31hHK7nz9yokpNN55Ve2fFfTkipTItg/
43ocMYcydusdSkU+286KCvtGzVO3Xh7XQb/tcqiQC6VYuyC9dDLuoTj/W2yWA38F45rdYbyBoyni
kbiDSBePit3URnULAu+8JIsfXMaJRkb5WicVacRFwnOa/cJCiMaD55Vejn2+p7dH+l4qttao5Ljp
OIiONh8ASQcvk2ATNGL2ZKyGPHeytYhUrw5mgWwcOkblO1J7YvSq+hpb18W7ybFC7kwheOqyHXKj
3iwFUp+xO8tVpBdbQOEwg6HrN9aPkCnjIQH6uT7DsagLuKlMStDPK6G/+GQIAbq3mWzdRH/mnftJ
4SKs15pI2lvrSrXC37MAm/c9seUXaNVT56qfz9d34jOdb0MgyOlwxInqZMCMqVhO78B7qFAzzARb
CHTondC2rTHHH1hgyOfSpA1gWBk7TkgiLDmVHCD+2tw/J5bYTqN0/I26PojEAiz8uIGmViqh1rFd
iRUMrx69Ygn8Rz+GQTkqKVZm4FsBhethNp0Ms8GDoUUHBwX8HyAVBCt0Bsas0Gz7OKLrYvXLCeHI
/ClDZccVURnRh7YpSTa/zoyBBu6fJeqJ57lRKTgLh4mXN4NdPHipyn0DT+i3IxPORJRzmjudhyO4
rOJgToV3jopsjkOshph/BXNNt8aJhkPv2eDv7biemcGIZUUOUYVRGiKX6pkNxJoyggMp5Zt5+WWn
GlUZWlgKothMahJkPiP856JGSOSnY4K8irVRz5uCw270CxgQndyoWB2jbTzXtLh1aIc6WodYFlo5
SfuimjT6s+3xsi1RjAAED1XUGATv/n/EvpQZzLV7nPbka423/vYMLiLO/q8khwWxQ923qdxAF6Uo
JTwBW3iII93+H6QQq9Zo7noVMEHv2LiUDiNbKtIP0F3Uun3GpaWEkzA8oCBaby9tkWOCIQ181uBq
CC0RqHYv6h3s92puf10ycr77Y3WAw4KWzZHo3yJWYaQDtIJ7SId572JWifnQmpTP8wW+I3noMoZJ
VjMuVbfNtSf1qGxdZjorLgkPxAvu1KRPMMq0mD1Sq0RefN5Mz2QQsa+kcHV0+E+XV2fyrJb+po4y
GSa9yGNZhofVjwLWY9uBdcfu911RKhdtmTxS6qOs6v1eLYIO1pKFXB5jAU10AnVpVAKasahW/j4w
u92KsUz/FKljng74FnyVTLrGyUN824otNgqOC0cZaRNjObTHtwS39e7gUsjz1ggc6JSXX8NfUzgS
sga0u1LRAgu0fzq+lKoiT3b7d9ar68q1UBIanNCSlbJ9hADU/MK6F47gf/7nt2MwakLVt7CqvF5Z
u6sFHPCE1nm0mNj6CNS+77Y49auxrvkFSp+er8MtklQ7QwWcZlvnqw709OQtuwoUvtZZbBZpq7lx
N3QPpfpG+YR7+2DbAg9mLKdWrT9oG49FL3Djd/g3nBAWyAyHNBR5lBFVhmSZHtQi/F7FJk8wUg/v
6pWVitlY4Z9/4EXhHKHPzRSwnggIP6iTbGpEjOeh78pMyZW7FTU/FfDpkYv8rS8wkGx9RkErw15W
9ONdZj0RusOY/Qi9d9J18a/d0Wjj/6ieaTwwmKXFI49YnPe/LZyKeOdzere6d1NNMP6Jl9Q99ZeB
chpH+K7/tTaJZDIwsWvEsmbxBnDfFNHA0f6NBnAwqRFb1bWx5DGV7N0Vm8nAkpt8BM4iFMCMTCH6
7/8PulLtI6JqEnvmy7HSyMcFgYPscxl8LUNfLk67QlNR450mLjUd8W1oI0QwCD6U06XhJCRh5G+6
hG0zk0I+7u9DCjaEn60vExmDqa8P0JiMvEuHgbDY5GYcgjGU9iw/hycf3/NoXbDDMMLiUFYqHeAy
BZYB9yekHPXKO5r4ylDg6BIYGYHv8+N2FYP46FzODghIqqhbsrTR9gOKoCYGYEr68HCU0VoFJ5gc
QK38XGdLNNwv2zleWZdqlHb1ZWmIAwHv9NGBoSi3WU5fO88PVQqXC0RnL3OwYJHXrlVT+pbn55cR
Vpsk5QD0TbexA39vfs26Hh2PPGlyRA2hletDSH9rf9oxVYriBNHfIb2J1ZrQ0pZ55YwF38t3G0nj
ld+v4thYZ7PETi53jZDY5+kG19b+5rljqqdgQ8gO4iXpE+dlCvX71idkC7TPFU5Frwmjyis46mfe
1N9/7M9CPKCNrSoJImATTBS6DXC0rFhcDelEdwXKnEmfu4EqerKBOTnm0TzV6v/8J1XRDgHzmIdU
5yjrqgGViI44tMWAMYbIQFD1A+k7EYLZ1wVh/xRscYRaxyE9/yuA3lQPtH8h4Db8Bfjhm5fsKew9
irhbkXetxfv0K8xgwoVH1EXMod8Q1VtajNnJxMC4hkph4TQjbcqrBLT3fIRxZ758SXS5brjnJPTO
O1OG4vmbp03Jx/HHO8jwriDUVk9HxrfrUYhFVM7s5Cld9cr8hTpoScvPSKjAZ29DALA8CZG58DJB
3+XBygRbNZ0k63SNAjGPh956KavumMa89hbfhPMNxok4uNXIb7AgA98rpRTrCxBo/1DW9iUIRLiw
2XHcOrb0+S+msEJJbTw8qaxYGyW2AXtrpDpgHYs/3FvxRQnI1BKpMqP1KLa+DdUKmYyNgC0uNCNZ
cq+Clhr5ORc5nciul11dMo+QQxUMHhR3CT3ThYujMaBXyNBgsviNaJ4lb09OjytF+SzSri68KGiu
Cn1K1mTvTysOstYmb3pgyNUJfu/YMkuR75x4sv/oKRii5axiFQfiCkcYwxbPF/dW4lPEQZvVLobj
PMXvaO/VaKe3IW0Ovxi24sfQzDJQ/H5AtouI54Sh91FOLwG7I6U2OIphe++9lQRZeAgOu9mvwZAE
OZRTde48LlY+6Sw9x8dQJMIlAR3YCsT2n3nNAd990RAl1OVkTSUuB3hIcipwWBqSGrmicI9srmVf
1cCA8RQ+wcif3Kg9fw8J20Crc22eeobGbyY3KAaTqrHD6k864Afxy/zSjG72TySKMh6Lt1vJggFH
4Co72XO/isGUdruDpAfu1XTnXXEFkRyAhyRTKx35tj4nTGY/VaRVaxHDS4l50zQ7QGUfdIvAim/4
T7985P3dkqmWVfSgCUjbtCymdHBDhPnGWqeLe5X/Yzx8vF4ZxuenbG9C1hkSDiUI8ztHQ1yQdJQY
75CsdliL6OfdsgXf/8maygKEI8uROa/LoBzTRFJZlOL+q4u33BHQJ1HCUYwDBtHd1HQ3IOO0A3qT
0jOk580t07QA28+/D21q//UFSxJexxNHhe3Juk/kBYTVhaY0qnIfYg+fRMuAAdsvXlqoaWQpbk6F
kkqmNdj6Ns81z2OmI6/6Bs33L4J3q5sezF7GpnyyuEoLogc8/Z6t4sUvI+dbpribCHAnwy7s76MJ
N2T1ZQbgkn7+XN+FbpKE+f5a2ksbQIx71PVC3iEoPDWgS469Nl6eORAO1HvshbnIXnA7eSFkwngy
t+UzMCSTTUIIfjGQVJ1fZVIAwiUQR0QaA4+Hm2nxq+6lFkjq9m5evvtA5wGyr4sT8Aiyxaog2d9C
o0tSK+5filAfbkdGjySaSAwss7MdIgVLjdtPyceGk4zVpmBCVxNSQ21cie65Kj4MAqxgjSp99a0Y
d3hSN6QoOQ3K/Ihka7MPdUFt++VHuMEriXNXflSvz9cpReUaN6GvYiFHAeaKLXCUYLyKRfBm/R/5
Aji24bwkRs59j3q9Bi1G3b7ILu5QgNXHzAQySMpY3lvszfKjNBjsUjkHHvjXqWcg6cQ++qPAy02L
6uJQ79G6zDfjnZnX5ntuZaPe5XfUep7RVqMDMGUCbgNhDHyCXNtIkomFB1NBq0uadFf7faaDXpWJ
OEZVwqzYjPopjQ053EjyZ9EzJle7PbmyriS5vJfJJ9kk3VvN8e+PEAn0n3mGsdmv2otADnAlDEUY
/2WrGe/Y12NkAEU1ndtzkIW/0fzIHtVeUKcYR2/8pFiQ6XehA/+PKypPyKTlo1WltilRn8oSCcR6
4nFOVKH894CLs48EfTcE5hngDQplScrM88GVY6hSwVhsNk/0mFoJiTZRyKeuQpzEZFulDRljPdvT
fVe6gTf0/G8vGG4fNAEwhA6y6f1UhRznKZF7cIYvtf0vYWYrn4teaVhdYTBVOutvTZb29/Kunihs
YGqZjNfHEiisY6h4mo0nUovFYbKUVghIWfn7m47NBcrfuIByuhywke5sjoNDDAO55g2ktudLchP9
UlOlspHe1g7VRhchUk/0YL4Z1lnSERE2TaWGSittC31IFGxiYB7u74YLSpZx/gRYwH/uFgXhEWKt
6kZaVa0jwtj6CX+qi6W6yCaQlkHB2WP2gNK/Zz/AJt/qnUDz1MzCAaUOOVegAEExeXoZsRsJwUkK
vBAvHap0bOFrJC4sQrsGkgEPfzqIvcBDbaY+RKpeegrcaDwZ/4SVTBIdKL0GzxDd1XZMXYv/nw46
tGMB4twf7P/RK6Cm5XmVzZz5YgZW/5c689PaalDawscYwgbG1Cctut6gP1t5jbR8n/Tk6X83pjyW
SVJDyTRBiTU/Nns+08fWX3FAKf9US+6wwkx4QxmnCexQMNlsp/CC/kGZ0XmevUg78CRwVxHiyNA6
wFKgRt3glpN0XXtM1+5QRk3nKR+QAWgAspLiIBDSr3yICBtZA5U+z1VaqAK7STVc54+f7IBEq7Oc
svUucg0jWLsQzVCJv6Bu6pcPT048SaKbfd2M9kZQZcE529IbnubRoRTn3/eWRFA+pijF3mzOn0G4
ZApBSO+/0F1CoK3IlId1JeQMm6b2WYklbNXLGmjT+Ci9QbGSwJAvxw4pzwJgz221OMWofBN8cxKO
6xZdWFusRcwNelQAbdg9AVVf23oxb0+WPvrNPfWnevmSZAe32b51HISN6FpYl82/u2KksOM2L7x0
AW+2Ltcs3hVga8EJjheqQcqsyCB8YG0q5wZKa/qW4RhEU5k5N6Ty32RWsIXMBCBvJb5of7k4O0O8
ReBdtZWCieauGKsk/jpPgaxvj8VqslFsgb66LxxXU8qo1ZoUSh+DieMy6D9WzkFhcdE4/MCEM1+q
12zzGNJy1ehum/TR2EUC30DgUAsIQBJzLO5N+ghB/g2Sz50d30lbgc42eiJ46cXbcyGPt8hUQ/c1
qkMDuinA3/Go1J+uhKCY7JAvjeYy0Ecnks3aBkGi9xXzDg85WxYCzXxIO45/ASbseNb/jTN5XhtV
biLEhQKFQnS10HGhozPv1Z/NeMf9MyID5VKaJ/40/ctu+SguODoQveTSytnIQoGeoxnCkO79o4e9
48gBN/oWzw9nfLrCTyuS9QjhoM8blGGP1BwhTI9kMz9tVZ9k/5F/i3dzwHyk0tT09rNm5LCr10mP
JRIZyVrtrFZtaz5xJ5l1iSwtQamDGiezTmy5Lm3RC3S1KwlN4SoFgPgEbxWQrdQPUGxoJD9rqBfa
Cb2bvsUZ+FBQNp4jvivJx13PuKzMg9uKwkn3pzz0mmyKVWwETZUcmsiuns9iw5B/sH3vxVf4Gn2l
ND35AzP534bK9dw/6tS+znEQGIp1Qg6mHMd1uWdZIoJ5eIaH1PVC5Ld9S4DU5PovBBRtk4AmX4w5
Ln3IAQkC5ZjKucRmG8rrb05xOmFtzGgZ5/a0kW2dT34VQbTmVO17HkTW3/bYONQRyypYlHFJQO08
aTAlGsT2JANK5ezqi1GGYNC2Wd8ge5Wg/Snd5ZFOQ+yI+qV1aJYY+ZPtvXrA452OMlilMr2acRVu
0YyEEpeFrDLOpYvDEngpfnaCXM0gqC+MYPB9gm+qeYuk6KwCPFP3fLGqkd28HLonFbt+/aMmT4z7
87kFZBywNI7TBUk0zL6tXAG4DItlk62Mnd0SosmCl2EBJnR4Gou0lrr1vth5zbC5a76C0PqWgq4a
R4QFzJkYSBQKLz7eP7dZ5jX9MALSX8DRrIcY3XKq0cKMKHqs7yqidKPsa5FjdjJBOl+fVAeqU1Ft
VrnmKQAQfuH4Y+gXnQyhn6sKvtl3Z1Mg7+SFtcfLcyCR568Q+F9z691Ccw+Arwxx7fJZm7ZLl8Ah
s6t58hCNYCwYjWglR9+2NLMs01PIpcbRR+B3rE4zCVij0MarZExY/kyZbVAljViWlpozO2Zdzcuf
BnPWqvbnRIsELmGyuCxmGB2FOLVZcTpo6vJ0S+IXjjeHDszr8Q8pKbkJrye9hupCnNMA77d9BvMT
xeudD//HzSEOSJtkjlCrV3WhR4i8Pu2bgrUc2clZdOhSXlcVlCvkcBAeGu4sL1zbM5RAyQtZPVJ4
GQLXV1NGVCdpvM4LAe+5bc599fSqxDtWBQpbXioQ+JFAil5L9phmX+S4S20aWlGKt1D/MNXDsEcP
WB8DoILJOpNdakU6mkLPnVKPvBPdJFgHYXm+2n4c69H/+sOgrlJG0aBwcZUME6ZXRSHPDUjTvjuC
MXH2m8GSnYfZSIipKPry8lB0Kf+NEEXWzfFuc2+jjciuLoXEnM3HsHM5s+mdKIHuWdSIRntsk19w
nw3hFk7Q2KQmKkVVK2PuPKSnJu1CHTpa6PhA7rhjjqe9tUgFaXUXGAVVf/XB41Rgad2M6aR3o4iR
SvVrevfTIVDLOy1OIaRA3zGKZpT3patDJME90ePMybHFpSNxpVglJcbRQcV6dmhi025arYc67I1S
k2ZTyr/+CWOjLoQulhr0+PErk1NPWU+1tUFLNd8eraDmckFz+iistzpp85G0EanPtmAm2a68rr5s
BHy+W16Ra0/vepsocmQn95rBlEwbySn7SxGYoDL2A20m2lar34nzu5gp9kQ8Wch8NJTTC3qkxOe2
ALs/KuYOPb4gi+y1NY0Vcz4ONRywOYgtWCkGCRjBieMlamVvi8Y0Lf3fglkXowVislyOaHUahplI
dV5Le70QbaGIqttvVAfpl8CcuKVCluttnpN1IwejdifV7hM2j8whOShXn/2BNMiWnSuBPrtKiXw8
OsSIbdsPQY4wcTig20VhpiNkEHoviiIZSp7MJ6zsqITdyXt97bB+jmOOWsvykCQueuWqGHy99NyA
R0ctpUN8heO5Fxb0F9MyQuXGxIeQnup+ejV56iQCdHrZmfmyBWzitiJWag13CEYFRr2dHck9c6DR
JP5yKp7M+37sHVWmYj8Iuk0f0kSWqlZorgUGEnyIJ7/jTGQp9AbtbUrj2zFzC8TS7TlKcwjtLQe/
ZrrzpSs1QgwT9B8iEJDkDfD9WkCo4gLq8v90fvs7hqf3K3ANJ976KPARH5NOG6+Haw1J8J7azows
1aloiOXjIqOTX7X+bsvwF9N8y9xeTK69SFTNH9DPuKf4O9zvmEue2XE1ldBwxtKal0hpAYxwIHKj
rS00EHR4YEVYPCNBFgP7Cv1M5N3F5cnx/uXf0T/k+6+icWYd+kL9HbETfcEDTZxJ3uuxtW5n530U
wAxB9Wy+Gu2OliNV7PHA1x0eY52aUUVXyKDJUiPzdw/G9go9ZgdFNwEol27Pe6zLhz5QYZriROcP
uZJw9a4RPyi5i0aDSCT+/XIxm7q/foq6EHz0uImQKspAwHbOesomsa93grrOhjWWiwebSXfDcl23
kNYEWVaGMHZoVGB9ipHXAp5uzj/0PH/z3HjxWozI35jc4hbzBPCpgygO/0ynZAq1j+CrgFwOX4Pu
p+4mBemHSqpFeFdOnDAeG54I9iDLd0IGnkaXdgn+DzpsqYfA8Hk6rt+aqD8oOBCoYbCOBfU1UXbp
e1ZNufV8SBOA7uvhIDQ0ayzfv4+oLCNCoVMd/StT+Y0gGsE62UB03ASdaeI/QV0PGyYrTk1qL/wy
c6t9ERkklAGXeAxzkCZ8MH05PPvSFb19kplGByqecvILT9bJosk2TpmtuH767Q2VAXIMaebI7UM0
og/+mmnnqgM+VY6UxcoIZEaIu/2MiUcc3nONPzoFOHg/4kZZk782BkF+TdFiE8iRvkvRDXv21LzB
7NY8mRpWICwPUawJggsPVm9jUf/d7a5TCSfL831RJ3pHCUV9I3Qr6AUWzBGdKrrHeaROZ972n4TD
ZwXVmbv/dI0YndBYHvPm7PgWm8lQC2Gj52XHa1AYlXi2QQd//Q0BkNyV/f78wX6r8CUlDP8967sy
KG/bYBPyuptTZtgcrUDUBhzIaN6mE7cLETCU32Z/oi4+2s8IeR5NWWt2oBdkoW6sNC8vRxF4Jj/7
IvnoJseDVyV39JmSdUmYmvkHRDjbZFmP9MYTq8anO/cK2atpYHlPNCnuN3tXgyw2N1Hp8tnYhUba
w2XUOKubkj2K9vVwTCofehXOpFbOWhdF8kuDZ1EZsjuDkC+91CHQARLE+9Gs2wwIb3PHpQgsnSeW
V8Cni9wVoF1pMnT29te4IQmpKf99ivb8gxWSCNQUwy5WNJhuAwsOkbUw62Dv19IKg02cW+r6sOhU
T4ZZFjUJ4/Xsdi73BXZo3k1fGeq2HR0GpNWn3OKU63SEbYx2Ftnu1n5Mq52dM0xAGPZBK7s4B6cC
KpkGdyskDSdgoUkTHVJfwdM2CtaKWpRCwcbLBtilcK8t1NUSEb48oWFb6YoAdWFhyX7adfMZmxfa
HM+O49wbnZ8lrZy55HXvAfYD3X1KJ31VBc1Zha17T3uyWjH78wVZ5WHUkhqyxqb2yMiN2TwE9SaF
FtlbqrEo/E2LhyloF6BF47RqoBMW42lqlAXAWVI/JYpxCsSh2nGPx2ktlyTvpk22qBBl8G3PbPFX
MBiz8MzPhMKfUrbOPt4PDKNcp+AEw4ge+a6Ma/bOMA2MHUPAjj7NSx9L8LMWzIdjxIsSGl1gUay5
sx+D5Gk5+uijP8cM3Fz+qlfjFaapqSQi/IKa3Z7CdUEANTm9tdiHAeL17WpuFCkc9F4TWudXfGZZ
6og9UPwxIaWm08Vg64zh0TAmCLxLSOqFw3WaMYzVFLrbecTUxPetfz6oXg830KYOJKDkVSopHmHm
hMg25D5zmGvL9/i/sndlm0jDegcxjGn0ZfCTBEVkswd6GeOJutPrFNgqZ9KJrDovDIK48Whu9tTs
iadr2Sa7a3OAdHcmoapR3gTC5c6yGvW/7+Kz0j3DGbhUSiFow8tNL3nKSef98v/M4lQX03D6SjA+
UEXFQgj220oDPYsRMqxm2r8QCcdwC0sbj+u+UGivGqOEhKkPGJjOF4FPUwJn3p15n0h0i86Pof78
REyV1g2gsHC75F7iHIGxIs3BQdhp85UP0qsc2R9bcrsoKc3oTRpB0iCpxe1ehJ1GF3ctAxJPw559
a0iA2N9CB/1XmuCwfjDgQy23lgYq3PxxyvxM913CgEfR63ujbCHZcg8tRGlyp16Bs2KGNAVcUVT6
nPNxlSrb327IVKj2F07cAPiCZPU5iBsf9LTapZbWpHNu5x4agRusWnPLEdsMxTs5EyriYVRb6EFj
GfzlGNQAES8NBzA9zB6pDijLcGdOYXkRubDe512oB4UqBcRNMGX77lAJlVgJZg56kRlKtcSZ26gr
Qajq7C9NA3s0LMEfKxF2IOkFnlvqupkn8gnICAQygoholsF/r4r2FeUpZBJkm2PoaDKa8bCCKA6t
y9wZRlpVp5jRJP465hUDVf264NKvNUNzd6KIWcsSrTVyI+vwybXxLouhUFq0PZPaGzmSAUYIr6iF
A9vWhXA8z8ejIWhdqD4apvyWZRAGVsbUM0YlBtV7xa3/m7zgFUblp7A7w2VtQTjC1pBgWK6TyxzM
gMaUS2qqF27IFc8q8ZCBSThS0Lbn4l5i9RzAjhgNZeIRF2f+FMbM/wqIZKKUAPbvXBlgTqbsI0wt
+Nurfpe/x8its/t9oPofApuhFuvPceZWDX0dPcVGokOb1ktMNizniD4zrSCra19hZErxMl+M1FdU
PBxoCS4RmFbmjfI9GLDxs/EyKVBbNTh9JjVPcMTnbxW87KRfuA5S1FCexnuGwETmXAdcdVHqovuC
DZZw5QGKL/Rhjxnv+uIzLew8Drhf98EIAPm8/WWLc1IniLAEmj9qa/TjWXMEgfxUpKdZBEdgmHR6
DhVb9x6L+OCsh3enGgjvGUWnwVxkUTURN9ia7DEB+CJ7YwquieYvJC8OREGuIuG6IDhvgcoNt2FK
XJRx/sXPI2f0bdQnbhZ4KSHUQWn7vFMz9efxlNJ7v4gjk0I8fUOWUh6YhROEF2Q9qhMtRrSqRlrG
O/QfFhZ5uORJradIOiIBhZcaPrVSUEC7L3j/E9mipmuTBWGHJKhsTG4bxq/+pgJx1KOI4O/WnjsU
Qb87V94ySV/Tif+OXJyD9EqAp6RGwJ1HRNhmYRoZr2QstSiA/1xGlW7eNjY1FRSfGGspI9djJe9b
FN4OvfxfTvVBvRBfApYJbxsN7vZk1gh/VLzoIFVxRRK+ZmZN9YFy+iDqfOtYiOq9CYghcIdUWwT4
Lhiu0Byvv/5VQLcN5GYm8vzyK1cMZ8GOh2vGByqa1F0ZBRCJmedCzfCNYoTV6ajRud0DsTP2xS4c
wJS2RkIen6eulXTAfXKrHSg4ut6lBWbccc5cpIeFurqLsIHS992obNVQNv4nnG5yZcYU84MdolrT
664+jSSIo/6xI9XnTtvuSxagzYXGcZoWqnNvPPTWAxRY9s3WiyotnQ25bcwVFGz1If4y2+KJaghA
hCuBid3hUZL2Eo3eXd2Ymh3H3Gy5hY1SgwXx+OZjKjBC35VKoyJdIFy+ur5ztywPVOQ/0wVvde7Z
lWVtZm/TIqyRKvQCcU5cN+8PGXh010XqWYiEFa19Il9Cc2PvJr951z8yIJIlfp+uwJZFfovMd/Vt
xGJQ2nXLoFMvk/l1UQHfT+5tQzqoizfvwDZuW0Ju0yyx5JYcLhGIKRs36dgayvdm1t9r9U1xlipP
83YZlwCd1ZujIjpXjZJHqGltVdoYSYg/msCWEwh5MzNWxPXAV3mHml7YC6uS3AMWzGFfSijMSvY1
s1EQ9XV8XW21USTcJQnMg2zDq903IQ+XYTPHLCKeo+a9D9EX3Ik3V8M/UtoB8QgL0M5JXTQ7dSoA
TMEpgAHN4UjTYv0ufCRWsgo2lHW9mKjZTMRFYb5fw7Bp19X2K0kr443rwV1AiBldh8h+w5PsFC47
4ICRvLFypM2caJU5Sl8ft23+NBA2XUh/v2yDlVj6lqQYdODhTMl0DYiGk7HadRxafEUg3jQqXJuw
JJgzGb7QaQgiVg3kIdyc2Onya0cfTR5ii10XO/SAclnwcNUUNsSt1MrD8NAcBzWv3GYAJz7SAI2Y
AXUlzFug1QWWizGgTJ0OIzl+AgNxqluTIn8rshaUgtAEGryb8PxQIrepdzpToieAZarT99AqPpn8
clDBgAMw4KJD0VoGHLNPrUXwjQXw1LMMlImI8wjdSWeKJZSHtVhtDkP3iG/3a6T5nf5MAwmiS9I9
dF4HVgghw9vjJOfmDF6DCIumK6AdK0zxQ9LwI5qK14hWoz31bCms6D2A2xBkhtvo+NLFzR4kV309
KKjjmySea/aQweZcbtmr5JuJPZqRNJKOAt7vm8Bi4aAmmzEW/cpjAqZ1aRcOYfpgbE+UFDjDAptX
fQeYlZ+5mEqKG2hdfNXMqRfoqQXCDR0MKdth6iDolppwm6LckTpJrOXWGEpMDBJoXco4j3M/UD5R
eM8dKqlV8LfOfiEZZ0+SJISwbjseIGY/s3AOzX9xZG2GFn1qS0of6FlgDZb0I+MKCZsxvhMZDIvD
Z0Hb7c0mRi58QU/XNSJ0dD0NkbcPjJzEXKDy030HtxWujtnRjs4QB09FJn7a2UHMURDd2rprmJhP
DNbMtJkBSPSRIaLs4tHe+7p9poD2LvCndqx+rU5DvuMAluFqSXz02FVEa/hIN8Sy2AlBpK5FBV/4
wjqtaFp/7Sv1tuVq4cFD1stTiC1VD79+lHVwh251aolH+uDIDawst8uC97y+TKTYW5usQN3kEsL+
RToMWZtPaNOu/nxEgEY+DutEEjtx1yogIHoJVm+L8B8NdNfoW9zjR3nbB+/kyDpslf4ItBUlwpLa
Ar0K1W9cQuWClxkUvRk0ZGUQBROhrCaxCo/BqVxCMte/eYPqM6wBzOCEZdpH47eEn+0PNWlA0IBw
ZgJ87drpjJD6MM9TFnzCkIoePQyDKwjBN32tALy8l9gurhMyQgRj9D+3iPkLkxp/pErxn0FhKbKm
59XGvEZSf7+MakhYkvLpyA24W6EU53nRQcSpkd2IzVafI2jU1E2UgWcr3PLKdJL1sPoZTmqVQ2kZ
nA/69lOiYHjUHL4zHBnXQBNXUsKfccr9Ui/3qLdFZzCDLCF48juw4hvnticsdK5JVQz7blTlDcvF
Gir3RdP2Y4WuqoLTcumrHB1tlYhGV8u99eVAFzVphUTADr9itW5CQZ/iH5CAa1Qy55GZS7B/5ihI
2aZfUrVRrE2WEZPZA0S6MZde5INYZPhPDAX69qaiT0zgx1vXdia3QGJN3upi0axMflqhBx9Un/Fe
GS02p7kNFlmEBfc0eSl6Gox28Mnqea0bm1p5+rfmhzTXJfB2JzZksVFaX1ZAAmN0EOklRjBSG5UK
F4YPGGAcGMM3FsspK60MiZ8FtIqvIk7VCeE0b9zvj/nG/07StwqeieOUWouSck+b+vVnhfTXMXKH
JI8r0TNMSPWls1GzNj4sxjECya3bbJgUQK3tdbeEbBEJp5qcta2GscmA0HYEzTAXzdgi18toP/1W
inELYGggnU6N2WMa6XP2nPJIlh9+H0W1LFQuEdwFm08/FtmImtFU37egDSJ7qL5x3CaVWfXuzReS
WOEXp/2pG+y2l/VvYYyDBBRZ4mFRUkt93tU5K2PWtLUesr1m4RxtOmRPsM6QxbclPm7yNUO2ZnTw
6gvyatj+z40qcUFavC/+qOdhAxnuaSyHEbUxkuGp4UntDBCJF32tJrJI/hVgIw9Yr+AXQVHLYIJn
WHsDeuNCtlritlRfwNjodEs+AA8FsSAziE+IOMPWTUcaV3a/dVCZLZ+rrBxx/O/4t4tRpC5Q8aWW
TAnJex0XE5BRw4KFLmeEzb3kZIw5e5fQAe8UzkEEERBTWjsh0CGX9wq5CgasRn8miBaQkEFp1VAK
KxqwgNrTiGL9J6JkkMRjAyuEVbZwGpwMIjFLYstAl1F4WBEQVebjlN2hZlVaK3ZITBugnMUArPS8
FushQ151sFaRmgIsZICkegyh9LM0Xe6CYFPvC3wjW0vU8Iyi2A6sUANe+Ihvl0D7+40L5bPp7d+o
fhecibj2gt2HzM7e0+Tnjnc0GV0rwPBgQhX/sNcMS7obvYFj6U4sPHCzJlHPqq0URUqgbzcernjK
+Wo/3zsst+dLVAFSJcljA8nCHTIFSwFjMenum2xa70eoE04JSRr7KrvjBslWL8H2XjgqTLDu7eq9
ottUT2NHDjnHuaBMDPGXuIqRJmL55ozr9SsmYbnrXHHSOe3uqeqf86+ibIycaUscp5MHbulheAa+
j4PDePk6Yo2fBKdlLuoVmR6+qZb4G4TDcC38egJo7k+dHSXD/Rbw8y80vg3Kv/+lnQWjSg0cT2Vd
8bxoS3JtfZBWug6Hl6EoZdlW78lXRJicotw8U5BuyxVCTUZAfFs8ZurgZecepnAHX5zjY/CoETHy
ApD30Eor7s44Hj6ZopksesP3jo/6jIBGpK+Lca8a/JCPdzxlyIdVCIJgW52f04CFDeiky9eOUb85
HHyWI5FDF3g+FAqb59IRqZv7OktWx9xOZ4omH0ZqxHSO9KJVyHRVDhKXPfod0FNPC3gHqEEdzG/9
qOe3nGiCbe1/GkSayWTWFuFh6XTdDwcGXTnxu0bW/2fCn0tO5yr2F2gruUlh+cXI0+jEn7k/VyAh
dARygkGuOUQNeUyIa/osF1XgRPYIxgtM7UIatM/a+V4tV7vYHufSGm0JFlIsNOrXNRqxiSwufIUR
3Yot2TX67oJKbirliUsKDm1EJUDxKbljblo5VAN5UCiS+uNVTCpLj/4UqS/bUT6MW3zhELYLzHkc
2x1N0VpF0UW+Nhv+nGTnGQ8Nv51pYqsg3NjZqlp/gvWGcPIZXVqumfMCj3pSOiZQ/5ySMPH0Id9s
Mshw0KIk5xgoiymzxg+o8TtlG3DWxZZ2WXFNXncqdt5td9pdr5T0iJ/8P9J3o7Iyti2CSE0c0xAD
KpjpCQCxoeqzF1xiNU/1qyxB1ALZLw6VL0oyCPKal5H4DnEO42h46/NSzqH1L4Lv2nU1eqMTouKO
hnQ/CtySqJpf08iZ1KB5liaQdArJpl7gOqC4mnybyZF9/3hJG3W3n+yfIpa3JPtQHbBg4Gr1iLP/
DDdWguCHJOgmZIRIpFfomgkejwngQUPAb6XN/OpUbyBR40iqFPVYjnjoYgN5kujkKSKIfXk3/5TM
gB/C7iA4Kdgc7sbyeZMO+GFs+cc5KbDKOty6BSJPixQut5W78mgZaL0U6Yfc0ez/dfRrhM27zuo5
HbNknWoEmL6lDacq0mykIh+DoLL48wIVop1THfLywmCwDYTr/NWHKULo0YgDRcTDs4XYpGkLMV08
Sm5/5KQ9lDdTK6vK9PNEwe3kZ0zvPhpBw4TcM8oj7BW/uVPjJN4+9WQYEeMJaCyhzqb0Pc9LLJoX
f0sN2GCC9geg1gSg7DI357QtXUVa1YYsu2SiM5Acq5VY9vQ02qZi3C/wjMhxzFMoJuimnY2Ziq25
7tDWq3o9VB+pjrS+hIe9nK5DcMaN5IK/U+INXOEkSwOj90ZgfLQH64gz7DqKZdQFI8mz/jttgAPj
aNxAnL8iwF/O0igvCT67fOXCpbQa9yr6O1k0uqeLGlrx2EcWbGwxNJBQciEkdcO2iEmx4rfVQcLc
/Kw7s0dcp/P5H2HaPwsc4w2oWaybKLATb3EksAq6kEMURFbR9/NFN1gTCIeRlpW2JYA2NIYB1m6N
c9vf2cDR91WyNigi/C/KjIE879c75Cb+N8S7GAp0m2b8aMJ2RcuCsvlgjSxqdILCENGFoQkylnIA
e6guPUGFlRyGdv8QiJL9oSu3WowDvZdbsYglH7Q4RBrxuJrlrtAL8xK3n/WhJ9Pn1RlCMRFt9Wte
64QuhQisYyXnANk1AHiM1inUrw1/5EnnE3If8yAACCuc1W5wqTx8LcLYjNmKj6ym/ylYSMdBhef9
2uc5B9kHHIzEIgRCPAWOKXUNr5FroL2qlfwz5zDfQP/4AIhbAPM173gpWyXviiDloadE2wJNKuEh
rw058Cit0RVnPAVq0sunOuzQjfGO3V4y+aPKjtK98qAP7qqh7QlSJYrHLyvOZ9olbw4Iu5PVbVWF
O6Lxk7NZONstPXqXQDnm/ksuowZGo0ZaMXvEgD9phVy1vZSX7ImVBXB7j+XYj3wY7lH1UWrSLscJ
c/XM35c8LcSTIWE1QkkgSRVtb0jhXgDrC3hQ9A7/zRcBcUYGlGtzi7nKfL2W6soTPpHc1ZtVrHwy
ao/f7aKlZkc/XEkhGH2F82bYzSDkuE0ppl8H/44/2LXgXAgiKMPxoHmQfgXqRn09Hlt3zVrk1vIr
Vhzzg86RTno/sJNpdZ4gijYkCFIGAqvi5MO5iwlEdCjj7If9wYvD52JNUByAyOG8by1Up5GXhUVE
fF0DCZdzmp36xvEodTDs3ycoe0H8o3jR4q0QI00Ua/l6zktgn6tmTFwV/FTL5QGflUK0nUBsR+Qc
g0nt6htZIVxqIrVl5qhE983YdUSlEdxNzNzTidnOtWpA/XP64k2C8MqSQyaKsmdmh+HROck+Capw
aEasN4S8E0KbKWKfT8lZnjMegvW1FV0TcDdxWniP8P6ZPkBWGmjhFyZp9l54najh3WT6+ZaB4Yjr
YdC8cDexs4wE1gYs0837cJrqO/VHapYNPIjp6nhaW55JW6nRPsP/xibOY0vcSG+4z5SGyDsen0wQ
kEUXebVvHJMvWTiIH0k459Wrep767eClbJ/a1cm+9Ih9Ha0sZciCaKy2hm+z8c+5XMk/PruYg8M0
R1RYEGV1/MfdISdRnc2UvLFVFcIKJSoQbtHiQYj004oVk9Z3RUMnB4xGwMAvmEklOk+pLF1r6PUT
KakMKzNx1pR24O+RSE8KBm0i4djWYVuR34gwKx4uEWzepZ7VQTITOdLkbVVf9i1cjHuGnmKxXMkx
mHaMVtWO1PsdkCVMlnxilL3AFLfEBzkbobUHZ8Of6M8xSU4ksocdS57NWmh55WGl9VoFGGJ++QvA
9O93Y0FUBvzyShAYy6LpJVh0OnqnUtbifeOB73RpQH6d5WWyZhDY+FHmo5rATFsiTRkXnmxsrAbq
I1Wy/HeRUIap7dunhPgA304M7ZrJRMvc2lmCK7IK3YrNtUcw7rfzqCNbEheBRV2EXUbpV27ppb8D
PUzG90Xj1htN1MIpDLuneGjHblBjwVsSXU3nDOZIwZ2ZjHtQyiXXZUvqgzo0fB84jT1nW7WtjZ7L
k9j3WY8ftIGUk0H7RSUkKR/3TFyZcez5XcOGqKBuq5lllpoxgNhkaF5zItugke8pacsy/XgYnA0m
CD6phbw+ktT9nw2EkD1Fo75rs7RM/EElfUpiG6wq0ihufR9XdNIbAXWqixopAg0wBymwFSf54IPX
VNNbYynWHnXXalAvOIFHIH6YXlVjjNgUqAJCT0XcVuS64fV3xWNQEx48TF4Q0oYMtGFYVx+GZdv2
8jplw2dRUXwjWyx7uoIWkkPJDbZ+zd/ydhG+6Fobfmhg2UxmwETIY1Dvwbde+vRPWWiC4pYRpGBh
fuKH48jaqLLC2ZwDQ5kyS3PZe5NBoax/2NeV4o2Xu+wudAZ7ABpxeuMeAnQWg25XZ3V0HAzae5PQ
JatAkQmD3JyDWIUnTbKYFA5y8vD+b9Jv4HYxALXeGCi3r/al+TawV2Mr3rixqzfCDNR2RPuQFKCV
JOCvuh34Vm15ohIcnxFPTUyFO1AkriW8qHyGLwDeqUoYsiT1O370DdyrMh8KJNxIuBWsil+7ffBv
9laF32CQ0HZPgmx7dV0j55LkYiWtA5xWhwW6kBnWddQ65rRTq+XRVCSgXe2BTah/PO0QEIDv3LBy
cDqywW27P3OI9rwqXUsELF4UC+bFzgXV44ctx58KdDTv7DmL5L4VKrvN9gvzcyc/13tUGVYiaq+n
8lx8TnMLI9hj/rEetVLqnv3yIgKtJ9gf4AWkYmjiAvmFX2KrNV8oEY6qO2qIu6B5QDzDVOkIE4Jm
kCdFzGCfQSw3tYbH4sxS0WpTcFcTgiEDHfYMIcQcRjYKpqT9hqOG9MHzQE8wGViekeIJwMGgbts8
ImSRg88eV6v1k4Uz8dqRGuUoT72WbXzkv7ZprYz3gredKAWiIrta3knC3YyA6oZe+84dkg5imfZd
pDsBKFrtNLgTq2GT7+rPEhE6U4sHJRJWcE6CaEb3mFY50XjOR1Iw+rtGHQAPyC7MUuIMdnBcB4oS
4KpoqhoKDwexLhdLq2ip46SKcqXjMmBAzuw0NtdToWvWvMRVWz/Db4v7DtDAP/84QcSZibH7pH+4
MLtOGuFhvLeVNAx7NJgPzRLFnGs6euVo2jbT4uX0der5K6Rxv3lHg9dC7y6ZrRyT8PvH9Cpfs8ZT
Tjnhnjl4kozwvX5IuOjWw4yMty34hC+kn9ugGENQbCMhMLAAP2Z73AMQmM8lj1Ws7V4nronqYYve
zdFtcCRm5xsUQIQde6apfP91sUC//uNvq59NCqV/wh+W5cCVEDB3B2dNXq+bbgQQaKxDWma0V28g
Qflb15g3QXv0ZKb5gWpdCVnyoFXLrDSB5ta6oZ4F9wCFlLUA5V8G4pUWykDA7k8zNiIHFmZ8hKfv
B4Z0eJPYgpFS8Hc20vPQddvsUXScOkIDhQvyxnDuHbtvSJmtPZGgOIsVw7lTMK+OmMxaPAFRw625
dHTnDM9SLR/cPvdtDKgmYiRSitWTqetEZcPRglEdWL31w8a57Ub8AyxkzlvgbODB5jujuCukWRhC
eI7V959Rybo/IABZd/Bz8fiAtRIMyNTaZUVlv8KwZ+kHni6MMfIoUMVWY48LyxulvHQoQgvPM0uW
gG/eTqHfyFSomkdnW5qFwd1EL+KGao91WmNUXzlXHl3Lz/O/WQBwOIZOVjRO/feHDOOl7NBEFct2
kEdU/6XbOzvQAmHYgCbCTrkM5Wl4wuPgclwUREDNG0FwGq/4CszOqU12tUVpO8Br37+1qbJ9DtGZ
0DGk3BAMwWv3bzI2KxbB7m1sfwzofcGo9iBVTyvomvGmXODR3t94OuOXGKz+CutoTnschsxwRuUO
MdXQ6tdeIGNpayaq9eyBAhtdNnGiGaCNJlHZ8bDnlFDMCRMFes3pCJKBxcPB7Ma8Spqim1x7mVxV
GpSoGyMAYPs4/uCO0aE4NZ0BO9KFkt5hw8jY3n/CGFB+eNxPkTLKW2N+ex8DBBt7MDU5n0YbDE8z
Zn0e+5+Vzz1W8g/2LJDST7r4eYKcbdcxBqhl8/edeKgQxax1YWnk1tTpDWUxM8FpsIk7NaTQi+Zu
BN/Cid5pZk3J8ZCUqGsL+Im9Pf3xUB2BWsXoLTcrvcOloeqJHQG9RzSYwovLo4gmJS86AKOWaT1g
JVxOrATZGH02lyXZ+fVBTNYo3tmx1uh7VEooLFuDauntDKIlANHIHZnGUNlaIQl/he+HNvbNtMYH
iZqm7lVmRYMMFgQ+RjrGLcnb8rPCLUHVsYehI0gkx2sov+UIOFPKIfeRCYZ6AACEMaocosggqefh
as53R1sgS4stoZsicZIXp7SwBC0DMKuLcAjob0ZgW2oNXhTlI27J41YjOvV4AGHM493y3ZxOgg6p
BhXgJKOtB7Rshfwa23TPi64k8L2m8RQ0Q9Rwxds44qMtyffhRCIkwykiSE7hZsd3vI0adcABepUA
QMYzKVJhuBzMfwq7vdgb29fFJu47SAIIjjaioMWdIRsHNYxT+ZC6bDC6DEivnsVj6stk1SJsY4Ek
vCBNDoRzVhlp+WfsiF5LihxwQGI4t8BjJtD44kG5xo0aGGNOTmC3f7XM8e5jHYUHTQGn+8SIaRc2
nIyc6coOzHVZAOqdw5AG48kpD06o3QgwJ2esvQzhroNu8x8FBGTNSnI8Z6pubSxnnhtiukdRRvD+
djhzFL1wl0H7M6CXd9OAZ0A3gYfCPtCVNPQLfXZpNVMxik1XF2eJ+SSuYegZYfb+AcATKh9j8XCN
7DRPOz7r5VKRdpBEyofYiRFjO07F3Z0VhhMApPohujx53D3km/y4tAQJ/HaCrcRUP8SRZOIpU37T
E3ZbZuKz4DnOpcyEKKCD4PsqrQNY+nGW4+uIEjZTcg2Usl8HHB+rbZXsXgc+dSTrdE/iunmT2dmm
loQjHHRjklHUFDs8DZRtxkujXsWmqhXUGv+ml0EP9VPTcrGDmSDVQi3pCDrGYKcSSLoe/elUFWWQ
zPgk35Rll6/9huCJlTD1B+ntvXT7GZNP4gcMJYGVbGyOJntnSfrgg94N6fX3tZYY4IyHxVpisevu
8ldKNw07f9HFxmcie25zC9Qksbqp/Ew6g3BJPDkf9O+TEbI195uwUyYFQH+1yLt5vut9DUHRT971
Dm5uXKWR0S2i/726nSELNlZX/Cb+Lb9qq/uMrdGSrQji4m+lZ2rluM3Lu7f5n9vilmgsUdZsrd8n
4AE+5mWSz6jFR4msALBC4Zu1ukJChexJTuagFBBqPVJimY5MINnSPvsNcQYKg5JPIf64lPU8jTNP
BM7kIVC03hZVqDcES+JfXPMLuddrJZoGkSz42wXFF1Qait9IU91Pq22tB/+v/lYVu6eX5Dgr120h
bFqMLwm/xq4i/kFJHXEDEG916qREDTO7hIerCIPtuA8jyMCxTqS2o+XBTA83aJ/ZpY4g8cBzaqpj
XiPa7ea/Rmu9HwEBO4EzMAL179YbhMmseH6FKClT/pddax78J7/E+LbDvbTGMCne8JLBW5IBa37X
S+2pAV9u6oePmcMPWorKRxUTWuoJ2ZGOGyRnhFP9Oeg3uFed134gA9gzsf0giJIgWrK/1wfwwFLL
pYgVUzGEA0N5VGiExIVWto+qOz/sjv3xF262KMaQZf93nwm/qlHaGL/FuncjWN0rou0h0xw0yxUd
q32V1XW1TK5+HQmEZ2AtnjLdiRYLzmDazrtFTDpy+47lmCJBO3k/n6dWl3RyyZ2EszSkp8daA0Qj
XtqpruEKjE6DfiaivPFxLEArQkDU1dNpiT4WkbmLRk+ppgvsECdE4UqwGbKdOvPWEC85fQPnMmdg
tB4GUqeVSQNY78GmeA1fG0jfteoFkZEE0R7+qblm3gj/9UdyzUFYwZj6blUA7+iXrwyblBQp2OAF
0Nzccz3cKYNy5QOQJkQerRZfzkbZlXyCRUf8lc3oAKq3hr1e46gxa1Me2WqegzdRlAqd+pK/hALp
qUKZ5JZBeDvyJdzA64xLrvfeazOgVq+TBO55FBS4uD5lPynOs1LSkvsJ8v+5W9mvuGWL72oksr6a
hs370szCj2LFtSSfIde7Yh7X4geUhJKdtsvorYg9aMkFzs+ZSLEeLObwrwdDCclicE0CAEzOf7fr
3MGIQ3TuOtpLESkodgEXtqWRoetYHG27iNQhxkOErmE2nEV6NTZkhimwtQnemjfkKSow1/WHp+MR
TMSvO+diNLUp0Y+qt5w+m4TeHp+GWR46/X94JL/YGsPK/Jh1YvXTz2oR8nykvCaESoamWGpmI7y5
rgICNLz0rHvyhxkf/YzfXwhqTzxSPSpAELqOGqKH2hTUTUJVl7y4m/mVvmnU8aAWkLsCsLMsICF+
RPdfRX21oaJ03SkzERX/5gWlmvln8C2/ZVWIRZPbM2cI1CBCM8EOVkOxC01lBhiEndgw6zMn6Yle
MzVHtGNZbDraBtwPq+KrNq6LKbikHwvS7G1fou714XpMWJWUwEOL0wLCsBMcbOY5LwIuxectKEgZ
/JhbP5CC4cPhRs1P4lHVocEhRIUz4SBsTwJcaX9O9/7L06g5oR9HN5SuuNq7VZj6d6psGs2TtVYv
BbRSiV3Az1zKblsH28KZE/05q0ikp1XzjXwDvDnkFeJmomQS8SOH0IUQWs9yFZmG6o6y5kVJgdE9
VNiEnCqCXMeQgUMuzm1F42UyYsU//GXMoun1pXz9AqSXhZma8qzzFqQSXRjuetFo66/M/H0i1mvn
u+SNoyarAdWjmTw3K79Wy9czFEuMe24nu8gCIpYXOn/AJ0IG6UV3aRXNTqdG/D30H6mBj+Tko9HD
i8AvvRdY1+m6O8wQCc/U/cmlhErKzebyj8ujKPABHwZmbDfO1DXDaYUacWHIQyQkAcdvqBDYWwW/
oGCblnPupfcsDG+b++F2xVylTFn4nPRA1mVSpJLQmiIR+IaMAX3PP3nk71KdKswySBX46XhJQ++F
lHstcuxuk9AxYRcu+Fd5kKYQ+xt4uoZzSyATMgYEEQV18DmbulQ2lNuqkxUeDAEGwgSgYRoUiBVQ
tnrMvjP0uMn1wOYx9g+PCAqTjbCoSCQh72fIYnFnonZT+RvIRFWrFk1OtN+67PrVnjsAXPJGsSKQ
De+P0PbdexFeZnfG3oyFdzo40mkTIZvigzGSoMeBwWQi4DFZjicwCgy5v5V8gIpPexmCODJRVc2h
7cYNFGcKkaLsKvNcSDjyATBcGkx1u5XLkj/fhdo4FYst9XVu79T5iU+E3p6L6XQwDqhSKO6sfE1/
+rNf5WNb47XjIKyBZN1Xy9x2w7/ft7jpD+jBr57xo6spavF3XonjsZSDGHI0Qfal+X2DLLNCF+h+
H/Vt75Ozh64Ke8527ojbfBs6i6/btryuAfmpwCi8bm7Iym3FOCQKlyrx9117Z+wui3XcCZjgVidV
1jp5N0Pl1qT4Xh5ra6f1WFLWRjrnBVM5COxAbYQHnLU5tLd9bys4hQKFdcg2D+3azzJKmnONWdMn
BQoLsU4ym74FJBH0i/+RjG4TQFtBERcmnHBDbQ3FSa4o2QXGyYcsLnVW7JF+MqDoQ0CPvOJcWjwQ
vOQwaK+bMVzW8Fxvxsl6EBHz/scrkwyo+WBVMpZSbIatgIQZi2KDWxcc8ZpN+IsvkeiIf5OltXZj
w/f95bYtCfNbpSfR1SyQbbpO3m6h7hY7SPAxKI6qw7ZwF6ageXv+wW4SnO8DzlllnHTJBY7wOa7p
eWus/nluPD/QXI6Pc6jv2zzmiStaJkQF37SLbqcJ221LaAHfJTE65qD+SqqQHn0fP7TF4uO9JvU6
+id+SAoCvar5jrCzasHfjfRXai3+/7vStnK0CRBS+k0sHqHaIM7pSotqA6+kiABqC78aY1bjKgnd
9hVKWWPgvZoZ+BTym1enAUonxLKItu6MmAkOo0TtFkKdycYaZg2EZu1mniBUjxfiSkiD+UL+oK5y
w0cPn8NT0Y3B+hYYMFBUB9N4RfpBCG4X6xg/EuJk1trlTuHeiESG5SGugj1ivbib+97l4ST0NHZE
Y1Gw6hkYnIvRHaMa79+65ldwbOW+WxxVpoKOA2kMZK/ER2SW1DafvuPbPYxaVjo7nMB/KYJZdand
UII5fBOocvvl764xdha+MZ3B/H6hbshSV2TE1jWECO2+5f6UeTEMP4/9svhfbWggEedVFv25+fd5
dmAO2czsfBLY8Uzr/PNFNWjlroLp2x45RuJ6oAiQ502BWZxmtXfkgNbTdDH2ciUDkqX927v4kOmr
MhGU4WWwJhQ6iQwEbQosH9CMPMXckHzqTz62dBKWmib61ZKnKUc7C3pZZIZuVcSFT5cnqEoTYAxr
z7DnSXnk9dagttHhWJcme+C/bID9DzkhS12SgO+pzusi+m+Bphe/ni2txdPyWvsBg8t5EOTIn25q
leMgTNoJmlsiJE2qapFvXHjyprCPMVBgzo41zf2VGm8MAis1E0anW/HdlI1NqbrKuwFYEb+bmbNZ
mWL+xpwef4f8wwQYOsqIJ9u8P/CeDlfgPlhMKbztCNhmjwnoARLMOGi/vU1D7bPQYzHI5bh1uG7n
Eh1+kbdR00WXqi4KGufmguMHPcMIPw+gtDxpLcRNH5yIPvL0dAqvTWNZIpjNczRHmE+G3kIxapiY
ajUPcCnG83nbsJ2CJjONa6B3CFMg1RnhnpPzsHSldzEvVEGXGQeVwUqFBI6MJB2XTcug1jS+BLwp
QmXPcanc4NMzSZ1kaIP1I6VnrJJOzWn+A5Ebf1MOr8SLXVyakiCJNZz1F4xUAtgcWvTkLnTcRXVZ
MEXrZ+SCBmqr5yTY9cVE8l4PS60QRH8Ln7MMtmzX+2G1pdUowHl6f8RMJgnTq1Dz1IqbZso0Nc4t
259mzFA3VFRV/tlRUVPdBcxQvsQoJ5wwXW52EpgyrDWV9Kzy2gCHIpO+slo+e7nlSrlKkB0YppK3
OWj58FIzqlelfI6r78boIxLFnxPttFzXj9wQStrNiqIX0Ir0KsqDfK58DmAncITjfBgfe33qcqNd
QEHoesJ0sNbv1wWHKV+r9aSY6u7I3tzSw3IUjhgLo6CYt+yVveNG0GZC1Ys4Tv4QW+J9Wcwtkv8k
B87WQ4wO+kZgjhpbPodAzTStJ0p6bUEdYqa5BkHSSu3yRirozNXTeXwrbG/7JG+4WO/vriQASq52
ZHglPNQKIGn9vf26lh7p/l046DAQJvU/9ORF/2FyEhL8RId0qaBhNb37j+lRhdTzrYmo4WxbOsem
GTDMlwaub9yZ3JNcPQM5ZIMavInz6dpnhDpMS4n95yFjQr6JajYyfzxCx49kjGJSRebYc1aYbfYJ
XLabfeVU7YAowStTC3E634Y71Qkd6JfNUzK7rzc/pXiWUPEJVG9BThD9ZrbHdMh3BoNFCZG00VzH
eUeBCZhbwrJlfA5KQ6x5ko3Z2XjNLdF82NmStbxl2HC+ZEFwvmpnl4P2m/pTkKHRZkTo1hPPMYTu
LQoTN66afnD/TtK44C3dTxrT2K91FxiggAIOgrkdWkfUkJBrQdh8v1ROMEMNwOub++sfU7BeizzB
glZy3dfeQkgtMwHEpO4ICWXrGrvwEl6jhKrGotr5H6wHnJ0gsgC/jDdAQybB5C+R038+d/TD2Q4T
mlJVW/0NCxKlLHRv8SysfFByK5hV6HtNCjjWrahOKlRg6oYFcXJ3Px69Y+ZGf41tFkFXvO9N9Wsl
qM9dnQjmNAtwLFTNksiPhNsuT0lLd2hPt5xQI5u6sih3cRgy5G2HwZ67LPShsDjTM8pSbJbuilYd
u5nztsDu1Jv/5k6Nt1+FDDyktOyUZ/2lxeFEQFCAO4cPJkanD9t4A85UEvN2tT+7OdZd3L9bBjWP
dlGws8rtioxc9SZCsY7Hk/tOLVMbOUw6CxabG1QHcK8XnuYAmot9ArJw8lzW3lFpVFydZ1LA9H6c
bT9udkocJYCUw8sbhKBQBuX7rTuvovL4Hx6TD/aNeJnjJV4etvbiiol1q7KkjAUBwmjaFPJcr7Yt
VcvZjOnfNrZNf4rVcL8WbLyYqEX2YDuf28D7ycEBqmJz1cxdv/QB49dw7awDNNS0jyqrFiWGPxKK
/YHgcW2e3zXug9OGy9tprT5se1/jhqhWp0tcUeFTheKXrUQiHfnv1IgkpQrBskO+Fa79hicUTL9Y
2qhq7bQIi/BIcPvG+PY1eAO9onziZKpwSq29skUQ+cfPJS6fa36fWi8+kP9322KEUndASzysCyET
xL2BLmRjT2EzTFfpM+F81f82MGadP03TrK9E27rmqFgVELJgvOsXLK7vuOsWgdhyadlfKtYbaiVg
Mmegj+5SeU1y8ExSYFXhgfvqND5dDNTNiSTbIqfk+8wTKdv63YlxKQb4W4qt5J0vq4uWa36K1l4A
dGLo9Pgm1uu5RKuBKMfM6FBKbb/n7vXqkIH+gS1zVWGzlfjoxlR4qJIRqzjc6d1dKncV+CYbzr/i
LA14qP+nuyvsufCpFFsbTxXo3gfFOoN/aKbinHE+lNtMhDLNNpXJrU7vmGXWoOPRKdw/DL7+Rdg6
k1uzHcXQMqtLYgpsxhgc9T+B7OXbNmJXM1XbMJu/sy4Dk5K90koQCT8/a1jm7nxKpJg6THrzGypW
29dxHeltiQccJvFUPBg+3+sL05hTP1ZjczPZsLm4y41hzceQQOMAxI+PK631mKa+R13TGYsxs76e
JdAvuArftLVxQcwhkP8ktjzKl38HkLsf85i84girWq/0ONc9e901eev5ILHjL/b7xh2SCPIsxday
0ZnJn0Osv52A2uq+NcHB0+jKGf3Zai09vZy0kzhRjbFwIJ3p7l8fmQCmftETJM34szqP5Txkig7K
Inm9lXIEUO6RcbbOXbz0u6SK9qBUErRDUeMcrjpinMjVXKw+elPXdjzM+vBnmAwqegrv87Jl0vk9
1iR/PQ9HjOi6Zk3g/NEwzijIs+o63SLhIyj7K0VRnEbkoED2lJKpLP8XJ84tfr0/1aBzxDufmRc2
OYOeCNH+Y5fRGBPKzTyOlqLRgGggrGq9xqd6cHiOTHqoQvQOK5kExkn3fLsjM/9jIVKBOcIntY3B
SmOo+4v0eoSmp5EXMnIMCdBjFj9MWRRNtjFojiYjhBOBA6QAZpg3rHmcq84s29s7ps3Fh0TAyCk6
f7IXQiR0bg9EtU5F7dB3iB5pE1a1aloxJ7899R7JlTcUmYwi38Hm4d51wEMs6czD56PWyPFIxPFm
CMk7L/Ugsw5EwxhC28gRYCno069gKb676Nr2cD4pP6xjxMeh3+NsPFlj028yt7kK9VfWlfRppXzb
g2ip4JuAVemTlxvffQXe4BQxfJXHqfsTZytZa0g6LkkcSzeZ2uloCT46Gm9KXo8WbR/Wwb3vSdS3
c9hQndYla9wAQAWgWFNoB4tYX20YpE5IVEu/ISrA4evlKob/0CHNVTiZMSc8sdUadSOkcR+k1eEH
8ig1/tZliTHDTaUlVfqYew+Ne2DXr7hEijo57DHVxacLDFeQdkN4pdmheBk7nKmw+IglWIBNRusl
AaKBA7xxz8NTMIQ8+k0yaOeV5TH9B7srapPcvqMFHU88gqhQi+xFNHmkGvwY0NCQuJCrw39lv1dc
wgch0tPV++ORS4zn3HkDjj8wfKZ7nJjAyqyrBNkTtw+/8HzY+ZmnrKZVtXvisUo+0j7XZShkd58y
9KmQLEdNVGTzwo5PG6C+JxZ6haAuBuAG5McB8Az0T902V6xqcHdkg4hqqFVxtce+iw2VdVHHAFxU
hDf2rzk6Wuh1s1y/5r9nF5dABlf69bp6WVCo3nqKXEP/B6ZER9HhMPv1Dlzsfk9Snvj1n0p2A3oP
V0CVxngpDl1jXHO1YC6dl2GsztmtzSVBJi2Iz3YNbH/m+pSvTZYERZPaOep7jOdcEbYGVsqOV+bl
rfFVkc63dsdNLCExMLYDHUjGHrsqwNjE9jzwLNMY8gNCtG2djVEoaK/w/+mzeXaiKh4KBN4V8ybd
tEannWX5qUjmie6pyo6pg7wzoQOY9dl2WKav52HH/MyxANAoSWtrwwYaQmMmoPL1H9uF577hAMas
q2HEzg3ivxq3aC0V/EeiXO5We0NVxwKYkteARLbmEQDEl0037lrN/FUGyoKG9xcpSmORZufmZaWy
J+UdtRZzlW6lCPknhYkREb1Ly1XnWjzRD1smHelvmoAQ+vMFIAb+OGwizyMJW+4LunabRVoEQgD1
UibaDUsa6Ws24HCOj4mgufCe4MhzqDFXLAVQLEiWV2bjEgtN2W415OuX1vtDt44yvOyYt9Z2M2kT
zpMXtHXcTIaPqxMjbo+IvnfzM01jl9sX1vtGFKaQ6oEfQrmZ8QUCpjnJvKoQyD0mhVVp3+kax/3e
L9Y+crLdMfm0kPBEhZkbX0IvNWtfT771tScSBNMMvpIhMxOh8sRYLUrkjocOATYl2q61T9rCnMDi
ixe1vl6pFcFJp9W6e2m+bKIQyQJsAXptxBizQd3b/pI77HeUC4x7oPWLsnBoqN8rIcpBqpCPwuRS
C12tS5/iLbIIsjL0J/oYdhJ/c3UZuek8ZkZ/51lh4j4IudHRqjd2czWhWiERZCT14m7WKd51gB9b
sdpc1Eveyu2gRDcoDM40/JnH7t7tqpmhScXIh1bZYO5f126NZ3FoWjsDObUK9SvlRuEb72qeZaOY
WTVb+PPevnSJasX8r1e9kNDl9kklF8zv9BzYN2b11ZLgTVbdjmsgcBA7IBlmUq/tSjsSugTV1PSe
3fwuHY13P99KVo4qEnzyxf08YzfcUjC9l1PPVS5ls9IoZt4dSaFpXRGYN/77D1JRT846TVQ0QFtZ
TTwNytvSv2JWEbYBcNqVjB4REs4NaR5caxUVCLgL45Y65aK5OiLd5EFppZ4saC7ia669F1NL7+Li
bdWACOf144pSKGGvcAVStG9xrO4MtlnUlli0zhYyVYrGsxhBQP9y2JAxobSKC8SsJKnrN0dWtopS
iP7AKbY+JWL4T0RlXF1kGijw7ETdQfvrmNDjL9WDjFIPqxUn8h6+bvjhvvwzOe2GKla2qZesoyle
icIDceR3R63iSKMmPeOfXbCJ6qXtw7KrDp4TT55tEx3+Lvwqj2lpALDU1SfBXNdWa/CcfFYSgYbV
ZqXRVEWfojDmHABKc5bdsbjZYK7h7vWRtjebAOu5fai8rtg97NqYnjW2PdFxXztiuJAPtdRHQaLq
w2iPVLfKN1twKFkdfvTTpxL1GQip1VlqPDOHZ7xPg2vTaVrqBMclZ11iw2DmM3tjXFOq2olHdayQ
Ev+d0njGwwluQRpMarqcO4mbwe/gYQteQQo3SsLE3/q/3kbaCR9flyb9Vh0/qYH3soT4407Xw550
Gqs3vihxBqlWBIrNxF9G0xU2cDzeiC/ZwPlKysCmntiFpbhkk+rppMIWXWutBlbNUo65Bl3hViEZ
+QcxzQP8CVRLQXMjMAOv7HU/bOkIAhml+B/LGqo49DbDnDcPS3TH3HAEvEAtl32z7i7JNd7Z6zrr
a25zs0Vu7Box0b5svzjXUng8zNvxISHNgw8Sc8WfZmtzTW+erd0OMdH9keWWK+vqb8BmQtr0sMH7
yZaibmNC6Su0jlC4EVYriRzCnNOKfFpK/5Wq0QJ9/DNj3CbTxvxrlQ7l8R+sUrMDm/JUDZ3cnik/
B7RfB1UTKjqzvclNpGynHwr7QARnPW/Cu0neaV3DqbI6C2RoOGzaNjCAx1q25l9bGK516KwXv8Jn
AS7EHA9GEji8VeqQcjI9F79kgv4godKTgamBQP+2CgIl9HumEISr1ogtezTn0fKB4uzKX4gcWeeW
+r45xjtL45pNEjfEGj8Kot60Ad5fixaM2/rzkbeYpEpqFf7cEaUw2pBgTqTsumM6PD3vn7omhz10
A0fmJKHBjIw+S/YV7zFn13Fk9bOgDYGrozD8M7Hmb9LnoyWMQoQIJ/sOfx+LEsvgq0xCruN3sm0z
cOYk6jSq790LjHUclavU+d5tSr6qe71avY2igwi9ocjhiW+m/L3GxT1Px7QaUOjZSe0GtuMtuqZA
DyqevEYwn9lZ4IeAMEifdBRlpHf0dYdV70NrpuIO2/4NyfVcglWQqb1GNkweZtucnU7kmO4kYLzz
RY0RvMYXFdD/jtJoPmu2kSkyV16PxEZiklFWy1jTVSeYnvNEhIogIrc79BPloL1QMQFnVz8eMdV5
xMT/Rm/JA9LRqYX+Jhe6k3aIhTMXG8sutdBWuQDbD92MqtyASdSLM/LpZiUWk7zBF275YHq4YTga
QgAHZGhb8yXFU/AQigyD1oBaDGrxkWEW6DLVNP9JNjQyl3tkNYQO+fDr/Ir2jyeDPeX2ff5rlwBi
nGRQ0z0CadXLzEysd2TVwJ8z4lVJ++iDkJgw+jgqR2O2ZdNxUCzoz9mxYiFEBnlyp/AsEY5cV1lC
E8h7EwSP3KUA9walpQ/IAWUB4TBtiqSt+T2PR9WKtE1DeaNuRGnvZGxxyW+O1FEi2aacIJIsH1cq
c2zFMuS808Q/SBZFN4Dww0JYXbPEZA6Dyn5OPSFNXKyLmaWKZVVHuqjvZAfLHDqzR449v8DBgiCo
3KjmEGU14Lq1O49LxiQCtH/pUusdANK35db4NL6YLLKXApsHs2VIfB+Kw+Zm/35vXew3JWcTvh64
CiSpmWm2jbMYKvk1LrCKu99CzMOGsb9SyCYbU7W3Z2KRvUDPmLzc/ortcTCm5zBIm87OoRxG2oPX
k9BCiK4HLAbBQ9VEjAkETregfZQPQs9Du96N+Uz3PgeR/ZjZOQr32lYNCFu3axvecI6xb9BnmscP
Weyjy8xA6sFvH7cO/i2aOfJkV/ztJXhr7XIP+QLZxJLPfkZ4wjvt6HNAoSQlSW+9/4UhbhOqAnDG
Mv+j9WdWZ78cH7Sm5XoRafFgv/xUR+79izuh2JwmaXInAGu07cAbIqDFbzbGFEsTOsXUPTtMdpm7
D1Ipdpz/JAH1P6iu40IxWV1VqbB3qHL06iJEEkldaOn+ne+v0DOCtNIdxB7pwz+ZmAQv7U8ZrDOA
bDQUkPK53LAtqlLMw2hUY0yukMOphOW+7GMo1mcWiNPwgGAtQeplUWVsn7FLxPGbHVQxChguOe8m
LZdth6eJk7of/koj/ck4l0XfJFBy27wShc00hrj6tt4oWyiW6O/SvTKZQ4ACaZpj3XKOCPtGJzBn
Ei9S8vH4k+VewYnTAslKoiWgECbhsx+MfxozcAoHVZvC5FS2XvwJ0Z1W1b3eLLDrY/yZ0OyPJ17r
vJPIS5PKnxTniIfvlf6O8OCV2ndE6/WoncOIkHExj4Ss/Q2vwYVIfXyiA+ZXdJK2PFJC02boL9aC
6fWJN8GYoRlsZyE0zS6x6wTJiuiCpnlx20PnRhi0lZyALp19hlSb3NxTRGk9G9moRvd0zth3+mI5
mP+JHiYnzuuELeHE60qSixzbZduoR97lF/4Lvw+fP6QVC6dLGzHuEvUa5uGn1k9gq9PgoDvvcf9v
1EG2istA7TZDuHLX90W5GAAY48ENCsJ/R+5KKw7LEgk/G9b37a4MheZ8CImysMfL5ny3LzzSaKHd
7m6NbSi6UMtAeSL3UOYwofXpx+Q4UxGYX3GP7l2YnXpOLWV8yQf1VtpPGvIqICbCScHD56LhruSo
Hv5H+rPnAseHktn26OW3tW22GQ9MsjM3PBstRqr52DGeeqKTUEATtk4DOSOS522op8tIrjnm0chm
pbLQrfK0qFnk+PP2bbMxL50AUkZ2k9eYUDtGrk9yRDJJetv4jWfSZWAsOe8MVjqYFoFsoGwCc9d6
flSh7xE/6rwZdaJsdBgmbph96r+CVqUIq2q+uy87kkl4mlJaQAlzyPB64dzKusQRhFwJTkjWLXas
4/FclKG7ba/xfW1Xag47RvYGmfnoLgPbXkp+VUEBy84xULJ+P9brjhn5JTFRIvP1+LFfu+XZovBm
XY1fvXg7y2Ne8EPVEVo5ZLZhNh53IUbKYor48/S8holDc0U+gOdB4gRgeEQo5qtJWF72l0DYXpGa
IhqayTxuvhyviVtwo43BJlifpNnFk88569k4cbDaG8YOfdHN6bKm3ZBc956rDX0UJuY3dIYl6qjv
RfWmgoIpedr+EMLRlsVZayn8zLxwEQ/DMPHGExiZdq8m8tN7QS+YuAb3VWaCazNmecuHRhy6DX5r
rmBWzwlamnaW/FgJfKKxB/zt/cjpONAH9x3YXBAMMPTKw5wnO4lLeLT35dK6ouXOZjSk8VrBM1Nv
xhl6QODA91hn3uQyrx8Z0U/F3zc+IL7cLMlHrke/jh4TwC2VmlpfbVHE0EXjRt4oohGSCYA27Jtq
/bma7iVhgtFxmdUtXHGHHb06bAIVBRM763wlvMIbOC9s8ZM+Y1W/FtS8q+Xw6mhSy4+NZ1bnNxnD
4zWyTAp/ksFQ2AGjgznIrWdW5bL51nUntdQgum/qUEEnP+Bod5c2huFr00KhRPBa45l+bylnKcwU
AlAM9M/FpeWKYEwjRQic4NDzn9gyomBM+5ak1Knx63BZDwz1FTEfGFeGgFuFEsS+eyonNSANe3yi
DcXgIaVnZiErvyCtmB5dl+vyEEuaxalzVIwDBm82QPFrts2TC95RjGVrZKul23ywuK7lvgpdVHjL
jyzdxh6AtLR3HaabRBN7Oy5n0jxZmt3m6NGjMtSDfxZu1dkpdME9HZ4LXUa3UEdXuo5GSKNbTWVS
UnR5CsD8zgRGYJevai3yf0asJ9WbIiwc0+4TYR6UHq5kR/nYSDlS0d+2+j4qUOT28yCVb5vgWDnC
175K777Dw3BxGdjMUnHofVB6JnmRqtBiIPbVMDMcMGzJk+2H5tFBye/bnxcwVcfu4A5PSlSSVv8m
qcrBe6euVKmCriV8pITNC4BA0dmobODrMILX/cVQQkpWqW2ubUnNG6BS1bzrNkyMZPEbqOWXRw57
XwQvbQV7ij04E2Aq/adR/uSOqseGmQy/hb33U4q6T5HBxinLLrAhcYIA1Ppozp6fTNxJNB65vXMu
1wsjMR+NRJIMppa0B3ChnKWzIu32CAq2bMhb0ExBBYzJA3sh/fdUcr2SIOI5t8qFBoC/HIHUADfz
UBHDXRG1g+5VEveNteg2lFS7+aZR4RPhCkMj97DLN3rlKENNG4ResJPgRpeyXeJ+TCFzi6z9EPg4
bG6MnMxOrRR+1KFzka6tYp2XfLEdWsKwDpMSEtS7MUpvgeNRMYORvLWNeh4OCgnzWlssLJxEgxuA
AKamZdrntOB0Uh6A4+QcWvzPnyid2FXdPrqTZN0YAGvKxbKBo9/eC9ClZkAvtWQj9kV//iBrQia2
6DBXHhycZ9gMEWmpRqin3+WBu8Ir9flJlMLIq6hgeyH16gpdvNykwSAZRkegNEqkEp8amLnWDgtv
veA2MVb0ocIIPsgneiBBCvOxQyFgZroFsKb9Ey/drJ/4HBPn0ZNUWVPZHHAOnLvNN89vXN2dQ0D5
cx98Svz1u0cAK7Uv+Vvl7BovjnzuhJeQ9bWDzvjw2/PhxG6EaWqcc8XUU1iKxsrRISSPDRlQln/N
QF/EYPuUs+k58t1jHmvwLIxqzZnpl3+vqgqn1QzBOQX5PE/H9fVyZe9RtFU+T1Td6qyeafhkHBHZ
8bxWVppTKwxFXt2BGxKlhacZLhCjJkzRJK643WZQb0Gn6EIo9B1tP3GUM7pNAhPhgMXA5Ort3F5e
jyqOcWy771XZ/bSVFSkB545j05ViW3giVlWnG/VPFj0j59aNLyGFdIa01782w684Ck090wy38NUq
TXiZrg2cHk/GEDkIgsxYT54wDEjvxIdpnCuCbFdan0als9dYyDEoRqdpX7Ea+taOIhQo9vsOG/4U
YJoyfeeHLxtkEs1r9I67oQ+YnO3gXSxKxyZRK67aRA2UWhOM4YuLklMH3FoGLnWn8mV6moyE8i7V
tZYNFmIozDzOFgOB7WHgl04K13cLGR6NtczWo70K1k5lt/BHmckwY7fmtZB1QkJ1MSkhqajCW+aZ
C0/Bf5UvUxEfhjSJu67rcXAhaEOF/WVJq98sC7cTbo+AgbF3KlgI9LRjn3i4ajM08RIJP+jrCALM
wgtl6YArb+fwOW30SpRP8Bh6x8n8rcizpcLBbDLBlasj7Vh3ynTtQD9+AS/2UZkbzGTjHn+yfXT0
M49EGT74Xo4i9rXcWLzckn87tGA6s7bTqLoGMfQoGbw5H6rHAgAisGes/hYh1Fh7kORBphMj7BK/
PCdq3z+z42Cf+1z5r4vUoC+77QdrP1YZ19xE8JCHZZ2lJwqeD+0ca8GSiwp+VBKX+h6AbJIUy+l4
YMRm89otuuZzUKaY7npeEbEdqS0VO4fY2HkcU0yzHC49RIsTU5eGXHCB7h0TzJgHg/eW/3AbBPDU
KdllKd8bzYjRXB7PUuQdWZHRCKzXDaeOQNJFvABjcikBewRHFXXY8vaKZybmrYuPLfWpHUZJCv3o
cj/1oK54V0rQuS1H9Wc6TrNrkNEvkJKRxkvPzlHy2teWkFpuhWcSEVtBtth/5nDCUTA9iC8S3akk
/KNHVE2Fxj2VygtY4Oc6LkHWCKKByDzflhRRvKeem9CbM6wt34SsgKv/qEu9ZZmWMgzB9ONK3f4x
TQ2LjpDY9r6dkSN2ueKTPTNc8cZKKoN5tMoCzr/YV0d0Ys34uLTQEfIt4IS9A63cCKPwgdC08bzL
9Gl7U3syqSeFT1EgXW7ZMcWSTEnXE/b52D1zlbvYkjvRERV2HyWXYzc8RHNjvmSQWLSrr6NAOiDu
cinH1dPbsWMQQvLaftxuBdH1x62e/+i5JU+h9uKTKdEHSf3XqRjhSH09ArHIQ+WmEil9J0TpaLUh
QgxcFbc3dho8pBeh9T6n+VXaSlqDnEiwALt9s71KQFJlbsb78V4fqFfVc8sMR0Y1bn63q4G459xW
X8bA5xB1FmfyEKCptMz5AUS1I7Jy3Q/nkUoo8dvlDlH1oLF/MRqPlLbfUw+GHjP+Fp5pityZTneR
/7V6I/FEGhf46YSdDRBSWxe3+0ij7LO1+f63XbXADwr00126KJMYyINef3IHmDdEUjVkDpvL9qGI
EPFta6CF72Qf96E/MbnQg3Bu/F/TEcfOR7kvRb1kgcygojICcQ1joE8lvQekjimO3rwpQTen2C37
AUTqn5o7Ck03VdBfEUxYXE0wO/yH8eHQpB+F96B1+3OkD1Fl+zXB1BORHCSqPTlG5LSQdW+Iv4Lh
aL02k0kfyYgIpQXDVVePPFvjdIufWVgSlfbtvJmz3PqCgP+AkJ2vb6Tgg4GT/0Jo59NWTfsYRL6V
BfxAqjR0RjcTRvBnz1WyKWY/ZV342fDTAtxKXuKUUBtUgRy+JcdSsidzMCTHI2GEncXOp0NpbXVv
FqnZlPGTjfGBxRpIROTezvzgSQS7se+mtMnLbSuxOfT4F+7GE/OzXfOB0N2JWa0SOSqT7J2vCVM5
Z54wq+0oOMecQbdYUZHcQFvvbJxMgOhr0Rd6QFP6eCDeCShjSvJbka/1r7CExVnW+VNsoFgDBXn3
BkQ7UA8V9DLijFdt+aQQsNS8B5Imz5arB8IKap2hcsalSnM9U9Wdulo6b/VNeD4jx4BwHqI5r27I
7sI+xNfGgPB4JD66uGvq5ceshCJvp+Y7yCWeyP1+Ff6lb5p3enHZdfZYS9Sm0nkixxgaOGk4NWE2
sz1HkxT2OGBGHqRrQA/cjCVbVylz1sDO/JllAvrdUjfAnm9wyG5gqZYZ+Gpy/umqu18Yc8m6LGdM
v6jWjKisk+CSdCxONtrdxoAu28ADs8sVnDK7qyC4gN94hbrn+sRzMrbUX2IeIW7hrBsD4JNwkjit
3sCVFV6bL3lFpXar7WQWWv/PBDL9A5osKwAELjTBGDavNSMKlVKfjoPYjWEoDny7IOhtiOBz+QEA
xBYVnRmQypxU4hBO6hTfIo6uEWT3hjbIxgXy/QObhKrrRnTRGQ+9G16W14St7dy9kCLobo3Ipld/
Jb0uOzpZXUCbEhQImuUk8OkJNPQoPE//WM5H3bbXOPqTXsYCpUDySjNviwKTIfnlDbR/QTpF7J68
CmjOphwaU55WPFbz33CJhV+yDY0ADaNTs+94dFdWxjLvn4JwSKGiTe9nL+r7rrCyXzicmRO6+c+M
pKrOduy0hmR9AHB0r6Fe8bJtkgTC2aIG9JAxevQarFubORRrMOyDY2XO1SbfxmfaZqtSuYWx+T+c
UlIQwQPqhFV6TnthVlM4WboGNCPc7vcJfQIohVkMBTU/BJhDY+wGVLk5xMci/We1sy+TFwC9n196
q8kjE6fj5XnYaIMdiBkfySrZCwKit7/vWau+EnhSfSppKWlSsod79uXXXa69/ZE+Uj2GDmnSfbEM
lqEfQTgnRPKdjukIYHy0ccYDSR3OgSIh+SrQKLOE1vdplM7at02+0gwK2T5URyR9DokSL6ke7Acv
DJmk+LrCWRQavGm7iSeK06OyRPeq02Ej/wAPzhNV4OqVLdQj1t4inLJb/29yz7XTnb54ZKaxogvt
RhHyqyKkfkSnnk/waxkmCwGtI2+5PeWGNgLC8jgcTmf/YgfsEbEW4QQfeLuu1BiWdN7usHqO9PLB
6fVK30ROkIpxPAYJn+X/T1T9iM283mDuWlZZwsgXJusuaoapH5lC6Nz5Naa2izxert7DjA3H8N9M
tRkg2qfvydVdwK7i2/Nu/EdaXtHyZfJCCVZKIKR1hn6D3veCPb9o7qWzwCru0mV5oyYfbYgxY78z
AxyDq8n8r/YGtq60Mh9qC65cC9xAdQDyjJbX4mqIHZ8hBW/Q1vxxCV5r9mF57N+KzTg0XqVeR7gs
Cx9XyHz/yrS2CDo7M3TjIcyPZtv11Ct5O7UZnYHADJlOEtwuYonmLDdzAu1zQjaeAgtxUwiRbYu+
dwa51vUOMxhOZhKURud+pck77j526AOrdT3D3ihJS0kzSOtosoDH/ygSi/XxlbrI1c9zxiupmey0
IbF0nOz/rVJpZfenui6aF4khW1ru6/4FOuF+qHkjLgE46Zw2+v5EyDRFRKn71oMiGVE3p3Q6ugwc
5oaRESRVNGqA8mpvAKkFvw7/rYIuZoJLTdShPTyLclzUce4rAPx5zHUxw9TjovIAYdzekls88TWj
21OIAKy+i/BMSsI1q+JPNgYGrIUd+FyolToweVMcfPLEZBMgyXS/293pbG7+6pCjH3dxM5mAHSTR
xPKZK+hcZlEupwY3rP7ASWkpmcr4JDhJvpizV6LnQI3UCCkuNAkXslAYBW/Mix7oGG1uEn88AGcQ
T6I1SX0kB/JTDm9kEKGJqmMRlgzA/w1E2ImKdnOhBpV0qdKuBDq+95aVosXiDJt5lD2HEqmFqwJf
qcPt89sF3egLg1lKbOeirNSURhRqGThpD3yLz5qi6Hhx+TB83vRz4/hqQ57QBT3szJilgTdu8PYu
WP5YuOiVlUe7y/ZlV/WJyXX9MzZLhXNaN1U90cD491u8k9n/jEpMR4Lbl8HB/cKdIm8xAFpPcMaR
AfMnxHdE97RvEwH38OHuPCoEBtarjSxWVxdQul3iECpszUBhovBbw4cI8bUG9EATUR5xlPlvshXn
qW7X/VRmbMSJQszKEV7WU85Bv5V2BwF6EKMeVkDOO9ozS3uVtBxQyProI+KYTIokZxSE7zOO/2Oq
6KrlXW/ZTzUPLELFtjeYf+xLWT+DFNx3s+lK0BV+/8zOjDPFB+/c7aSmLge+x6fAKZeZnkUiXTuy
43nbbj7fN12skuD8a9IqLvgR+KU59s5Km/BUpN7ZhSdgYcsbd3WpJuXrd8uNElaJlTEoPxxWlEPW
kV7DUQMPp2qcn7qXfWqUv8elyd7i3XToOzNhmPyiD6blMiWl5ZY0Ye9QqUfLvQMESx9IbR2Sdw2G
j0WekR9YnT3lMW3KvO2oqjx6CUGQ8/OzVkAyzJQ2ZRQIiykWpRJZaNuNtZzvWBe/k/XnBKpBNZbG
4DNboxY+weCYYpdXpXNmV5lkGSdwQ6h7VrpHJAPFW2lJVAXPB825FKS1los6I2sebXw0k8ZwNLfL
FMu6stESjwoyGj6GPgWTcZfUnRI+QQButAerPHV99NsKpV/qy4Q2t2ZMBhdzNfgUAvJp3L1WTfNj
SBkBjgYlc2uLxCUdriARpnmMjhUpWYSBW33mOpWeul5U6DDFzPRAXexEOvYw87NrCg9rpJ09wDmZ
k+pYxV2kmt1yOEbq2lsjcchx2qJDkSZ9ai+FqXZ6DX3MIqOgznlIznkQKmrQDhX5nFKgoSFfXw6Y
CuaVEzX+gFmwjWv24ZOoCKRzWFmcrBxK/WeDmjICzsaNySpvoFPGErAd0W7NvXMcd94jN+Gndq15
IGASgtsfKDeV8TCpVB817vcdUhdnPqZhEFD/6FZwZPzq7vuiRCWB5D+XzCJ3RtUhPro89az+q5aA
6R44IFn6AbTwrfhYlQ9gHWTM/n3jKx5hQhxGgtS7ZyQy+JPfPbW6nMCU8TWux0Tp0ti26DIxVKkc
AT1Z+E+8JRb/cI67GiMNnP3ZQsV9AF/p759XTqQqVJ86NJ9iX77PpP0T5llVxoARWdbw/i6iSFrn
NyjOE6hsB3wycpoQfW5D+C5NIPdaMAhb/YmGu6PY5bbUtZWBez6dH3ZqXUilW8g4JUi+h+/3Tvrv
1oxgQaPLK4ZrNUicMs/5Pzc2JUVJ6PAdbUsCpVkNDnXhbBXlalqG+cggmNSc9R8IIM1CkcxlStzh
PyTKqh2NwSVHYiFj5xlhbsiSTDD/YUVGeHOzhRlYXF7QjDsSl9dJHw26a+UlIw0tP/XF2XL99LQF
ULPdkDT84c+2j7+gkOcAu1nm6ZkKzRkBtmLwkVypPvsVdHn7hh2GWkDY57ZINPMedOlpJAd/OJxD
OKENBIcyZTDbcgrS31xPtgEMoLy9dlof9PZPwQ4KDRvieeAb2PsHFjL803LZZc4be2MemREwn3ja
bg7UNke8eFcH2dYHBaQrg35/XVwjhJ+BzkF5/KaXgTEuzI22VGS3aVeZvqAfZdCbkBzy019aMsGz
qFGmrMH38sQUli3PJUrQv73ZzuoFmV8IuwFhqhz5iguBw3eB6wm0xD7F05KIu2aDQxKldBglFqWd
3Vn8YXOinRQ2dXC954wqx4dBXPWzDk/HqBzC3vyd6Yib/aSkkmasFq6tYr5HzN42yv9u+SjJ41RY
ZZxwsGjrFCp4rSgjM/K0eTjkclqvDVCcRmw9PfIE6Qe5znMH53Mnogse363+PH1mzip0VRM+KHfv
4Ea9xAVCWbVS8YQ4piNNue0G26HpuEaFhE/XmuDShRNPd1K3nIFX/8kO8vlXZSxZXZveopyTHF7+
aJbluEWFp5cUsrKGTBKMRMba2nhdbuPZokXYsCRpiRELa8VaB4HNqbdtCw2yE9xmluonYXOzs7AV
TATtxcdgkcD1HB29Y48ZiTGiCHat6oy0bteoS+3llZS/Tdcsoy0vC+MQyxKK+9T27eOSEDvIv0Di
PNwqw3ewXvl9v0QBcM0v0nBZiFs1acXU2AvPDln4PhsMyQs3kocL2LHGnG9v7BKQoiRK4yWMtFNq
JT9WkobZM24QGdAUy4uLcKsYHsNOjIEfBQTfsnLirJOm4r53O7MjTLj3ehinDUaqNWlyju6J/v45
0+GA9CdQw9CEldZfFJwpss6e/W0eGNC0JrUR2giJDYxM8NtgD/T2N0qNX6xuBZ8CcSMj0q38kxv9
czSXlP7chm/xBJAqSVDuLZSIxXaC1HKg92oAiB64z2u00TWokbHobGIEVvlyhbGUK0lGHHHK0Qfx
g+ve65QyxCSZPT6klyaV/NatqrMFVhGMrpbiTrirHu4TnGFJkskrh6AONlmnugpPIkhyZFPxa89i
Wl+HjYTKxUZf7N4jpBxy+1BI3FqWXDOQfFT1Sc5ERuFDOnZJltQzI0LuodpZsojLrujNpp5txDyQ
TVzzVWkwmcl66IcyP7rSGdQ7KxewGg6oGs5ntZ1ZS9GGFxwWRZrqcndMw647PpOP8BbJVx3r0w2e
Dyyb0ER0squCm+A3SROhFTWEVQWAUlPvsw355NKIAIk0nPeQnGGqQnRpDl2QrqfZengaugzCoDzH
rBDN94Vk9RNxfpfySTLN1Ibi5dfin0wbNO6DjHa+oTTMDyUeNGXphSuFYJgZTRwPzD327w1QGdRg
Aab7x6jXqR3wy1d1H42W47osTgZcQLJ/X1mOZ47Uh7VGV71u8Rr+0WHZuVPnNYwlkwWazEDPNAv2
MCNPBLOGJgh8D3nV9q4YbytQmYfSk1hScI9kbs9S3fQhDERkSY0kDhpohfUFg+YtsjHoqkrI+doF
H5hrwHnVgALmiwLnNPU74n0Eu+WS5rw4vCg63GO6ovIkJXNHgRY1Isis+PuLGnZVvoR3f/W0KjUa
+KnYIUWsRcsd4r2Io0kw+/7pC5XjsSGR43ZKlovYDy8ZOnMvhpnhPuaQSEEd12Ma+O6/89iBil6L
+beihjBytBIibTKFgEzYfEmGgr76RHUP0IdVDCiUbNkugJ80iX2LnaixwRprypB9MRziNmzRX67D
fAXw8QzeTuQv10j2oeD5s9IhEEltcW1cGQg3pqaIJ9LIrNTrmVOAc9vS/Y7n+dTwyoXnMGZfQ57W
BYy3KhCfWYKqw9ICgnDltFh6geeFHTtP5Oat0ODPXxkjeyHvLXDHeegEu08lcuWVMiF8vo9a60r1
LJLXT5JcsZArZVZnRhx8/a+CWn5HCs0+t0MIxyqQUvbLfUjAOhhsqI2VtCoeQoXa0EwLSFNmL5d4
BAbdZ0PhfgIYZorSZ6d2YLLFsCXFz4ZSPLgpmp9C7Ka1ZVZtxnrrubrPE/YsRs5OfaDMDl/rkq6C
zLMt0vl0nPS0Ych1Zfwg7/AhRmPqCfRnEH/j/EFPfe4XOOJjtyb/g+++TIfK8qXuscd1W/VDzsQF
LC97dVJZVoQdSFygwso4SbLpQvamLx5+XUNY9lA9ZNM5tqL0Tm2qY6PTske9yrrtP/gAYnCxpW6m
w/jEOHYBsCl+v6JD9ZMC9aqRSTgWyj4Kk867HJfmow9FerSaI81BODFleA8jSxrXKe8CqJZgx/J0
OIST/54Y07I9ePNLUwDs2oE1n3NW5f8yGjkndTgaR84EZ4LxWzjFBKkf0MycQv9hkZ6wqoymvTgw
IwYUUyD8D0klq9JdDSN0c2Ts45c/IWfDvM//X/5K9lqE/daFQc4JL+DyQAkd6Pk3rSYhXDQggcGP
u1yoMsJ+QwWEFqw8vtxzYITspbPh8bsUXEQL0jFt3ranfJfOggmjuIZKjghTW1W5rz7MU47XYXHD
vgyQYV11Lta1CMSc8xWmC9Tn13EDfXU4kJf8PtMKwSOnbaJ3OqWotyphve/UWBn+Mla9qpe32dM5
YdkbL38Aw6gDtIDnVP6n8Is4PqLEUI1Ln3u1JNrtyq9RtZCmU1ERt2cUKArPPnoONo2+v2G62U9e
GLflubqqntoE46AUnZTi+2Zktsyf3t18sTvViFgQQKKYSZrpEo38V/OwLsG67fq0Wjsb9mJCNBlz
NyFp0pvWcWg2O/K2xT6fG7Y9YcdQ40DUltjCMzOWhv12AM07yn1eegIk0h1q/z8HxWW8fPmi6Mzq
8tT9neG0Lm6Wjq2OaN/XMxr6ziF3Knce5V4riF83jmn9vCilNkRyeoWdbgQkj7sD6oXRS26YDoI5
d/qSx3uT3Bx/dY5PnHNHJB559RFCzNqKGeG3j9Gh4Laj0Le+DMQ54JrfPUpqF/gaAn6X73uqnNXb
WnMh4L4My4ORG5m1w8eQH11q+j4TGUx1WnIAlr9lDDreI0x5BOE3e0w6u4SxIN3/avMN+9C4ItmS
LzpY6xDdLocInBUjsA5Z7fJ2h0NAsivN8OEO5r4N/7qRxEfoxy8QR79IPxS9h/EfuCUGXrXV/ZaQ
/GhXKrbnDSO/wa+kAe2dIMqOflcGSxxCXkZjC9Chkd4WIfSbRuoFZT2RR99LxNKQZNi+ocXBerU8
6Df8Foue5fYmMK8yR86TTXBItHJkSjeiMBYTV7gAld8B5EAT6gDeGrCv09tE5+a6MpWUSVWGIcjI
jaFFtzW13av7bADs+u0mKmNz4LaMoEWsZWf3wzOwBwOZV6d7yhVHV2iZKJ1tSUna2WhLYJwFdBgO
6RmkY7g4vJpSeDWALj9oXxoi+g1VhqjEq1crPzFERgm75H8A/ZRHwLuM3vvNGkuOKiI1hGHfnGw5
dej+VKHIkcqwjoRyKwh2JUC9wEgO5rG18JcyeggOwCeytSg8lUQBmh+NpoHuYGN+T/W3A5eaN2HM
MOv0HssTmem9y9abOw9jk5a6cnQiEYosXa2EnzaC3heumInbL6dcAIzit7YrJYif8fWhH3utEsN5
CrLCcYk7dX2FDNo/DOTDFJvXR1FX++MNJRL/m9UITnQiOaKiZW2DEw7Jutzuu2kZ1MWRPnZM20M/
PL+/mlqYh8bo1g+H3mgzJdI4jTO248uOFEKsOD9ON/kdc0tCzUDNnQKI6sg3atm+tJey5T1y/3Pv
RHN576M1LdHd2R7OWe+jfhiUi1XGZQQ4ZxvjCJjdxMR1HocGQ52imo/BPKW9b4YOufZVjWJB5vvp
WgH8kekmiyiSX2Na4Rkb5gCWiCHEn2jXWnrOxbuOIr1VrrtAL6vPHVZpc6Y1i37eG/7uWolEaHOG
j3YTmyeQtkkPP73GDonitqA3O8nlA/cahNnXw+jQ0MPVpUyHnlD8cqiVBdmOUTQ5WEZ5sTHw8SW7
BVKhbHWGXDwmkD2MffMCw+Yhhmj6g2U/p241YeOxuyOgZ8HywEif3NGTyq1YNgoxVCXOnzvTkrRs
Pft8k83snxshiT/96MvE6PSvH0qImCDZXlDDAjvW5CtLXuB0iniPJ45fRyyi6KZWDKMo4omH87ty
bDnJkR3F3JvI0QX6rJ/WbdLJp0mycT3NQRo7EQs/hOfHztpyCVtZhYbkmHMoewwn7hiG5a45OoNn
ZsyEzDqpJ4YMInW7/EBw2G9kUKuQdEwU/GZD3TmbhfKJoH7lJjfdfuyM0DgWzYyxWSs7yaWZLXIi
bCMACcqEm4OFHz2En49++uOpswTqx/iTPtH1OAG9SI+b1hjZVRfGKiVcY43N5l+G4YNbpaqfJUGE
kkX0iA4lqJq1woJgpJnnOWU6Aoj4GJtdhGorqIltS08LTqIjgCLozn8JntB5O80xNsFAQEj0RvRR
v+eHqNRbcnvv3EIN7S3/EGDSRNzpeMgc+kY+bS+iS57IZZRChS1P4zv4ACwLqe9Sw+gW+IK7GpnD
V7EUSi1A64RsGSb7V9qbxQLDsWUNI7Js4ZaqJcjV46MNL+MNGIXqCAoRg1Tha/2s2tVLovVv0ffx
YQaheFZCn5ONpmaG3jHDSV84HwxLWxUAsBKOCaJS4Tg338EMeFg01zpZoH6jRIB/H+VEffJ1H3jx
StPvCpQSlbD4Y96psY0e2OA6KAOM45TwzGNw+XNASBT6MbwkMh1gAYxCiFfkV+kqWHEEIIB5/ej2
P95P6t8KdnQ8YLM1IhjuRlH9oDQmA5l7gHdnQ+P/7VVxf2PTT2g+rUVDYCOer4+kW4rxc/h6ZD7r
dveYnKESq7w1Q8iQLCxxhDujj70YB3cm4sWDucosuHHjlx1O1T/+R2am4Yhktgz/q+rGQd2XMYVC
pqHmf7gKDnEdAIXDGTfH5dK6BBisJYL38pjVZbbSpVEK0uUZtSHrNCGYfiUYZDlBWftDB8PeKh6n
kRFkHtfEL2I6r7VKISJcS0my87lzgcZWQ7jQe0WdU7XusuWR8MBytxTc9qrRkgm6yakTXl6bYazN
80aRRV7tUbAf9i9O9QREJq0e4xOUJUvYLSSLmzCDrdQysJ4vOka6u4O8MaxSmCeC2g2sgonfqd2w
4zbMVgGVP1ur0ELh49Te2o2h3w8cmJj6vHjyvDOw1s+OfE4PbbJw9qLXEHi9Oyn/OX4Hxw3jBsmc
xwq4Lv6omMYIQHv9RL5GOBjBdaqLFC4Nva1s2PpGil65PAkKQs4AfMrdAVDUNg/KItXSRNYNhHGs
OYe/n8gJVHyJBxQivsmpogIT0WwQvrcK1+Fl2YC4m2N++jHoi2J8AZTD5rk05gtv8UGKDoukR+ca
cX2RjrIjZnd4avLCWsnMMA2QlP0sa8eB0wdcn8yLXtzDJZSCHW4PZcTu528FN01f8Crkz3XsUpp9
LXOK+zAUYTN6DWP3Bweoo2kKE7AMG6CcIvgNFU4BIo806CLkh0JGtN9Vr63iGw/6/mW6VzX2xXNe
pFZAAIdcjTTekg3aEkI1g3lwc9717SeVDEEh4+h7bJY/uwB5Xnx4fjJpxERBjTu+0ydUMbXnyDKy
fNU6ixE1J6QdGjplkrdeQ3qJcI9iKjhnwvljuX64Sy2jo36Q3Gb+roDodRLIcScQrATPSxHMBQtc
5/ufshBBXczczLZsOKyTS3tfqNoMI4IZ9vBtb/bl1tLScJ+mYl2K9YlavUWSUX2kKKeNweyWyk+5
idLmxc2vWCjxbtkPas+wE5WanUxsKQCeFTZ3OyQ4oQzPuWCeCP3Bl0Z8eYk89Vf9/QDECug49IKQ
bKTx0Cg7/kOtfulRSuZ6PnLhClGGkoGtauPdb6bxXlkGT1cE+uVM1VuGE9cg9lTpXt8NQC2B7nRH
Df3tXYxnl0tHpAa+SgEcb//5FA7Ks71qIvC3QybttXrm1+TzXPq8vFDQRL5HYX/4E7tdEJOJz+8Z
FtERS6tcClKONMPtlUlFyQq7m8zCv6t+a73QGMF6zabjA45xawGIWRSudTOt7pQ7C52N6BBQiKuY
OYfX/FD/UOJ2dxuR/3TfmQxDHFUXoYNBmpkdbiQeTL4UoGBqChUkyyghffIztYqCvV2584J3aob1
zMco//sYtk1VVzOkAKZcHgGeAktmb4CiAz6gRfKopdTMFoG5ns4E29yafgXLoyGN/QLfLY/RX4WT
ZJkIdp/SNd2AF5DBLWlpRJlOGqcey86zb60++e0aZRxQzvGY4M3W/RtDlzXXrmxRQ2Vz0YkYPU2K
Oh7oyyKIKFKDkGa6SyRUuKIBMokkSYnjZ8exMou7+9tJ+D7rn9jc/27TsFNr3EiZabA2oQdWA348
LAqm3wBRRGV4BGOcxXysblPMW0qA+32rKvZoXaLbCBbJJ2jJzqkS1sAtRLJ7L+Xw+IA8pVZKxyk2
11md5v1s2A9wlidCGPRI0g20JJ/8Jm5YOhimmT7W62bvvoAEEDidNq8RvHdwCfvdoAuEa7RXNj96
Kmm4sfu1vQTmJKznrvTnkBuvJ5s5bg/XIJpLVk82lCC+xZV/e6Cq0X9A0Zv4SrOhcaXDNZEeK1qv
V6QFSAUvwCCkbOeeF5QXUATOSAF/cZHYrLs+f/XAmYguPAYsqfoNu7o6r43MQOhLveIOSIgjo9Ip
TmOAweA+l88N3+YDEBZ4JMKCt8ps1P2GhGHSALfmcQ3WgMM+k19LaA9eYf0rhfqS+3owBatSQp1q
TBFfvgD54ORinDxHPudgXpKpqwNwvZWVqbk2wzjjKsNqlzZdsGumJqMn4vpF+2J1FkbMT6nCuQxd
TelHnnVrzrnenuXQjdsyTeCcY+mnMs2u+czFV1ArwHzOXAhG3vyXhu49UeGj9mBgWC0ID4AXkBLm
YVshl+2hMa4/Vfn0znjN7Aapf85SI+OcGbmjx4BqlEyAgUpgRfqK/yNqVw96M7WH+GKFjcmkpoQd
Uky6ILhpKwjILfQZtIne0niJhf55I3gbuHEfIfqdF262zZVMFMtqqTWXleg7s5GR3FHuoyEgJAin
yvvAAMXXKZQIdMo7IilCTqzbPHWXFkrJK78Zw1tXtvOT7s56s4rUl5A2iDisLvRhfy1TMX5lklrZ
gic36H86ZKF318EBQPaOJB+ZPhMjRU0qH5BD9ZHaSFtPtZEqn1OfVMaCqtv6dw8Sg32dVNjHFaGM
BYM+7N+Ci/dJecZQtA5dI2MfA/AdokCjHOh8J4dgS7SbxTPfwr7G3f9PLBYFsViGDzI/zdKMfXgs
h4J0fZX0WN+GbWYXxAk6R1peYpRRiojlFSn+k2w9u3CL6LfjfgIB5vEtYB6k8zjg7stHj1/ADs9T
lWZB0IB4F7KRwczq8z+01LTC65D64bQEPjJhrSTABjV0Aj8j6zKtiYDbezyFNIjyLgstF8QScaNa
Lk8biibC/AYvINvxxK1OF/aJL9BFy830QZ4V1YqBGu6DsphpJlB+otppWYbBKQ9mDwBnq5tOWTk/
Ia9uhrbfT5Ij3HpxG48+spUMd3n5+gO4O+acMhjj3TjNPTKerDlwTj7pWuByUiSwYNJoYDOfrm20
QecDmo7HNU7jUIhFeOYLFN0uLxYERqwsdRlwvnKFdIYb1qsA+pX+6epMZEuYVZooIyz5iMQLhBxW
Eiv2oiZFqehxCb076e4sizzC2qmaT00nDItQkXSwrRMucJTo+9Fw2kG7ZhDSt5X2rrIi2zQx9QvL
gkUtUkNKtty2s6r7crYyUlSNPzlR28gEMT/sfdXiCAF/HuHV0SPdxNXQJcQf+BGa6xbNhXRzy8TL
Oofv8fz1qJGV046xNJVg3winOwCo9zITelA/o0WyRW48lL5/7DWEchyEjYQ++ha79lk0m9VfHjLz
PBpY0tfhUm27Bb3X/BVrgMquo5chLnrV0Kc7cgWsxqwsI80CljA4Tn7BtATuCkWMu2WQ+lVPlq6P
NG17GpEH2uOCd71Ee+Lt9bfNC2X+KXsn/kCw3vRoYsE7IcsfdJWh36QnVz0BmGgZrc+Inqo6JdLg
V+t2UmpKm33QYykr8hOtYytrxZAKcEAd72rDCTXgbWzU3Z5Hdiwi3tedN/hv/bbzlUAXkei3NfXn
6GSZZJssQPLoWhts0oyb1YoqXiRO70bWMAWxTPw9szbDOocWrLJAmpzVlHHd/EpApGgoOh8IKdKk
Zi7cgKpuVMoWtfyXofL4OdcXkoszdB2fkJF97ZL0/5/bRtTZjyM06R8oRFNC6t2D2YT/O4NUTado
zmmelgXlRBR4IG+T8OKmddprTLHdOo9wLbt3N2PfU1qWjlCqc+LI2Eu8q9ViH3v7gyPYbS5eDfn0
xXXJf2b8RKbALqDCbou8EqGqCBySJtNPpCqjeynbq1c6To8xGhIVbXTGWIIKmDkhHI45H/Ug9APU
/q2nB5MsZtZwWphkW6Be/yTCzpehm3pxRaicFfcA0e8ZxDqiSIaH7O2z4fB8SrQI1dBs3yjta7Py
oZibtT/dIwFm/WsqB9kE3IF/G0LVv0v74KKuJo4j3efCLMMkjXqMjIermT3K7NFHypAQEJXYhpgZ
1of0jEbWqBLD2/UnWblXjg1GycvfIokxbtYSO4FyfJTmQgL+d28uBxrKYNp+iDIQ38Ln+n/PNWi8
8qhXI1XO9wTKqDOHdHk6VmBJsOe/rzqNwMLp3bkBqwyYCMY4/sJSWBKZwgsX/EAG5Y1sYDM/yIFH
XukV2qOd/F9Gv9+dU2c9IKceKqt4zXl1vaTF4Sydb7Lqcq00LAeKwgBzfYVc0HXN8bAzFYNh5O6q
YgU28DIMM8GjI7CsDwpANMpuVCcW3a/2G9Tz7LQuIl9pCDjGlUnWxV4a1Ujiexf5xCKSZSsptJK/
ZBKDy5EDxNuB92mUcA2gSJ41o3zgtni/tH2Z87R0wAwmMkJJItK6TyXEZz7Nw0iR38gNc/MA97NY
zAc8lrIsWg95CEp0aDx/xhFR60RppvrYc7w5mEZ1kpLRE9NfaevMOipM2x/Z20VKu0Yi+bgVuuMS
IPIEnbYW/rKd7hKkCGJN7rTzKieK7BdOuZ01B30/aNxaFdpTTuY784qLsLSmXp975Lzfb34DEmsS
el24W7j8DdwVzd3ZQzv9Jx8VA9Vvcmwls2o8xpPiWS7CnNqz5l0Yck/T9pkldRV/Tt10CV1sGtY7
BE3QzmmKfaY5dIwMIO6El2tVJKpjWHURhoBIAFcoesOmhKTb/f8Nqmm8S7V5aHPwe682ggVYR2xn
plYB4k8LJKjY2hunyNVSm+nnn0lTgRxEzMEL9vyxH8ALHpJLJePxORg393UwCqpRsi+zuRV23MB3
yFajXBi6+jVwN3kRo79U4UBR/pPDygjw6EtSrEvbl/cPb1P7gp5mrqaCtgm74aY3wSymrPfHi6Dn
kuFdXtAjtmO4hIHmfYTKjTarQDu7RacksQd6342VZcFSJgTfg8rRf6FVRAxMZ7Z+kWGMLbCRyUp7
tdJv7zR2XGFhLOaomG5QKXFFk6Ezad3xvRc4EZn/zJ5uVZbmllHD6jcxjY3XradJDbwvsCU+yzkw
ElWae7qmXKjMiX7E7bKnvB8c8zwApW4HgPzuKDf5uEVgCu3rI1rV33AijKbk4PFhb8/R5SICoza6
AHdd4VX51qSJV18cepAwS6pRkLywd7VVxo8wRBWWmJZK1Qb0GFB34oy5eJ8z3OgoGrT+IZionUBO
A2D9a890gvko3rHNHYZnfGajEEYr+ycI2fQEaTYcizTlqvGhwuI2FMHpWar4o7V591dMvDoBcmqK
g9rjZf9NHxOm3B/KChWTRoLmvVKSZHL42joZlMU7YqdVJ77RQ8GoqnQ0hJcBsojvG1jy9Mdiv+UH
WoGs4eeEKNsTPLI3izOdRjrGPfzqm16LzsXvHeBOWWMM+mmdy0AO/Y8sGhiqX1HEdg4XFKCGsVSe
nZWqmR9rSKDuiqgSVisWnPP/yJT/54dYKz3zlTkLuaaO7oJwvbgoYBMUGqwmgnh2X9II/xGHDSKO
nbMTffQPQ6b/fNvTfC4T8e0yc9ZNhXxo5M5vhE8uQAcr8oDJLWFT3UNuZhNl1O64kX24WVqmoRp8
qRB7gkPdtmnupx4Z5OKWZKKqM7VSSXFu55TVo1pb2gTz2GvTVWkdXCTyaOyslRxQ0vMdgCDcKWQb
fnIKrhcO8Sl3gOAR0IdUkxU2X5TdUQtVm+9gKgszuzBGzdoav+Z8rlVybzkaPO1XRyjsvCM0400S
a/dJvH3RdZ8tSlH+HpGfocBltgekZRI5fcIjXjSF34c98iUSJ9dZxtvXUTIUp0DRdySQPUXMzcOB
tRsiDlddBPEOtw+yh1L7uv0JMwnWDUnlpgQQKwIkPeG+WJ7kRPNHq44vmrIYtgqBjFYu3Aj54gSj
9hT/0+hKRURbcsnQoZu68G69FRcLIasAXpiXHyreKkimkwjFoSgKX8pjijxStjqgRmr0E7+2nE05
qh+PEnJdTkNKHQUNlVdzZwOkNoI57pmCCrapibkpiiQ0WP0/PaNqpkj4+w4vXISiQxCXCqx9mdZU
cWLY40BMwl/qSaIFgJaX5WTIqD5H21AY2J7sMNFBv/2cpRoKTxEy1hkdDFkFckJD7yTWkWGZkOec
wa5VAEgIepK3hWjPU45FOvgw5rZRYw+ay4H/T6QLuE6/KePIplbl46lO+70IZAT31OQw+SiSluLz
wbPLs4gVuOdbREL6CylGUWkFvInA2L64JzZ5gqmFuiCBImOkdOkESrXyNt6YoOqEJ60UcDIe14Sc
ha42EDKu0wyPNeZLLsVu7Khv6hP0EEp2TUhRaOfLGFunVDxBwJAEe73jicGOCYgH99u/RIEzk1/t
HbEatCOw8KLk2IwJXZ1IGeu+S9RxME9pFPcUUoOj7Yl0QMBgaj/tjzMSqgDxJPbjc4kCE4/Eu/8a
9qqUNZ9U2OYii6BiSCPU2KZegsoqgsf7QidUM5fJZgKQwOcwLg60SYRif3ZgX6so4UMa8REqoHTh
8g03vpSBOJYKbpJvBtREGAq8Mim1xz3/+F2Lye6s1cyGGJObFWWlzzj08WYehRJg3VjYPi1S1pHt
pBAAvktLp/SskZ/ohUqMgF2jXKroSb6IAx0IaTBLYIANkuo0uQ+UFpEXnB5GhUm2kXl0FrKa/h+u
0TH+4KHO8Pqfp7Vg7eTP/ismEUHlXYKXseGgqcBHE8Zp+DS+DNyrsCH0vG8WPYY+KpxI4wRcUTjx
ftZtdn8s4Z4w/nTSpY12BsUqUTVCOYIqpcCg/49ADhT8EuloFBNzXXzPx8oEm5AAkDMGa9bgAGyj
EbzBO/uBakRYHIVV9gFq2KSTst1XqC2tqdgE8cjHa2ag83ldZxv6GasSAzcFNA9ydTMC02IjgQKe
RGNEJq2YgNA1K93rRXO0O1WLrW+/BJywXddo0Zj0mI3OzSIVGZRCxnmUqphKUXai2qhCXD8wCXEe
qznZ4NHKYkxH9kIFpFrs3mHG0XwyqcH5Ak8I+DWLejMtIucG+HhHSAKzOW8paqL+h97YybVPo9bY
3+uCyKqDnmhcUUnkJrR8hihYLZFAgb5QtzlaxO+txLR62AWc0BB/QNEn9lGvlczjJM4jpVlHlufQ
AbgCdYpyPck6DeS1lOtZNOat1mwph+wC3wmemK/piku3bQqQpVDwU5nbqTjg5xyRKvEYFIsFs7WW
4QpOnrjAo5D8pXkRaWug48nskykMJNGMgkId26KEMOtg4Wg3p8q1aHSj1DolGQRdpnIS6ebmPjwg
B7HexZ5fX4BCUNzRZrJWDdrQYEmJ/wfsY2BHe6q1Ielk+vA5ljgTDWJPkwSoewOKQyZwV0MLCyzo
R1yOenIjucyrCSiu3RwO5CkuH6FdrBDtUYw0X1Ou4x62Hasks4ihSAMVqigEzm5U592JnDYPzW+m
2HuhqG+OBrwrKnncguCnK20ow/P7TWdepZnB2pdLhKuAdHgqAKENPBwXuu2VCsB31ndL0HENmrW+
uKq3P1mUt08KZi1yZ+F/NWtfP8TuGCgQTyOF6ApGsDAEVaTroSqvZZIKysgxXntioWO2sennHSyn
BLWZk/I2uYR+NFhMK5VwAKIeIY4y/BgbllZpnDiVH0oxddzh0AkP4AZ4nl6qd7Skamc8yoZRhqhC
h7W135ze+WPOFeo8XDxeHFdxdJs8TYkbOpCu3BZnmpDaK0JuGEeVjA+NBh8dQvvACKrPR8Xnx7i3
vK6jXPDf+D8xzPYAf/YvoyYuPSCbMUah28htfVAaGEobWL5ZLM62JnOcDwyzjlKYmLWVyZguS+ei
LPWLrm+ySTAjgRQ7W7XuuJDyX7LDUEulozINmeC5jvChLJB1afB/1P+K78apfDoFl/9H8YjbmnvG
kLOrTsd1dq2AqVVc7OFkDSWz3EAcBfjgi0utHcmndP9mQucpg5wDfaIbrFAWO5+uKOmX1s1B6VbD
Pbhub89IGnhONELOoYepfc+0kGF14QYbw9TpC+k+KMJmW0wgCslMPpUIKE60g88pxUSjSCrdybJZ
jW4xXMt2Vb9lPCd6dY7OvmpnT/o17TPzQHCsrVMXcNRqznz6ERUM587bMqcMI2BsWQct9UYH+JYY
oaKwLohkDuXlokW7tq2CdxqJIedaNj+tCIzVDZ+GpCXqVw+FmdX6ExW9Hz2r6ksUXwrssvnidl00
TFiFFo4gsNGRHwx2FVxLzcPACidvGOo58fabI9lClw1VYlA6e78cV+Qqp44pPV8CYN7g0Ir/LmoA
5+PfXSBNGpRnk+bcTIpTQOV1NJpaCFH8jVL/PPIlG6cMg/8+XaFnO4+O+Dsf2kGsqUK7i0Up7l63
dHReJQeLBc2Qfnz7S8g5MjLNNmX8gWSdk/+VPyqv3DRlQ6tthvrzfJrwUBmO1eMGmvEZSrf4gwTW
E3oTpdKvStIHSETpIN+IY7Be3ja3R4695kclPXjmPqP9maLblLj/gHYPZZssK+3llZHfoJxhe5nR
TzvbCiD1fpX6BOD38FMoAy0eJfK5yioS/dN/GGENlHF36EEIYPBwliK/gupr+VasZU0gYv6sNsR3
cDDLx/uqGVnY2cbg7zGcMrYj9Tpl4F04o6xHBUnxcWdtiLhQOTSPnxIOU05flyagN0qwHsOLDbrl
0S6Ls889m+deL8M0SJsxYh9y9ZSQ1PtD57pOuTFVemNOrCuhEYYa//+z4mng0feRyetMqMvGBArN
eV0ZptJAoWKJq1LkPHlZk8LME8xIrarHozCm8fq96N1P9+W4/kpSLyS/odM2W7xtTD4HGyEEp8QP
kchDAuKrEGbXjdKw8KaP1iCJ+EIHQ7AL+9MpZa+mh6R8MAE4YLen5BV1ZMu9j+me15zOToMtSntT
fPdUycK42e6s4EWWXbAOzj8t4TLrk13Acp1O4OWLQmkigjXEeishq9glpsi/4nn7bvr8b4ne5qRe
H9rVWdpiAdj96ZiYsBvR8q9wvhhxl5J8/pSnxslmjgyp0Udj4T/MJdZKCgl8Rf8HrSU7OnadfDND
tMKx0nXw6mk2MWp2iAdC02Ff9pz/pniO9/ZarQ8BhI6hG9A2wGa6a3kiIILzzkjttABKy846bL+/
zhJqcHjqTd1VMGK4df0TVXOqjt/9CnWZMKMp43M8ruL+fRZ/yRowd9Nd7J+WtwD5mvz1v8kDMT4s
TBawLWEr4BMQ/akorgA/3/91AZiPb4d+k1kHnlTFYemqbZ7Qg8yP59ky6asG613YgVWyAL3BdjIt
oKM+wQhR8rWyc2Pmtkn4IJ6Wao1SZnRWEYYMaK0Os7i8HpsdeH2f13DYqnYMSh5v+zNEAFrAHm0g
koWpnJqt8q9Z2fHfLie5mJAiKQLZPi60U+KtP0BYfo99cq9Z4UrfAZ7JpM9d7GMeP+GJAdkszW2j
eSZ4GQ4ENX35zI6hA4VTLvVod2XiS++wLUJ5Oxp7Wi+eGgw5HfIwKHwOV3ue+zlBEBY3/i/LLpY6
yumEtwwTeFZu1csD/OqICwgP90LZgOduPG0xioNZzK8Q58b3E1SvKNvC5XzlgPX5MJVsQFZsz8WU
O21Fbjnjufjsx5xwSn92Nzz4Y9gzLusEWn+XETl1s4vQLoQY+48aL5kVb7KkmlHWbMr8c7gaZj8y
lGefTXH9Nqv05bmUGxY8VBny+VPAGrrj70T3ZUKAtxUFZ8q5EKJ+BiQ1kCkIg/c6EKsOy/yGJVDk
54/yQSEgPbO6S/qxhOt6nXj3VsMgzewwRVsgGypihNUvMthZvzeBYfvEjQHtVXtZ2hFjHhiwOsSK
j20fLP87r78WPEU0+K3tbTUhdQyFAk+82qcObQXlXkdRe02bfcPqZ7UOYiIJBd3tsLOtzzqxNzco
FhZEzLRmOYysMrgYSRLAInjSzRdE9lLpclzq8GSh6x6FguOBGb7Bw7ombPqbTTOh1d9iLLWWX+Xt
oHIRsp/Yp3YhEQK3jezsXq0keMyrZgbG22tS9LthJOLKR/lvpxNma+U+KwnL8UdERxoF6FAvrbRH
uGMhnDh/2AdGMu8AeypqTX0YtobE6RJzutVXGBj3wmXl1GVk5+zP04E1+Vvmr39Po89vBfebIjDm
X05oPTikzI45rl/S3shuz/THscnKIIdbch3Q8cwgu5VjDWjuZtsuVbDgA5LmZyg0+H/46VjKPFZs
DDvLvvFfwi8jQj44UOQa0GPf+iAX5+33HLeZ+sOVOYGM1/IGGA07MZfZBAD1I6hZVx6vZDQhlTBv
MmBYrwIsX4UUWEDorI5Zoehy9w+V2ZYV0RFX4eQ6KGnamtVyJfgzZEwTjKimLOeXS3K45H8Emtc1
pLgL4xKxA6rGcrACM3wNYyyVL6yH76v3FHUzO9H+ei7wQDKL6g0zhCJgsZ6dioSMCxMpeht6yFtp
MI1mmA6pg9utXOQYJRX1xj4LUlmrdu3ML3XsyDiE81pghCepwKGtyBCP2W0uHIreQukU2KAEVFmF
rsfkvDM9Fn12RaZXbrYSuddxgNqansujDmKEcuj/JOI6+rQ3cVSlWejeYdp4hxPhoHBv+AcbUfMB
7xd9mBGNC0BDRrLUoO2P9/qJLG14VrGmwDJNv7W3DNdEbHFsIzxnHOmvA31CNiwq2uFUfpwvnFIC
dpH24OJw3p4MXkumNZ7TuS5DYuqj40tQjpdPDMPYaX9F7vxw2tWPulLRtCtP8iWN4mZwA32GCn04
YWnCsCFF6UxkBSfGGp0RqDDREqeuNDFYvwyuKNUJhueaw+nYgeg6VSMvVqzizbZkXCdPoWl67guq
aZTrXR/9g84T6eUQqYiR1kH+sBGhVShTE/oVL0tyvQOpg4EYPMb1wF+7l12igPvvjQBv/eASXgwG
LgmsQ0j6vZPrbieztUF4EjS+tlCM2lI9CB/udhAUJZXXEH8+T0yIMJktmmsVXfMHwk3cwU4miseE
rE/bXrc34tMPMoVRaT//jTvWHQJn0C84WJoHxsQfjszQ9n1QosHqZFKxc0xOqphQ5Qn80cI1Rekp
nYBjS0n1GZ9l7G+YdeEqHoJ5EDCR90ai8Vp1rBofv4vX+8ojDEwG1ExWSGqjFZaJPoF8U47ieXp/
AmJIaeMETjHC20bIS8lAdIj4oP0axVqV7qv5JEQRU2CRyp3Xur6Jn/Hat8S0gFCs3jLxjJCbsm1c
x8Kbk7uBGOh0XsbQy5zr3xhZWsclh4PEJ74w25z0X/g6kchl6RFf5VeonoCQZcJ8XFdHProbyPJj
QJV3kwFxqGBsxFQDJgU4tLhuP9pq/nMFOuY5YXQ5tCsTiwXvRcCscx4uuyYcgbHc7J+lnBvc9SLx
5bqiDNxLxxyuwcbw372w0XPoaQHVbViqmqHAEztboLl41z+OjM7pEZX5t9gqWaezRej56RPGWZ16
kZDiDvvcnDhSWMF8Axh1qU7+rRhSnlw4014uvw9+Pab+5NTCLmCeLujGEZIXtN7fYkZqra403oQh
qpOh5f76GzitkIVrJZjSiUv8r/Y1eUDJIqWxQcI8UGrcstrRf1W1UM0dVlHONKBakSUXWxX0ycXB
swvlFz2vTmLcBeK86IRKZenh6PeZxR3S7DM9lhuroUdq5UvtSaIsTm7uiz7CtdPAMBcH1r40azzd
Z+iqgDN5zmjZg/cQUJNS8dweOhs81QC+1tgIarNVDnqZ4JKkBBisTBFeJRPKacLjTX8/vQFTnA0H
T5uFdIJgzEwYDuvgxxmYS5wo1PQh7IO0b/x0eZ8Ebbm3cbaxMo+12V87nutmdeGLtx5qcIV3oMv4
kbaEn+0pSP7kf9nKHw1NQBfYGanj0fWwlf6R1RyisAw9xroxtQsXk/QAn17e4gcJC98AyvgwocFx
gj2vF7wLDRXck9VzzRn3FNzvVAkt7tp9G7CUTd/PblXIOK+a6YRN3BMSmhH57onNp6DcVYRqnzz7
3du5G1qh5hH5Y5N/xEGTcqcNGDOUzmaER/hJgucoUr+6uTCJBLey0qHu/yQuthnjSjh/SIWyKJj4
FDDzRP9O3SevWnN/rCspflih4621ZBwH7Qfv63cHJlYSyliC8ufLZshRVGjbetoohrdMvuWQZg8t
MomH/qv/ENizFMNbIT661nKx1nUV3M8GyT2S7VeplkF7DGVL32tO7t4sljURqdIo7WcTl9cwHEO1
AssW1C9AHq0E3X2hjkboQMPmQxiHgNWCqZtG8Mtm9fn8GvYc2Sz1B4sNuZMZvIpuV0Vub0EQlXDM
vjQxF9C2Oh/l4C8Go0MdFDQVXb3eAANa28cNVWJK3qh0gcXH0IwN6xpbUQBQ2ya7GTwQvBJHhaL3
U8NkJflR9MdOT6a2vssnahI2vnBvYv6+xUzSDHkWmbVdKjTS01Fzb+9RaSVyvOC7feRr2cOtfW9V
tA4TmbfhlRbUQAcBQkABPJmtquoCHsZkVrCteBHkgp/7rIsEFf5VSJOZvoNGLcq3ayYmzjWi6X4P
KBtLqHVqK1i1zh6OIKnBZG0m7JZbMyBtTyxVpiMNfsCQWnvSVzTacn9K4p2OACMYJrHriWXwpiEr
NWLPBEgE1mvMw4Jo10BIeQUmKod0iV7LvlsK+6wOAd59AXP/HcMCc+JbakpD8xtlL33OSdJi+Z+Q
hwgULGoW5kmn8rF8G1Qeqdkjq4WigjxglQahkzr7EQfCv8sHuTbM3cu/kiK3EkKsHXwppEMXx2I0
eH4jYjLE7Jfx0NiwAF4OmcLF2Hf5X3A5FDxJDPNExbIUwOyJl6e+UEmw5bW3dpVIw0RnxHlBb+Lr
Y4Oo2HVxVGd9KNp9z4cFs7O66KdCUAmz232JslDe/FFBwpdVYjWL3T9JQl3g4JppLMmQe82OdftY
iginXpjYAo+f2TIOupsN53lx8hNp9pAzGkuZTvpNoCKatkrG3E/j4DfVN9qwd77z5ZZqvLPN28Up
sTPDsI5rChfvYA7QzGxhakkte/330+7wtGCfPMqrdT9Nt4n+VNR4UcTGUI1lMlITYF5bTSrckB4m
jsUzBYggh08jSCrDeiKxgYRV8nyQd+GC/ZqIUrPPYSEC5pbkHgRjslW9rem24ziFpPWVKKQwh0++
nF3kc8n87Ip6TXBimZ2w9JukZB9IrdXYtilN9zi9OULHd/rkiFeQsE8yJK9EAyO5ioJGBsysTL0f
UeyKMy85DX9E4vJrCJSAEVDOByTNvXSus3wa0D8lP/Qg8f/VtuBSoUh09vJjmgvL+41ZzNdgXjO1
kpJgKVPfdYYJsaLHGeDm08pS81b2BfMHiOmdjMe3GebLZXBSODQIVFT+Zr77kNenG6gurcrrXEYp
iYiCGfKupPGnfHo9JL3GIM4Vcqy077dJHHg6MxljYP5ml+jsiUBEb1DvMVQEHrfAEVvXpMelOm12
VuLWClPBXIHICMUW5WHhMnI2nZX2A/9dSXAvsOLtTvD3aXWiqnswB3Gc0uADjH/Z3H6eu8m1oQnk
zvbQKumZIdgtm/9V4z4yR672EBhY0SSaPYkaUZWLt/8IrFSTUByuZjri4WSBeZzBujjP2+oOILug
irCCV4lQwKbNO71m+qCJaBY9ewTPeLqyvsXBbGnliOzbRbf1O+3wRtxRsN60lRC6XChRwDG1kZ5I
YWcBLmimQvUiobUhr9Z3Q/J7UcsNXXdMC5XsiVcp013os0DyVWLsP7ghCWACy1tJuwCA+9VCH4/7
nsCQLV29VIkm0Sq8KjClIzwb07750iU2SqD0aV1qMd0r/eJLmSt5sdC1wMhVQuVCV8JH34XGMkcU
36XCFTwDB255CsuDrM3AGlCvy/rKbf4V0f7FihcYPJGOFJkl/KfvSMu74IdT7JiioFXfRHp0nrpo
QWIb8fer3zZM4C/+cQRCwIrD21xg2WWeysbVI46unnzHINblfQOZ/8HClKubqa7GTU3jGUCxKa/U
yKBBl82EEUUfKNhH+rRt7feCC8r7YuRaFfI1xN7UK6yM9x+sF+mUCaNct7Zo6/2790p1yYmEVk9S
X3feDtFAT5VYC6920QrWk8OfxLnQn8cD+QmA+uBmTipzBii/83qw6IZNKlfNNHzS30uKt+6iNQ9x
3RjxHSJySh01Fjxt0HKPqqDHFlQICYnbepIblckVM0km8Ig6h2mOoDZ/kOP1ZD4e8wu4A0hf8fON
ArwAkOYwGepS8C09Xkcv3jpOTZLKzZYPVvPAbCZuOHsV6phlcNyIZYXi21As2cALTDOevRN2A70y
Mbd6iKfGeqfRfQrr/ocF7ThqqJ2uMY/ctTIbGMbX3mVhEZz5zstPkaxGuaPQTyU/bDrWUJfZ6lNR
I3bpjvv6rYUnmgGgbeF6uTQt7zFoT/OSeM032k9LS+iyJMEhHN0OJ70w0N1taJEnP44EzAOdR44G
pvIeTiAa6uHOVtXZ7ctybWcNhoiRsQ1lUypZUM9/NxVT0ac0uO5XVuUQgcuclGn1kSaZIp/gtWk1
jhNmOPeUnADbnSsIJTcw0sAVm1r6a9LotifyBBn5FBHXMWMM01urocLet7dkH76JFAlTt8ETqpYW
WXDkb7n6Rbu6lqQg0whQs1LqRTF39CQzzuSyfCuP1Y2zFsmuvMGt6tMheFrXKZtCW4c6HVU3L47Y
I7O4De+AcYh9gyRsVqe2gJXE6Dx4k/CzcP48a+RsHIICC7wMYxbbPdU0HAbPGEFDvlQ5k4ETjxp7
LsuzzpbqJWwfjemic2nqj+zAFUVjl8RNaWPSml4xK0f+YLZH8zVc2GzKtS3U89Y0jVqB7UjbY61A
N0dlWWcts2sV2jciC16tTWEAuMNL0R297h34ZaFCPReb8S2vY36xkIlWFsVRm2F8xfC8HC+32nZ0
KjrQDr8zdqiFuRCAi2m+k2DwiPJ+zePitBBELoMv4Pv/6Xg1UsfhbsKcuk9NiBHlWH/O9gqyJLMG
hHE72OVY7gba/PKkcUGymDPSnGBzkjDjCXbgenFPbL66hDqQGtgifIDdDYXF5Cgj9kOgvYj5TCdM
qxRBlS5q41jwBQJZWHmIadCyDFNx1hwMCFYjxB3a0LkqccE2tjKsK8D4coBoyCFkxgSLIJmxpMdd
S90uN8OVFaosHTyLoKq36FIiPQKjctyCKfA15CrHdUk3AwNzA7FVPuLqSeUdkPZB0HnYnIjkyIIM
Mw61RTT673811et3FCsusrik8vRtCl4hLbGoLAEaylbGe3U1Ue23rA9OYQRhAUpfbp9oHkTiE8/8
jbZ7bLXFczMTiGqTZmnzfn0WSGnt35vqpiDiqLB1OdtZj0lKhhRHHVZLwxM2MMeK9Yy3GH63n/3P
kGoI9TKjZ7jgNNkLk3xjCQvV+cxTcDQOOnsi1GUyalEEdxsvC4MNiJAujsK2KNMomE1ILP5BW/0Q
RRAgPS2cNb0i89z/aSuMM/warOEty/80Z3wS4qTe4bkTFPyQ2uOGimPbPJ6r4diR3UH1cF/vXGGN
Jn79y1VB3X2J+K/hN0RThG9Jau7Nd2pZY7cRbCLRhkwOk3ivgu2kk0ZZIKpksZNg4iHHkBtfgDV1
wVj4XnoXLyiaVKbjv7uKx3vBWUl7yjIc7oGIdgHNJ8KabQbopgUMx/XAdhdzGFFazvtfkU/55/pO
Xq5LlQxSKOuW6cPkPDJBoHWynuW2Ts6Mtym45rf/4f6k1eXhSUWfS/kKnuA7lNuPwPIEBtQlx6N5
9uYPJEknTZNtR2qhzzHdZ7JyGHsnjt69oLXPVTSPeXLx7PNgVQ8bxmRc7izYt6dEx044uN9Suw/s
D3JmH2bR2rKxGoDaF9KRZ3yQAOX9UJ4zho2n7yyrupb21Ct4hDTCAjqW1mY70cPH4r2Q7BX55hmu
RvT607gfj77V/aARZkC55EXtdohrAhqIailQd74RiygPVED6NJgGjdvKr1GMCcyzUqkgG7NoP76I
GhWMYF/2DnqnO94F6p/vjL8IBwGbnjxB885/pgMhbrI17MkL1iAxQAyWien6GKpE6czQXPe1n9cN
n1+Y8uhGOc6Xu/A5NBGNr+XjJjGvIgIybIlfmu2KqlS+RA3bCq/QmgjHS6a6jBRghn6r9SfJxUXh
ohV7eSqw+s4JNOeSlc+kDCmnqdbebe7otBL9lT1NDzx4FinVJp3JG+4WwXPV07XH0Jz+RG4QoS8J
m62JEMBmghbKueGycvkWYHfVMN9+j8gFx1q56ATmEndtIuY0t9anIqLz0GwHUHM5q46jIyj2cG8f
Kjnd15qbBtrpLw62spVJOq48xbZggQ5rV4ri16nQahV7IULg3ICYkBnUgNdeN5fU1NcJiF9z73hw
OkT9QNCeQM88TbFZShyYNPpCOL+r/edLKC4jb/CREpG+DIwafOW0mmRwkd+SQjusoNsEzdixjRUd
Wdlyn1dT40IK0NlS66BzU9B4Nj6YwUj8RTbSapZlOGQboK+THyaYywdKoCwW66NFtkBvJXT/MQ0S
YB/GpfZ9z77pY6jGUqtwWKFlHQM8aHjuW2gZKSKdze+H5ZqytRiv0Usksi4v5B/2OcL5CzsZHPK0
64yVc+Hjtf+T2qFVFxGWEzDWdMSGaXu1muXllxRsNMAxYZVYEkfuLiHcwy2B+OePdbdUQTW0xOX5
uATzygnH5Pb4gFEcM08lKh38U2Xm77tgBXBYomB3V+B4UuWlY7AO3ZJWtA1GR2QCq+ZJgmsYrlWs
sKv3C2Ri/y4ep+JnciuSeVJUKYg9ztfPpCGUQNLhCgd82m3w32mWhspzON/U+MLim6glEV3pF+Pw
9a7HFj0rEl44Bpn5+CC+/S/TKKvmxgqc4Sk7BB7GDmBBvqdjEaX06THSn/vvbcl+VNH8QkrXlK4x
yUara5wgc/6vzV2/TIfSKxvBRRSfqjEKl566ScFYvfYGsFJcLvFLwrvQC9qJEY8t5RpVWzaCDcCt
xtkfInHFFVdATVMX7blhP69LmpF1p5dTaj9CWdxBM/irvHWpLeonkmDvBRd7wD6QUjjGQyzj/hRu
W1rrtvb8IBCDIVPGBSq6mGLyaM+Ch6ZwADjN8JvJt7k6KzF18/WMq/MYENk1MGCKYUo5/ztFEZpe
mSaTyM8MSZGqcOmAtV29I/wcpPmxy84kCY8EF85FKZsXAFq7fZQkx40pL++HjLWFZ6UVVmhnRIiy
/LtpBWp5XHdGq74DV2+OkC4EYOFOhFJnw6Igu9IEOD2/de3++FKtgN9ClRSkUvvGn2kEs7BuIR2Q
wSjyx3bKA/dDddAkAVNRs1pZnLykhsUANGRrd8naIOPLLHTJVzYkY5vjuho6GTxopVbGFrn7RPqK
aS0/KpQC3ysED+TBI5MEVGEJxHTs4XEpgQ2X1WXxgtUV1EvM6Bif6BD02VtePHaUBZMgHXWx7j6P
jjMBkMzO03m9XQmFincBVNss9Qiag+BmLdUDVePCpMXOCoo/ZAfsF2pCPIwD915sj6bzYfVbjcqn
r889xoHbZv9qFuL2HYTQi7wB2GQgLpm5k880lQxMZIm/VeaLmp+aLUa5j2dvggsY5gJ4il2qotex
Sa1Ss8gXfVzBhNO0XwneptqnTleq00DafoXKcgLE7zDTwd0gjaZq6PgS9yU7a8ZjlVS9w44PK4qn
LvXuc+oZ9iDn8rb5lKJ6Qwu/lmphUlm9IF8PKroh0LGW2hkR98QCWgC0/T/mtH4oXbGcGiHePYCn
ZEn7unuN6h4E/VhGDPjOlj04ZGvW6aD3+W9PSkCC+6rEGEHOTXoMWCgu3Ik4VWSiz2su2A8m2fJj
tvAxkcmJOiBNjiYZ4iFgJ+VOM1+z7M9mmmc3T0DgHXwZWY7d76wcXwa9igaLYztzo/wpiMTOdsAO
lRd+eO0Dpk73Ca89mu0LY5p39QaW+mF8HDg21WK79a8/9eiFNog0oXnXEsuykXenOyUVeEOboGyZ
w/zmFfx7RW7B5ubGOflbJtg3R1+W/4xcE/TluN8kmw+gagdMsH+p7UWAJZfF6XP1vODwcePMt2hl
flQDkaD5bgCojBWq45q6F1kfkJGJfCM1YrKbecZnJxJEUta918GKXcKVAH8wexwWhBpP7CohFWUP
EJESl6bH9fMoMhteMRn8OTc0Bp/Iwl11947dFsnFDgbIYmTmhY7m6DuAMakQqPWLtRerkwuaBspC
GuDsddGzKA439/zZZVlBFYRR97POxPfoK74P4nKWofVCtdoMgrKuH0hSd6ZoApH3GoPp6P4GfSQR
b6wlgWkflrW+Iff+5PwSLVE2qcShydFDlP0tOsyYEkushUlHwxVb2swNT938+I+a7FEwDNu67+Se
aOsas7uMkH3mUhfMD9iW2+TAis8ksXSNLUCy7Ec4q6pE0U3iax6JJRqqQ10Wgn/jjECOFXFfHgrF
vu47LN6Skz7EZ9gcMec670GYDEjOjbyFJiO2atJYx9tOymUxCrRk2xt/YpiqhHG0vYAWH7ugWRIH
gBGx6x9vyLo/IDawn6PDwk7ntsO5Uysb3sUckzJR+c+y2QLTMQovSLf+1QArek4nc3jtNTLr0ZJ5
XeKzBi6i7iYCVSNSeC7Toyjj7PCwlSkMQ9fyk/qj7jmZJpuJrIhaYbpgwC4dJ4U5FvFT4K7fqLne
2tefKluIJY75aACjVWTmyfzAJGW3wJVf8p4tuWQaFqPUkc6fr6ZSRgmfB8I1qHHRJj277q+ZSJC5
5mnOjJaKoAr508Sb67JvC8pV0Eht0pbEeY8nIh+64z8MkhF8FKJsSCCT+vBUYJXQPxvBBGSeuTxD
qAN1DTQqeDyxRnMd94f7LyLMZqb5qrRkNCtLmItjYHsejuQAoNjZ5arlb4QgBE4GKZ314qvbIS/v
suCc5y7KHqJOPqPw2GA9VutPZXu6ffac6f6KHchTKy1y1QaKS/7gClQtHbq0vxcx9Zl/IPQIxxpd
u332BPJvT/gKZHk3VrS5OTFihMDeSA1pIQEIJoYBk+WFaTY/1xI9XrZVL2BmZgq2FuFEA4egPy7+
umY6UnUf+9+R4lvapi+yZceojObQPnM7Kqgq+V47EsqQE+R9NITuCKYP6ke226F4lx/LcgV2c7yD
iXaPZRE+J406jxf0s+BNWRXfhx6Kmo8lx0xRo3xMyGeWDuF+dcRA4xy1cBsVeDeTKq6U8vE7oaWt
ZgbuwZ7LNnHojtJ1EzE7/+0BTthfyaBFEc7Wz3H9FNMX2BwTggsaW1eG10VE0hgUcEmFkA7N+O1N
UWzcX/TQnEJ/YwWvXt0AqdmwFkGDPxxK7WNXuR6y+05k4TWikLnFnK143ClxF+uoE5egZdPDBwTb
eNGN1Kk67D4SVybAg3hQPy7Tcg1NzyJgAee59ia8Gu+PW0JsMqtZDaRrdW8KqCFrUCKY9HI6m2gk
PAXrHIH1/VntqvHIw7OnytA4mnnTv4HrNhgEA1DPsatOpOdkJaTCpqeSh2Ag/GM0yDruMyLH9BZv
dESnfmNmQPPkzPR9I3HERnLolXB/XVb6hncxoW/3sXQsyIV0SJna2hRQoJznD3F9pZwH6ZLi0a87
ncKhEoZyikTkfqi8RFVFvyFSEOOV6ZRWKSNX/7fqNIHdkGDR4i92zpdWJmnIi01Rc8TDQAGsU4+t
yh7n3DFB/OV859nHZkhhGwZ+ZK6ZqVrelyHxGCBr5WbIoW2tBL6/xv2Bnta5wC91Bo4ByHVDn8C6
dMcY1UIdEjpjbJ0NZUMhcSKmRYzbc1ewP+MaUd/MQNRAFdDliLygPRsKj9PymzoQOP5ymbHJeRkj
6ack1TRlF52uVmdOGHRAMzCmQrXa3dHO3GJso+Ibet7JzD5zgPm4Lv87bcc1flssOVOtyx3YgcoG
aChScML3hAWsSjESUkhYGqjVBDTLlbuzdWT+kg4s3MjoXo2whahrb7kozL3LSeuD9PUW1Uo9BoWQ
DjPVnOpACBClCEIRgmXSzdWQHyQFn0h86B+/w3cvVFTtT4rnP4ysg7orjGQWnahVCi+i2wyORtn1
Fw1ruTaPXkiNBDBqrY2xNitOeOrjgxRhJSpvpnCcmVpcjRhuroaw8CLTr+1qM/KwFP9emf8peNwW
pvq4xI8X6ncnAVrvW+Uvww4YKSIXHPIGRdpj5SfS5FDoRSEVutEw/fEvSl2jd46+AgEhrijFVBuS
6vlH+SFufHMDY0dhK6GRPghN8gbXZsr9I4fY1+9YBToGF7Prf7G5ynlgoKCVTNMBROCFtCC3ld0Q
JuosttWb3Btknw2hymvpdrg1tuO2M4g7i6W0e/95KwykdDJNfXsLbsnwCgVs1JNHlhaRQ7r1NEl5
oIy+yL4u0UZoZB43YL69SVZxKIEsOmFABwiOjNllH2XYNBhBHtaMsqh4xZi3WNGvzYOFNpfLh0Bv
z7ANjpxmp/kDWxXiE3qDHBI/q15G+TTGvZs4BwXJHG+roVOKkJropbX7bNIva9y76qrE6ya1OWuj
jQbqpceZ1qKK+AXMD5r3JctOpWfZNZCOJ/suYPZVMCxFFCNTojLlxkmSDuEy06CyfmZCkM940ltK
s4bhjxtcTqV8f+D0Ts+A0gzfvX55tNm5GtyHZFf0FcULnNnATDo0/drOGLCAbp1HLodwyEXuiPmC
MqmP6onQltOM4Q8Sk4vsokUmN5sFpKvo8NIJugU+cQDQPvv9h9VE2mdQUsy0xZXgKDggjXodbxBk
1TKrb913lrV9PsKPRGCvSrS62Y3RtSNtgytM1+B/7uPyKsOSmA1RNEwiE9mDAXcDE0f40MalJxX5
hCgBbJyntccYD/lpKXLFMRds+No9JrE/GVrr19huX6AbmyYboCxDYxoQaWYC7885iHbewotIjpsI
DIammqME3zO+8+qnn/WXzQBk9VaRcn3Xf3YzKmGB6ti5cQ/LFjRaqEsNu8zCfr7Cns+aR0ny5FZY
V2OsDhAD6L96uEYv292q4iwCt3QGLmMJX6tL8mNNZK29xbegB2BdWhjQSkTe8FcveBns2yfsXdgy
WtPXCgCgVeljfn610TxrT8PT30KE4jdH/dsgbGWw+O3aB7l3Xjy5kzhR2NCKjRpY6AWokJmxJtIr
0/5TDM6lOYSNZzBKHdMdit6zBcZ6AzVWtF24NEGl3KMj70i6v/aUr1nZhhvQLuCrhsbH5V8IHNp+
AiMe34ymnQ/wq/txxeJWt/GEIrp4+3fseTrkbbXnNDxvf16kRicRGj9eEJnm7yddzQrkgFQlL1DX
L0o3hGHePH/MImRgv9LPHNSkL8q1enGNSMpzYBWh9zwYe2wOzH2khOIXGz9zAzIP9LMOSIlTm23q
2R9jGzDlOcTZH1MfMV7uS8+DAFB9uDJS9r8GXgwJbhyiffnxg4QkzajeYuQrDubaoU5DeYzjDn1N
hb8lWSSrSlhAbOiMC1eXpkZIPe15TASlxwi2WFgf4eOKuzKlK8ziOJ/KbCL69HiDkVtU5c5EWLYA
ck4skgRfk7AskhmGh8Qb9Y3vTFzJsK0znIqUdBki6AoKJ8GpQ184zqDF9tAKl/VfN1vaDUhBAyJo
N7wUmgZAz4/FLUX1dztqed6GHcJfWdOZjBEJm1g4QsIhFxFIFAl0jpb5+SzaSBZHhfGFToGGp7lP
W+xlbpMwPkLe3OSLaxaYHxeP9IPkLS74LryC7abGg2jpPwGLLpngxPcIeCDxxG8NmBhKEdhFmIIf
APkktyLUnrgBLLoc6d5UorFOcfkv4RVd8DSeXIgV4AKYkhct9OQOObib22915eOqhExfUxhSLhp8
an4EdmLpomrnkEfdgPsj0O5Bx+LQrdteap7M9GrFfve1wUe/ZBuY4s6jVdcfYBtZAYW1PbGvWWnR
jXkxyoJHVnf/Las8jjJ2WDWUsGfXtWCwUb+EOkM4FKdhJqvS5W0uaPkD29S2uIThufbtPof8j90Y
CipyOMx4WPUZp3KsjMpfRc2heiru1jcSnpfhd/XPL0BbHHxZSYSAQJ7S3guHAwCFGA719iCtVWHl
D6cPDlW/vt5NqQsYmeOMYp4l+6FQ8haXy22ejLqAYjhRgEY3QpciJ04yz3qGgDy8DeW8p6wubXY/
Rw+YgQlMBW37bKfs/QEtkjSCnOwmOBk93m5MqDmoqFQw8Z0R4yga6UvtVehxV4Tecx76EF3sGVDT
IgzsjeiwfQivzCkaSBat7EYS09206VIQP55/CbKg7vu8GK/KUS8jnqXIIkSn58P3cAFVh9A3vNyC
wQ5GJXB5uoh5k1xf4GDZrZ1ms+S0OHgHDRdrQmrrurhR1cowRRs97mv6Lfg4xNYPe/gfshzwdDQR
dpJmGwuvrzvemvE/P8Nl29wKF6zMAI5pCbiPgDDVRS3z1B2+GzHMURl6embKNmk6UUjGgtMzPwJI
jvuf7orBOvhsuSFPGiNWgAyzkStSFP6PqlOOiYUOcSq1r0AIUJf1z5EQ3I+0E0GTK6XhI2yzX1GJ
5JryBBLlBx9tSp+ZfRONWt8bOZQfix1fsVsTHc4nzJRHWWCLBajklPw6SlDyZURQSwB7csugWAQx
1lQoKs2w2LmDDrxxV1TOWhfpHZ2Grnd9g2D9UwpRWykY+AV0NoUJmQ+p69pR2fXPUNey7nWPuj9N
hkjV330lCjeyrjSVIJsbC5V7AoW6V7dzAEgODaVvNZsnesZ/baZraVqCbbdfi0+rtTKsz8IZHtrE
DHQL7E1Ts0bCAU4tUe9z0etIiC6n54pktYcGyvzTtK55rXUJtWn2/0R7MmTMQsuZ7qvDsdINzOG2
gbJU81aMByF0+tu+EbSv7rqqoMbruqFgeOgfeghAou0PP5mw9wh9abat4ae/m7UFnayUdRArs4El
eBe7IeYeNYo4Vslx7q7sfLZ0zHsYFNQBkeyRcdL4LIOgz/fulVc2qvEmS11sqoeBdAkBn9tmSJG7
xBX3K3pWFE01ISzFUtXeTCIy9ZO7N65hDqZfE9QqK3WsL368Y2RqV2mwPjLDMX/k+JXKMqW/eob9
XxoVK0bmyZmSgQw11dwP8HqqdFudUK8Cz4ANdi/dEhewmPNZyBvoGd3aDXepV8bhwlDlLT4L3G7+
LvIsHCe6h9v3dDdi/dFktLQFyossMpE6VG4qvMGc0dF2v/pzhK3J3Nag5jGZ8IIcJpqeTYd1K7kO
FEWZq0SCFRopWtb6K1HSaQChodmmqo3J+8cfOMETHlplapxRfdadV0dw37UCZK4ozhQwuswL6+V3
fGUhBLAi/YT+Ufv3tOEX3QDBVOJARcpV2mX6jgQ3cXNiTmQ/8vx/E3SGQO6XhkCsnyaEu6o2cIXm
wdH1G9TiQuN+V+iSCO96UnE7PtrBKTi911efgUVv4cad7m7xEtEz/JjbC96Ju79JlGTklnh6KTuZ
KwJCKp+7POwflRqYIrp/B2ZO9hBd7+mujc+32WvpTGM5fHGt+IVts9lieoRkSLlyWxv6xo0XWhXL
qyxdTeerxTJDrVzVHSxC43KhO/oFEd6/L8/GooW+5JGxio3NCQuXdIsEUO8rhGHQ7axYZfQqSGlV
52i1Z1onyaUzrC4pLcIDR6Z37NH+NW9ZYDc/aNXMz74EBf2QmqP1WOPQgt6+x9kXRSpUcSWTtLkA
ST6wPcvSRSh9FrmyRKrJbLluIQUamQEbcrlerwhYcwxG1qMdNMDjBKc0FgSnZP+b6u8bvHuDUwcM
rSLfTGCFvoqPHSTyevkWunnHO3if5aeQl5JMpdsiSZXiukIRnC1ylLlI2OoFVp9+N63EGLv81gUp
fp+VLaR3Al3dZsVs1smxyE9J0/RsgTXD0Ufe756LZWmUYTMJHgCnog1A+ysA9oJuHnOysMMyjhe1
H2UfbSCQ1PhSJ7JTCSVpeWmGfWibG97J6ale66EiANoxt8Ek6VCzz+HcV+Mlxkd6WeFBslBxX5HZ
UYRIEEAKC/ti4iayQsX10z1u2plE9qgHsF6dGir6t3+QlXEaQjkeLFa0xPjvx3RNCVZMGn/UmIIe
65adFHH4NMsb9jN6KaIthFb6VB+AkubW5E6nSUy345aVRgn7DX96L/4C7FtHevxtDqPUG9TxJvtT
prS4lqTM5MQxHtOH2QFG83QVISDX86FgyBEN79g7XuS4/l0L3WmiiqXE9KmAX47mIwyVDK7BJFC4
uIyw9TMcU8/hjwG0rbBDl8uMlfe6VCmUDPv2mm300X/eFhSHtFrdxfcVEDSBx2khgCrmRROciRg0
QzfbZKvupaI6/eTeMCHE0bSQGci4NfviaC1Y6o5F2bpdt5FGooUX32DSJHDJRe9zAJPBOSWvCQCU
fCxZvwOLJwz5QLPXL+5PUs9YwQXKhHFcgCfRKRfvYXgoxgOzTg9Em7rMOAQlpMJ87pvD1covSf3F
JiNEWArHQh97A+I49/o6WS6DD1jAjUFN7n6zQ2hLhmgKBpFt2If/kQ6OAa7zsqCDprEBRJyKKBhF
w27u35838s3Ej19CMgk0FqlkNTCJ+aIDD8saOyZX/kYdBOBKxiceexxRi3JN/FxB3YqSJMQx8m6/
Nb4icycb+eoyQhF4s0KBWcsX7KXeIpriiF44isDWIXfvQ8WFDiS+YG7Gy7T8dG2ygDFTwu2cqlfg
XwmGVG+2s/rjElarLdWNMhRD0/ULBLXAJclfbmQS55U1q7nCQcU8ozdyLjMyOyMnpJlM67jsceGI
SN2xW/aIrUHViRNenpsp0nW2Ew5y5Uq7IRmhK6/fGljetpVoGPqdyJlGe+mdwBXuXNSLEjho9r07
YiSUxe0kRTxwcJD8dM+G70vvzjz6rHCjIHEnop9bIZQrcmmGlLcM49Fz3T92AgwcxyVT9fTssORJ
B+v7s+YPCu68JFMv9rxAde/FHUJZI27/NaEbPn/kZQASogvqAgfpHn//JxL0zuKY62odXV6NGc5F
mD4BQcHG7jD5qCOMY6wFaS9QajO5Htwa6z0D6hCNPE/nAAbAf24AP4Jg9A9QQL+YJprUi8eaLQvJ
DAceb+GQe17VCHE14eG1gaLaEHCPMB0kSYaGq46W63zk9X+YwEsNiPYgeGMaoBG+zIajtygWMHjR
4gp0cyhu3Mts+XMgo3LTtZ0xWz3KU9s1mBgREmZT9ZKdaiolNbyka3rapP14eBY/DyYY8+pPN0Sb
A3hxEGdDQdWjdRF69GrsReM3tiMmFPXGY3YDg+Zqp5a+LRonYfQketGPvGbmZ6sdsQR7ydnI05lE
0+D3+zx2N4ZJ/22Vmexaite4jg8G6/K+JZQ5rxfMuZQ7ULANvBaTHu7hd9pBZA5ZmgQi1YafjxYI
05q2cKgzzHdU3i6H53zBU3QM+ZthIlxJ8EpeVu0DalMsECbOtvt5I5p4lPCRc42VZcqhkURVcWVo
cFlV6vcnk9tj2PfGepleeOhjlBJ/LF+HJ33cngcyryjI/zTrEn1SfouHvw99UttLtWkmDdlaXjms
SgRPPG/oDF0RiIROoxcS14C40DRN+Vuw19t2cXRADm8fMy/60nmTjbc/UpnQqUs81BgSMj6eRuN2
fcdrjCEsOEatdtKOKOkAGAUE0Ad/YUxeH54tnq2nBNC7lMOb1SB9GheYXKZ+KLVvTKPSOZVZXBUK
bn1G3IVBmTNhotttamyyjqPjMXz0JnPfkSXBIfcoCC8LmIUGhAnjb6H1h7w6J7fYQd3BT4SEdmTG
mrqI9HhdC/jKc33fUs2eF9BmBFLWR+z/Ed2Gx3dP3ujBdLoeWRMUx2XN+NFW/ZpvWkDmS7jaiFDX
mF0vS3CDWK93ASxtZf6smWxFzXwu8uXcv71z0bWDjtIqEpLX9+pZzFgldkcs45t/1GmKzbmoOMtx
ack2SQVVbckgCb0C5vZEwDlEel52xj0qfhRUZAGKLr+9rL67bGwotn+Y1C/OvDN4z9347gFofAZD
euV9N1w4QCMFOzfQ+KAInjaX4BuUKle3+GYP1sE8Eu0F4APD7LuJ/UZmdNO6dwrDZdutl/4AN4oX
6lKmh4Nc6tlSTIMSMJzIFDA+UNoxkBIrPGBGKX7NWLSusRaCwCxN0+qw5Kw8Fi+DjmnMbEibIKPr
pLNd1kb0Bdt3DytHNO26USIdTm1Z2+zjlVIyG462ORP061AOAbRos+bCrnJVQnbOb8t6ryZBpEfA
SjX7eAY6aly1n9lho0V1NKSaVRHuvUWkYGxMB2Gu48ioM4lXT6TzqP3i3MRhL8rEH3rcyi2u5aPD
22bkEibLlrCXK3D5FtdD5sfKx5INHnRlL9eHKHonF1thkhtTpFFwVOWYHcOteqyeK+LnNYtumuy7
duj5ihEFKL67eBXpv/LJaZBMsQTdJheg7mgdaIGeaSZYimBNZYtfpfXkSsZyAJnzjkEjUG+tDVJh
KXlZV63jriTVn+RRAKlKCb7lw3Z/TbGfVsffozofVSMgh+eBRU7fvWBTr2f+VwolKD2lPC+4EMH5
IFj2PkE7BAwZkix+WtZ4tme+5H0RxlNtZya/yvIskO8eW1irHpES+r52ziaOwxMjmaDVCBH2BZlw
sYN9nOPo2aejpWcE4Lr2bGkTXWF03Oxpvj9YwN/GDsNOFKsGVTKFs+tY9+CTrMJ75DbHFRpV9Cnm
gYgEkMb9dpi0bPTpgZ5AsHIiBXZcWF/1SNdpks/FYDiCExxxuLvqgjAtvabz+orMFR80ySEf3wEw
bc+e6kUPxmBUtSGMxQCDnkrvIgV4YMEUuYIj48RwnnFlw4XniD9LdE1ILVT1srtVHpgN8/Ku9511
qi7f0zXdFY5UPxdlti3WATTUvbY9SeaLopIsYklxlrbm4Y2leQjXFtUCYzoPTR4fjup7+ptksr0Z
qo9ZbT7jOlJtk8xZwRmLhYoq85Lki56rUdAsnYl/y08GW27xE0k7PEwoiF4aTI524y82ZSc64ovR
bYX4napyy8zqxP8OTFzi1gcY+/2fp7fm1Dr1krx8tmeFCFRntqhZU7yhybzMq1PBBisryqBVG6jd
ttGwNnBGp0FHnZCgtH8NqdxsUdK5WnKpgbTCyIJwz0HuAQONDuHp8WJKjcvfyd8TWKbSRQqoKRIt
mU174dKVmn0x6BmIX+dFqsamlaMyMV1qXX9F67ddP/bHGYHT4Pi+c6o6luuIdRvFTRGcEE2LZlPX
owLFAncCgO3yEZpqLoweHUr7OOvI+3waFeqax8eF0eOFdAytSNhmun39XjZLBqw8ol5zRmnntoxk
dQYcTQK/o9LJibFMNQx44j2hVkvei1OJjzZBYU5/0hKwnYJsKi787bQF8EV0TjWXev5Oycvayqew
LLCwe7ThJSYmuc5dh0gDmGRQDaizZcHgthbwF9qZLb23UfZF5ub8clfdpQziAU86hdwmuzm1ZHVR
5P7EW8QKWFnFl2h4Q5/3GOm8VRkc5KqZlqu7yR37bJcCYyPQUI6TiiRR8jSn0M5CfA36jexkg/Zc
senLb8QH5YSFczIHYIB3vBiyacBvVGYIc2QvEwfJPZJsVTFp1cuBDJQs3rtQVZ6hRm/PK6//Gnzq
zrs3NnCvdmIHRsckGXZWAsbw62k5wFKoaoswb0lm/sEC63Lfwi1umkyd6ouyBv/8V4637NdnRVLW
tNb4BkXh9L7fzg1wsYJV5xD1NTfQBbIrtMr7Zo9VEb252OIolVxdMMFPxD26yM9NRb9tBQyD0LaU
zQNiNTTXP19TQL10sQje+7vWDRFEYZf6FX68xPP192L6V4azcsMqAcH/xqkA7bIlSPARKp6HhcyB
aEoO+4lGN7LCXUK7KQUSF6yv1Bb8Nx/lGQJresPuS6dxWDVOWCiDhwTGozVNur9Ezvh87kuuAdZe
x3ajxQpwLZriWqlIuS37MAts7d14ZNjA/wWfivslpyReD14SeEJxGkNeX7GrfptbaWxtQ22X2ZmT
y6SpWIJ03J1knRi2hrHE6gZAWmGXB0Iiueg1oE3Qg9VxwLWKMuSWiUP9grQCUKwnp5drlMS7QO1y
HuX5XTlfRVn+1pSwSwt2mUOzpRFc75kGKzEUA6Z8WfVfjriIPLRaDneMAZlGrAFpslh2DsxEeA5W
TIA8h3yJUjyNr+sZrmcjVOMzblTvYwKUXXZLRWugUFaFxSIR+1WV8G5in2bNJ30ldd2zReV0jajl
TB7kA7PCfnouaaGjJgczmPwzVmRUeZzQ/Rc4AThx0h+vO2hOb4kmCZd+nJM4MJUJ6t8GikExDYeM
HP9X94qRyLbXwV3QSOiTf+7keg7mwxKRch6gUR6D03wvZ1Nkox+11RWVlkxxiq75FvcP+300JhgX
mWL7Rg81XbyzRVPhYE7K0jgX2ansKEVwHYCgpaCCoTEA3GiLX2Jv6oqSAKrMqRCnPQd+kUfQF4cI
RJFUdPGhvRBUj7miZIWP1/0/b+5wBXm/K0tWvbked5WwU1rI16g5SIzZ85X08GVbCCzGtLKgXXhb
VmWkUVEq2z7+A/7i6PklpUk99Oh4HoArBMnMCdrjY+P1iAJe023sR63C9z6GCKlB1fUqGqQt/dnK
IQ75R8UnUyEeSH21zpXaRSmqQPvK6B/vn+vPjVZ60dLBzbHIbZpjxDPcv5GmK8csAeS/cJyEtHef
ls3YJ7dO73FxbtdtlX1pndjtmkSXYS8bGpfWcLWQnVy0I4N2zyrDSOGSMnAuDatgAxNDGYdLLQ3c
xubzI6C3haVIsnSo7FTOlQvscnWNPBcpyyBpRC+tBhbIk730FtJG58FjKa+mJGpG+zJNHDK4VK1m
hvrJmZzgMBmO1Ijua8D1QGoFZ1k/nCJl97vnOhTJviVrielP7j9E4FE9RomsMYqUjS0IFHJpQ2im
Aty1dFTPyJFpronoEuw+VzOVCzRXb6iLwYy68n7Wq2jvPc9vr5TqZbmMdwbVDcFpgdfP+YuHl/xM
fDVsPtlfaexqFo1AJJFfGoNTCPtAXy9hB6jP/NDGO0KeHD+DSmpKmme2/AX9hEG2Z1euJmivanvp
9upVDdpOJreGydw85pTcxrbefMyYe768oh/swOTuewNokUQ60KsmCn7gM6i7tGfjCLn6nbAnAUNX
0M2Q1aQbn2jJbvMQOS+c+2/GilQo8+jQcXRii9L826HXmpn7zIYnL3fMvP61zKbgJTG1UBLjhkYg
VJjplP5jnd64PUMHySCPlEohz21jjuj5Kg5dRY1IRr9yPORocDjdn2A2byrGBkTre72+r2/gDL32
9m29K9RpJL1eY5NlytBM6VxD+o2uYYdJp1nEcKeOl+iGXwhKHJ6jKfB2DSmcvoXj0WDrk2vYKEEH
cDkWWWgVb6xS+Lnt3bLbpgB6QPE+AKB5QZ1iD1I8lWnyyg8Iqs9Qx8C3Fj28MT2zYPLwQUzUpPAq
on4Yu8GrBxu+hH8HEh99Y3pDotk45m4hdelZdMSpvx7DfpQP62djRJd5GMbtUWsBvh+FAUdaWM0R
yoSmz2RAMk1Azh6N4OAQfstT8NO5YjG5+D4Ll1N+nHrGt0OUIUa2dQnSkgrGkkhpiIB6jJYD+Rb+
J4cSjGJqy92I0iZe41HNNpc4BM8Z+aUVcrZjK1By23c/5MXh/m83WxQgnZE/nasDWCZxEmXei9pD
qWXzRjPhhnnFPn8KM1RU/6knOkYMQox7ERke6l7dAZ2Y1G4pB7iTvAWG58ZaArilUExRGltw7Wo+
yLXeXYfXcGcmAP0HNT1o5O/gJGdzes1A2kd0zDCxsIXzncPAK9VBhacJsrKAoHkDXYF+Yc+KD625
sr++siJxfKYoxD+u6DqvB/CPWy/hrPsX/Pie7eQCncLgdWhnmz3B34YgqnhpY/zxuNbeSnuUgO7b
PxOOen7d2Am4U79qzcwGeX+wb5y4EE57JgSR3mOqkdx5uqXUO2nwPeQPg0waBoY94wCjInrrJXl4
+izsM8dL2uP3JTkUbaZSOGZC4qwKvlc2Eu7V+/GAnY9CnkMo7jfGDu0xvVpvZEPbATxaQykdRZ2C
wJXSkAjD0POSYB8jhcKoa0s7GUijyRDIiAf9oF2E1WSmHRSWyalcBnaDL0yI7osqrraV++pvIj8T
UDUaRCXbEMhBs2MBw5GA0JrFut5MSXn3Xc7C/9+x96WSIPsVeojsUTHjIqBst+Gy3VAGLu6kxNFG
WiEwxVixWwy8m2B6na6QYLtWgCfzfZIiDV450NGUlMW587w93+qyIJKkdQd5lWp8VXlWTE9wyP3b
VmoLLCTLi8BYGlhvHnnVt5KvgKtlgUZ0bEdSnH9hHorDyBC+7BDamfxuQfkAKvOZMR4zR6brgKci
9DEnw9Z+0mnlubGUHyf/7yCZoO3MT0Jt4/GzNdFNzF2ge/SKM3dw3OXqtzyLOM0B2tux/HYKgBJC
q7KzHpqR1JcJ1YCAVx1iaPRnBkQVhlk/GomW4jcY3XA8K1caPgeKVfpexk3SGYxAypg15iza84ME
6rp30Y9UN9sCwwr+hOG0KzUS9FGYutbpaAIVi00WmVdFWsuDGpij5C3q1gmaqsWoLJJjE41UH1/m
kVa7dzR0OrO0RPSeFfYR8vtpRjZ7u7cFRuadWoJGXvffFRhnzggY4CWc8WmXGTCyiIlz3n+jM9qh
VQjjRNpnfWV4pLjPkfphpzTDL3CG3yOB7YJSONm5nSr4eHDMvzXvI06wbhFp+Ta/JDI9+5ZJBrY7
g2QguCrhIcVfPA2/Gg4XtkY5aUjdw1PiuDLIyKzlEWJbuZwN07avIG9PXHHgDE3yDz8XDOSqhY+U
uZSgatENFtSg2u2c+bw5qykPsePIWmVdTHRwtu69MIadpvQpUk0MWlPeoPgsGpwlAvmhT95XaAxo
TjurMA7JP7Nik1z66igYeTWhqz95rGN/F9o5Bzm1ohSwll9ye8L9jLYhhVUImKhqju8MAZ9dq5me
aMGT4Iw5+MvI1hGVPi77b/6SNKIipRvC/w3SEBI5TXidqa+glBrYAwu+sLKbunB/yb2RIVDxraCR
2Ohhfb2TyGxa86UlTYGDQj30x1sJuYElTjUUPXcGqYu0N1sUSHcYQXDIg3tbI3PMLiGbDEbya3uX
2/hsnAPtWSls5FR682aV7J/wSYIKapR/4NV4AqFLYPfBgW9ipQmrCNOm6NPzYrmexIoCaPIvadmc
Aq1c9ebkLi/jnhpPINlArHoYi+kKFvqeWdurhzm9FZcyl6jROS8D3f80gI4TPYpas/UCYt5UXumg
/vjb/enzkh8PArtvvPNSnQHeHjs6e+gVN3KuF2j+DkAqHQ/7c/grX6hpijmwN4wt7m/qF7n2Nzoa
mBxUyF3Qtn5TAt1NQmY2Bqrhu4gqz93Rjv5MTWLG8ckxtfvjJkmm/DIPFNxV5tFXkVcjhOQMHSO2
WLoHiQTITL90Zt+7ll+Dk5Dp/xGA1tZOAdKiqgDxpd2I39/fYxZgiZM5wEV/SECvnXXif5ZIEpBv
SlYz8mVQCUN6yoBxv5XVrgSZD4LipTmO8mW7YM+a4YTjxXbHW+vfFkJMUjj6paUABbJ/wFTNlDVu
gkgAULbykF/OQOU+nNKLn0P3Zqak3JKEvNVBtLZA95lSD+/bzxaf0oCop1wg/qKiiuVDMZo+KxGC
0a2qZUCDDHaEhc0ZYF0/XbdLGv6HLj+T2wi+BGVahx5PraZv/+alvky3V30L4riURcTfgG9BC7aD
u/l+zJzIdKJB8TdOIU32u6YMuzpYEbR3YK6JTE6FvfR+vo/OQ2K8VDwzBR3QEqslG1ScPOIOu2kA
49HgxZpPdmHJkT8NQ+w1HKf45wEJrUoUgAtLs4Zi9culdmf2U0TzFBfLOS4k7cTOfKlmTkF/6N3N
+RYc1BqVa8L/8QF5P58gPmgEuBCtAEXhW+uBu4QC1KxSknTFejUYfHjRPRqfqhvU8xNPC9wcajH6
yp3Jh4Ri5YwagK4aVlhNjoM2oGuH6NjnMzYXPvg7VpT4rB4+N3vI2PxMUN0wvs/B3HW22THcc4FZ
yCiI+sk7JVS5GI3Qk5atfTHxmX2Q5YQm5dcKos7RdI74nODuFBupl4dxCUubLVUVG+cfXCMyC0OU
A9aEe4J9gcPNpZ28q3ELZnwD/C79pZ1JnWiv/ko7IpTb6liO0YiIEIWAR0FAvkgPYa4UWZcj0auy
xW5AC/N2ANhazx01WuqrhOEbKl6csSPlhMYnOPBCtO5NYn497WrO8GQWi1wer+O33oE5SX00fDit
4R47wlDzf/Jf513/v0/iYT04daqLNk0vAa3nPrXZVpr4gz/vnsnDUub3xpub7vjEFvp4FVxEkWIz
l7r6RDbCW9a4KBoq5jiQ0Tjn4t3RmkNeqHa/U5QtW/BL7DbbreSKVjIGArhVaNgwcYbkDF1JNeuy
IyfWxqdZnoJILgL8X8S0AipAe2nZV9GTeQum5eog5pjsECSW+LDjmeZmy19dKq646B033YwkxNHc
i9mBREKELXrWB3EeX3soc+PrJWJmBAOgvUuwcLI849wUJ9wM1AIwcIcTrEfVQSSuJ2UqeMfF7oqb
dRciJoWefoLv0i3A4vtlnqgnnNyXx4tWhs0j0gx+Xydqdb1tXIMWCK6kTzDXEMjrcnzWVBPE3cvb
AAch1KM4gcMPTCsrDMtc6zsxBM/8uM6VwPHKsd988ZzaW864jbbXDT2ToEbxNR9Zs7XMpTlU9udH
FDPLDygqtbq83WAtar1IFd6078tFP1E4jiokmlyNb+XC49LCjKJjgwHpGzbXxZ+FdLSAiva3NZCI
VAM8wSeGVRWx3t3VCXaKGChTF14hgB+kPelPaA2mNtUwdHmviMBeOD6bkaaLRMjOZPCBmpf72ici
XoLKkCxZEAv0Qb5F5zRYHwngcU/xi7KmNJWxACiQp0SRLvAVmoglwVv727xL2ds1PnbJGoX4Eyw3
ZsAG9GnnUr7JjSWTQdTIT0Bz+BVnMiTD+adElaGTDWACz7rnd4sBUbxlcIhYeqo187pQ2zV6atzL
CzJjLvPkeXhrYlTgm4iBfF3pYiQpGtcTFDOqsruX6YmmURQzknrLvD+H2mYxcJ2s0Vl0aFjxt2rU
AADSJ6/XsipbuHUkwy6unfOkRS0uDb37WOOPBNmjWhFS0kf6FkFkuF7iHuGBYQxzYTx5LoFFmj4a
36rFNeiMvE3gktThLl3QJN7xgfTLttp35DQRL2kklbI3Q5tsB/dQoYt/hlH+VYvU/AvqFZPlz3wM
c9L51Lw1wqGAShQ+excsPYMlGNsh89g4nEcm3qX5IfJYjp3rPndMjyAmD/rHaG3dZ5Bo3Kuv9fPw
0sPFJMOnxIraR9LlkBV+1PqpF/usvisB4kJMi7f4OURrCaW9e/Du4LTHAnOQZu6zVTI6pQxXV5yY
lloCdcXsLzRBdukceSDwY6yD14yO828qqcTQLAe6y2PWEvIr8sqlsh2zJV+yvPIu2hv/uyfPV8KH
EjHZUEUgY9iPJMUfsutCIz1U30T+wxwCI3bGO554nvrKD5f4x76SDAI2I/NogDpHgfpLok1jRXTT
DPtPHW0fURFTEfFq3i/eTwFNVWrmTCS0PkET/YNvJpYtwGXXUE00Ox7M3XPevfhih/QXdvtrhHCN
tWebZLjMjoMuz2Yn3M87jKAZvpd9zrCLZGr1GxgrbbUOQqd26x6O+1WLHuugHRHB8MzbxB0Pe7Fo
desfrhucXTZ7VGVYmPLNJW2qGlCZshXVX7+fUIeKI390xl/s+RoksGpRPdL3Hw+rGQYp2OQWmxqM
5e4/BJZQQfpMSVvKPE/Dzo2lNVe6NZZuPLSskW25BEp7Ml9g6Gwj2bVJAMyZaIOfEjp01otov7Yi
ion0iB+fsPbRqpN2P5jrTpOAlxKzRudO66rbB5zEVm96fQfLj5pDspG/xpxs+VbKVZnyu2s6qosg
B7WSrOMGvyBd53ZWWAziFJHHx/htkJ44k09M+gsn8twl+AreRdfN+wr0z+TX2fjaD2ANsb1W+gAm
UkWe8oc0kpVOTjk1/JSGOhqN+7/BA6GX45KmHMRrVIIe9xAQ8AhrEEcL2VOHzbOEEScqpns4RIUq
NS1CMb/EqG5GgEjz8ndwbZOhLjwU0m/Iv468xPeQMV4dbfn4rd2llgj028nomjLEl3fT3TiKmK8W
fmU54J29I6BHig+Y/FN/gB/5cY1ZyWZOKJCPgPmhl0K3q7ZmNyOJkpk/CyEuOnPsuSh6CrxS6eMy
SavbbmmhyLsEPI6w2sZPCqf5Im4dNA7lfhyikR0GCWtDAcMR5CKZeNx/mPt0LXJr2SAv7jxUPVQe
agUpCiynT1h8PY35IiPn+xQwk/GYnjkLifUbD3c2YQnJYMO5VWoi0ePiOrpwl8kSSezINILv8haK
ex5k0FoAcYRL+WYCQSrsQK3jXrAYg1Nq7oO25SxeYtMyQdwO+XVCNZLenHxsc8bi1F9kV6t+ZnZQ
x9DutYJBLso89igmDwOyTpJwVwYBzOgLYDS6x0tKHN5B5Qdh4Ly7GpoQgR45M5DyM5iX6G1lQ5fM
hIwpSxvghBszfItb49uf3taYCPJ60zoF+37LnSYf69FFEfzCDNkN+4mdRchlN4JBCdtEfrZIUASH
BArNALnQXTM99UmPuYVyFNcEDy/5VeowprF1YKPFlZkFpMuhnZ39eXsOekTwRLrjHhlGaEOhWXQq
UD19bYwesVCNFeSO+IocAm9lpBZoBJi1IoRZ4+GrJPdyXF8aYBbzFzdYduZ1Eq4f5GnZHgekglHj
SsOqjn18dW+distI6pe7g2fMKFe3fXZMtc01PvttsUq9BOgoBfIp0L2XQLwf1vl7FQSmxLpomRyI
+FGrfAq4ImPb13caqfrB3R0g/DSaRGeJs5S0FzrVAhBcXjcO28x9euetSXt6+LRwtm5huxWBylan
pRahnBuJCwxJZ3+6MW+1sBgkbwgExd/CNTnwsXxvDwV5hyQQTvqBcc7d6ZgKPMNn1ixq4Mp+YNX1
aJX9S1pNYgolfNgf35cbmZ4NeYCBpN+RMhVb/TZBmUAlrJ99BOR9T/qin1ieW20TGZUc2Pv0BZ8V
v4HQGF3kQckySo3fddUxxevZs9oHF8iqSWf8mSqt/AvAJcjvyA1n8IFz4SJNPjd5M1mOEkQXSGTu
3nzlPYzdIKfH5DUTcLIR4rc1eC4KkTjmuElwtvsLOyEc5BKxOdUWrAuW9rXuU0lv+sSDZHjxoY0t
Vc/k9A6BMta8sVg5Lla4s0mP7BFYFuooFC5tzN813U1n7/gwF/mwFgSX7+dqkfjBTh1grZ4+VH+K
Mahzn43MmsN4CHHjqSmJNluOntg+q8Vuyi/fs49OnmzByllftlQCVRyoLCRdEHZ4gpgaj+D+pDgP
+eTGVS+h/iQV5fez9hKKI5VNU9cPKRriOOc2rLeJOnnmEoRtKS7L3zL2a12BYgXOkdADxpcFoQ6N
Q2tDpgRD40FymylBGEcweCaasjeDbyrciuwB3labCPU91jEGZnr1zytxt28gVblRcYNWVHqEw0KB
Sn2Nv6a8Ufsz9MZJGD4XyVXDSHZti6euqrBxWIAH7/FesNaMmjYZKJteFJ/bSmp1A3k8OCkzRqz2
aXW3JHz3R5BV7aRfoIuUws6zZQ7CBU5C/rZpLymplLe215hBrnC1wKg+mAB8qEPIJ/0ZHT2DmAqv
210eUfouvWZsntwU5YOMzgxQn9q8aENt4VAYlswTjkbw6QMYgnlOTAYp8uKOG/ASIvI+dry55t/q
grbLYmryIvTbOHol4q0+9lv99zIvXAkL8COTBVnxVlKjGMNPWbmBUAMbcIFQb1xGzzLXWtnnZ7bg
KsOLgnmHwur4rYJzeBcwSBQ4HkxQ5709Hl2L41X3qla+gZqT5P/xxokCkusyslBerrMdlpIg7NMG
FD3ur/PlcKJlPC27Xj4IARWrEwazDpXvj3Ds0kivQnTmaKXJhpcW1ZW/i6gLaNPTv/hN4tinqEZv
x1FndCwslwwuXMNAmfroTVa9F/tFjqeo08QV9bakU51sEvA5Y6VuvSuA+HwQ11ePgWrTv9Ambwhd
/mMrip7/+wZA1qKDgxZImj10DLcxuu3/AiTZo3ve0qm9PtjDlZH+cKyX62Y9JpdJe0AqvWjPTTwA
dSu16K/nVaynl1PvuPr1rLmbWCeNqa97yV7mMLpvrCKDgOEA/FhEI2AA6vqgBD4wQClMt3OzrpP5
YUko591kzSR17VASsd/Mx2+d7HxUNwR7wQpoY22yKBB1QIKaq8NcOzHywrkWQvMuqeKf9Aixjiyc
P5EPGt4mrtEdRBOLgyOJpBpm5LeZgCSIw7ISc7H+NIbBNdcVRjxbt5iw3Xf9AzzJJvE+C7E/ecfS
d0tRidYrmN6wYhIQabZuvn6pna5aoKhOzCLyreWxBkMc38ywPAmKJOmCLmUs8edmMguQAEKnRJUV
0qGP+B04/6z2X7Vfyql2wv0Tgsgm18Av0S9gLViKlqugKbcnK3UF61u+8db0vJsoKENw96eJ2Tdg
PkKW3796dAFGD3i3zT0GAy8G3RkMuSNmTkOMDp7rKrIYqamjA5Lze3lHvhK9ZskwDM2u7uRa/ibR
qLFizlIJnfZWOvga/+mu9GqvTsnU/oNjg/bFJ9vW/wplYtrqnROtGEJ/wAyf46rhWwF35R4vSZUx
TZLE1R52gf43kLMK4uvhVuK/CSHKjlUybGcqIJUqoJRmpXABNCU2WUZOmr2vp7R1Tb/8WfkbGTby
2+/8h2hL+EBPKW0+5f8+coxvyqjppeif2Ip0Mgy1CXWI0Zd+6LGt9L8Lbo24HEeYYEW790YM+6Fb
+IvgdP9VlbddfzWtzS3lQl/oLACgem/Oi22j1yDLwKiaMbsAADcGm9oxfVeZUjWF5IXZZHQQ84WQ
pByVKnFyLz0/Yh4PvLRqKvy2D8KQVKvH7VI0yf6qvvdN1kVzG576aQazPKscVyMa1l1D+21HiNRN
ds9WcbqbZXXJCbFil5jLxR3L6eBTGjLZtkmniHvLxva3L8rSgpP7/MewItuyAnbIUmY2E8PvryW0
5OPMrHcqkbtuyw4vZe1BgpMbxhfar3f/kPacJrvqnKultoOw/Gfg37tU9aQLRKOJhirRj90Jo/tt
mnhKdblKoPdbFttncGHisyxKBv80IhfnFDp0J57Mkdk7/zChQj3Q/E1vXc+ROi1JCdLEKGUJDeAl
W+SKo6DFWHt10Onc3d2+zQaupym89tFFy29AjJ/ENY0KUHJXA9Uhbbo+rKaTLW8esJqzFiWf/Vcf
dL5uuKFWTUwMYwBAXW7D0nZybo4gqKxz8cvugs51RI3ymQusBo7SkxqV9dTorTOG7TgLWFTCFZZY
BZ84b/tlySxb2JFO/6nmpuMRrQ6hd6/HsZiIPP6w/YFuJVID1SKDT+K1Aad53iOss+Negq+UOfeL
zzu+7Z9+iiBJTNUUv2EqDvaZLNYIrBeia91QJtPOJQ9nCBoqAoFxldm9c2Zm3nZLBThKoXKfmy04
8alMQl1OQfqWVIeyOj+ypKdRitEtSwR9bWbXtwwYK1z1rGNuCv7sYkMZESU2WP8m2DK5PK31uVZt
6GHgqmfaH/gYORruZhDThx7ow6R25umaF+2Gh3QIns/St2/6iJlT9vNyFjO2SB5B3zsJq/J9BNWP
yaqMMTTyjRZ047pXAUeyLrw/N/bRmXEAseRV5LF27tqEzc41tBHg1jT0o1UCWDw0kFnz8q31Of+L
1pOzTNuO16E60QjcGsMoAoS8ZjFcKcUshmwf1bCWvCxOtZPtQt8szG+dBpHfL9e7xj277Q6fi0bb
hI2vbXAxIZQEhsE/cUgFz/qQoE9YAkPir1ne9O/wuLFk6cFNYJM8mu1iWH3+t9/2kLx2UzEPHFgN
qGrXuWbliBnYgBi+GV4xEMsrHhBww8auwpSWm7ljilMC6lzqJTxA3rUuzpi4RA1yBxoDwWV0XL7j
IIfCQn1tQbDO1hco4YaE95xpE8/CqRLTaVKLmdliHXdcatt02/HBqcm5OnmovKrt7g8JFuwrK519
Jpz7eiWOqpBZxs26KQK3ET/uh8GSA8A9bRnOqE7UQRRCC59qqWj4/CSnVxU7c6BewpvOND5MxWvx
rUoC4GVwWIjYh3rxDMUXJiIAOxHsST5WoqI6KrIxhX3oF6yYhB/gKQ+7mU5ELgOTrEDFOPOdDJ8k
QxuA4Yi9JUI0+De/UWKh749wf0wSbaW4dXBVBmV3dYuddW1Q85Buvswzc5uxjSCs9LX93i8nDWoB
pbKXJGaOc7Qma7IQnJgCVGMVMZac2PSkC8Ye8RBK9tAIfKTwMqsxk67UoYu+hAuUCjuM/62ikXKy
yyO01zjs97w8z3btLG4N4abKRA+YC1Jty4UfuBP0cML6HV/ri4jeplh7EPOtuwkAIrxHo1I63moN
Ewp4iD72RMCeSysVu8riZvvsQUkSCwKCk/vWp6KGDOKsxDPqbkno9HB9jCRF5ux38WK1gBq7gT/J
p9aOxlnDHspgiuxv1LuJtVwEAreo+zMEBu1m5LNKv3ltp0aC0CkE74xFrOXzZHZTqtSEI7oqQkMZ
luoo3krdXd4A/FqbizX7meNeeNnqHkjT9K3gT5Lnqe5kcfSOCC8G1JtFVRaHP/qbiA/usmb5soy1
1i7fgCeokWlkqV1bRCN9SHeghbjtDPTyeov5WUt5Jlu6masPfxdnSQ00oKY2uTzTXYNZBGjTjhO2
JDOFkOj819ODLaE3D52UGoPYh/98LvmgFySPlyfYPcBfiZ3IEPieMyaqdk9kxU0YZHJMA4C2Snd2
8g0k2RNSmAPBbaM1N3eRMh52IzGOgc/AI7bL5tykkszNvSFpozSMxqFFVWBgiaWrBicaWPk7hIMH
74wemrw3W4q6tZwFw2V7bKi/+snw+otSvp2f1zvuesmPdsEsdvjNYJs+XIAZcSruBY4ZtDItmXdB
+nJ8jGa7wZN8v38qmDfqLxwAATlr3xDG1u75suppz4+IW1H0z7y7qbCErlCxrlRgth8qRM1u/0/M
/p8NTBeJJyKu571ZruTNhoKT10ZnDNka6ifOLHKnJsNBVmnr0l7K7ynu2gTnh4Q1js7YD8cEzj5K
BYx9OEXXjlJQeWVw6tzXs9rTKYYL67Tf9SP+PmvM7z7A2wfF7+2XMs8o3IfnbxfsvKUnyOOq5/K/
s8UuR+Vp6BS6My545rphanmmKGsIoIZT8Ss3YseZhjLfxhFF5bB+pVHqT9Xp1XlMkIPp/l3tBsrP
q1h2Q8bQcrDg7cEVSRtA5DJO9BOjcFgJIhdIAQZgYQPd8/oKdUA2YQU2R3aUp3a5MZ8ALGrxlCoH
H1h7UyRNO53ylPybKFRNizse4Fo4OjoB+y5VuKL5kFo4s4+Uk9tCForzks+urQSzr4gl8mDnjAtu
Df3P479FKz2nYKUaScQTJpnzt1EFYms6oojtoVbolxb5Pv/v3YKOH5ZUutNNwjpCcyw2h7xEeeT+
WciSf30Z54DJDmLI+eGmClCU93n3OgRjDqoA1Pr9qYJcY29clOuRWEBAErFpsyZEtlgCP6XvdO9m
dbjG0G2jA7+9i/K3mlPtGO0XjIVjEJDWyAFphny7TGhN4uSTeZQnsBHCycqJXcyYtNdHKMfRCrBT
nhSYXSu5Fl1KgsDuR8WO8Pcs7FwvCaWaxzBV0ZkYl/MCNwTnDFTqAAftpV1Ku/Ut1ZbpACGZoYf/
mQ+kf4DVHsBPD7DUh9uQI9MyxGoguXelnOF9wtEEDXONRvgUpCpTSAdQJ96e1zmScOjGg1X4F/7H
c2jA2JKunoU5LfRlbN7ANgy3CKQhp/xugwDaD9yr2ALtYhoYHhtbpOgGniUhly+yJhalMWFfKfdA
JpPtkCwMN5O+8bAHeR5MRnGSje/hs3QBUq8JRbnnnmQMVCuXMnGgmhyiG8Aw3TNhmh/XDVUjM6Dp
/3GzBEc+JmV94MuvIImEtFCAn8iS7/sbOIBDmVsuzbSTsBCS28eL4IxRh+i1AoQcQk+4wNf4pe3c
hwXhy+aDgtmKoEjslS1VjlvZlBMWV40R6sGpUBVc9wd9AgKce7Eq1nDPbbAiOSG650swWxCwzMZT
gGlmd6qRY/S6WjFvPvTOZTgPdYTpOs/+if4MVoKgyXhDNCDIGIM98KGrGghTWiUkQD9VicWgfjZu
As/MlIDRx89X683oeP7Q0U0K/lazuWkdwGzi2nbTNB2oJ5jTPSXLCwI+i175//lqsK88hBbhsSMd
RYA3GNPgFTwRJuKoNCBZFve5mImcHybfMW97APmirfFjdBeXTZ3LJg4Z5L18d4o2+/4jH262vtJU
FaAJoRgUj2gVJs8Ydqf71hKOekF5MTx5AjwZBH0jM+F/1ATrvkh+XCYmlMHYVCxGwAPBhYND9X4/
C1gouW7AWgOTWdAjJHXUJrLCKdfayttI3JC15bmo3KpsW/Pr+jBmi8HCGKiqel15knt9i4eAAl/V
ceyEwBccGOGtPs2YHBOf/ly1ATPNxtYecfy0aFz1J0Mp4uRxEtmPIObpG07g20Pa2pn2gyrJay53
P8rKloI1LmIhRUkUSbl+jNhHoTmaOLFahXJmidQK+0hmkPzyNwAJyrlZCalii2Wv6/BLgZD4sLxO
Sz8zp9qYTVA1pThsdRb0fELxuqw1K9EMqaegW+o/AtjvPZNqPm9Rycfq0wqaQAtFQ0GvJO9StfgP
Y5W3E2VsOaaUJ9zO6tDuV1fkjRtZkeC4wHk+IY4UM6GN7r2pnDQg9VsS7T99KYHyqOSGsAHhL24C
h9KLGi17xjCpaL9DP7VZnMyXL+drWvqmvWKreKf7SNoNFKpWqdzlHYST/0BW4uKcEfRpVPnAzAZ8
sAw78pDbxhivVvnES+O72sbyXgVL+KYBWA4w5IEAp9PQJ7QH0P/H6actvJahpqUJ5DFO12s633ji
Oznmqh186E37tO6k55K3zy61DcQc/qijNd4Z7AI0BFodRdRu3+OeV+NLLo7jDpEPkum8CUIUU0Xl
6WL+s1QmD1Sxo4O6BRVvf20Y458CN70jQ9TFDozs8G+pB5q4L5vtal69J5+3kIf+7LAhDRNDio8e
F8cqaEQ3INm0np45lvP3uby5X9/2fVfV1/7fUkHp4VApa97K7CpsLG/AbU8C57d9dXtBU4BXcSpZ
iKn4PL0FKxtV1NOeNZ0vqNjeOWaw7fr/LXEwdsB+18Od5j7eScDPjUjWoNccYYFzbw2yns/7VB/S
rs8kL/8HnV0Ox5QPAushQxzfs1JzzHJkPHBXimk5QvUTUPvMTCDRmQuPeckCAk8c9236b4RdeqVr
k/TgBhtFihB9fBl6kh2EAW8oYP5jiL7WjX7BQB9cdPQbXky0f3WTKhg3X0jgmB0kApJqEVYdXn8j
9YJZSVOiruvGa9oROgPhHIdO8qIneF0inRVLeiHaWIDc+LAvgbJWRYO7bkDCgt7+yac6k0XHh76O
eq65+4fQp4SyP6Wjyn/k3+VRiC1b89zAp6z5+W+glyRgijkk/XfZCo6Y+rUPmfCkUQusRNuV5PE6
JQ5j0B4PGlVBey+ELo5estnielS7oZaSa/1SgKmA+GqY5MNCGHzFqJ/T5OVtAyiJdxnFH4tCggMu
aci2njBX2GOt+TS/ky/dLqTa/PSzZ7aDjylnh8lt3ENTKr3T0l6yitR0pnn8kxcZ5eMr+mRe2XJ0
y8Pb8kNxmXhpUdHdLEc8odSfX3zu7zfxhX+Y3oiGTDkrzUiiD37gYAO8yBxXgUho6UwyLHq5i/1O
2YWcZxC1NoN6SZRLR8v80aqUtKLetJeHNqef8MaKAJysYLWBnKJ8j//JodUUusW8WB5twf1hGkIs
snHrcVQrkDNvYjvqEkkKgIVCbzuv0ABq7YgXoJC6v9MFVjxdk4xDK/S2z7N1mUIhxovp4nCl9ey+
4BF5Ht8QcuWIVPWlfMRGtA2a4TNTzw668rEKrT5/Pv+xSurXufD2fUv2MZvjvFojRMAGJEkhGJL2
B/YtgcvpwNTNuUeFhcceJbT5zpwmO/B1d3ox4yytpAq3SEckSKEaSqeDk4O1qeOV8IuiVkk1b+A1
ja3uTWOLeFZPhdZ84aux/eS9n3Bwq7lOG+70HXU7doEWqx6YD2jT8TJBotHm+RJKvs+EKFotSmZc
EOuEs4ZwpURDbf88hjpi/eiNpBDEPKtBDPU8FZJ9F2hT00ESzcuT4mhFmVjZfF8v+D7/CmaCoer2
hG8XBLMZX1DL/BOjPhTgQBfOZ7ZAyOu5k85hwJMQ+/edjDdA8cgXeFcjcKXljG6uRE7gbYpPMQJx
zgy4ESZ2RhWsytXCjSnMoKmnkitMUVTriYckul5hAOtygY38e69z/Br4gfF4OxvRFk9aEek3WtNo
08e9qtEfC0mI/mS65J151UJzi+YbGJndp4jSjYhM0wdnzNR0kLKtBermRrWBGcyTDGinlSKMM952
ZNtlOwxYO4yoQT+7JTJZFQXVuCw3ODqteZeJMZuo2iKYnLnGTbuaTmTj7IFMa4XhwKBVOMzSGM2p
k5xMV1RIGrJ6gB3Y/XTK+WTsXEsZyTkxjJw2QKccmpBjxcl6R12uaQLrHAkhBy4TOUNLnJGv5XCA
t7Pv6HzLDnC99pDe0QvEXhaz9gWAlKT9WYwMljoVXB8dU5z44ZwVih/XhgZv14kTPMXLycOqNYX5
rhk2LB3BExCyxe4pI9iGnaAWPlO6YK88HBm/D8QG2uQE0iklbvVYTxwphgGTCrU74+AxcJ7VU24p
su5s9NbCmOUJcAC9nYQVWxSaxL/RzMyD2UFn2W9hw+GMMih++CuVOoAKEiSDKvS92N4+wf3+MbHa
Z0dFUgnoo/Zie1MmqWvQBKfJmjer8iJBGWck2kPAALsnXzROTO/S1B77c0ZCnr0WJ7/SwQVStraw
4+aCHMq/ULx72jN2qcjNJ5b4jkr0JEHRqMZXBCJO2Fjpbvk3wrvP5MAfxS2xnK6WTQK3Xw+SVdnn
u2rcYOAvqGGKlT8xkDDgcSJ5j0wWzxdYKx5qHSppIo4QrSY7Dqe81uLi7/HwXCgYpzKxtg+a2IXA
PB9T02scF8KDBMurRHhhF7YC5GXLAUs64laDBnuNeDgzd2QxuklmXbkjogJGdO3TkQrwJiTgQ2it
ozGY7IW3rHzPo9RHCgBWO1XwSCiPU4dNJOXE4M5CRP/N6CkWs85Z6rmI/+Q5Xcf/S5yGNkQ1cIgj
ybr4bdGgfHAozvTLJvridUYoN6FsCEx5ILwczO2tYs0R0RoQNUzjtA2REQAEQwfMWwdJ8M2K89d4
iLeFdzCETdIT5i/cJZx3XUNM8W6OahlnO7t30TT7hwHCLHIPTgqL2RvvoJ03KzpfSrz2ycDvjfpN
hcwcNDSiC21WGYqAog9TKTTzaK1atg+VQI2RdV05lP4tEEij1H/A33oIwxOrhY14qd3cbX3wZezC
Me3fTz3/zdBS22chF063W58zoLGCsMpyqlFep8+RitaNVxbx9SsRru4a3W9YMS6eBqrAQyH0K1oa
nRyWxSdf6+5kAaa6+ElRCJsWMU8SKSdksLwFciKOA7JgGwx0cIapT5PIlCG821Bk5lkXpVyO4EAS
1Wemu5QU1rdBuMiHs/mGlcnEkeLcWb+bEZKbTUBzRjVBxUWg/FSkX9joiJp3C97NsVRHuBADNfWG
G8SoDt/X1ErV5wPZHun9qwkk+d8loFjEk5RiU2pnA8tbb1VqvUVu5ev1KRsQSluu+4sU2x62p/WX
80u8RqBDj9csyBotzTqUENGeQE8QV+uKNkktFosf3Hdv2h8kEO0XYqO3I2Vvxh6RM8sbuS6bbNkd
BUXPHjEchEThpe33HjyRR/2haB3jIWplBJH/94fSVmFV/TCcSKdsmi3WQdO+I0Y07F90ndTBaCY0
KRs24BQnxTdSLOkylNHmTpejjBfOmc76SUW631vpSUfKv1I/PemlRwzZXxpiswOGjVKqJJAJegll
Lo1Eg4PpA5HNnw81nJQyIUx8WljB/GfKOK5s/XVMze26UlZQBe6kGq22EbABtfIfHw1uiHhXLsC4
e/NTdB3w8EvRp93PNZ4jOHh7Zu4M9zicCjC6i+pYUfjxmAk1MSY9qIDPZHheyX3zrVj4G2OA8vXo
zbEb39JJN0M1FFcrRLzG2VoUtNIawZfG2Ue/C3AlhUrKXohK0Sj0Q1KSYnVlB5Jae5GCnCzGtJ0f
0zE+jNZEcRPg+c+6CGoDeWHjZ0VMjehCTo34eRn8Mekx+OJy097EnlwJgtcNrxgE0/WD/CiVU+v2
KyHa4jjn7XUhBcrWW5sW9BBl6rZ34W10rgOXUNTJoYw3q8gxvM4Qj8F+mKB8c6Yy+Zw4eze4zS/z
HntvxHC2ROhjXj2+5GudIwPm1Gn50xhHpFUxQ51qFcXulGz6US9DErgG05oCbqY0lAw+bBjYDm8k
i3TuksAZSHYoORwF6koNjQGAzNTP+rwGUAlymcrsFeK7RjQ0sseWcybU4HMZUzUzoQuD5Nkys3YQ
ALFqGM/uFXQpMjptSQSbPPGXcY3ontEhIzy+XXxQ7b423q0lKEkn/c6GL79vhkXqHU9fMsNEqHFt
dWJ2D27fCGECBwIWw3WuT87gWvnudjob6LVVHidrP7sXlZ3tPLmkQ3pcdbaPj6ufqslrCH32PnBQ
2MxNtDGoLhmrtiMXUZ9UPlMli7AvSmHARLMcKkiXey00iljWZNHbPU8hDoLzS5oJE2BuzWT4sYG8
XOvTINI924PxJMKMvdlMkBQpbCnpu2/AqH/AKRN6GntbsGUKRZBFCv/MECNCP0iF8n99mNIBp8gY
WfuCnS+z1lIZ61UxuUudMfVzMFTHrHmTDHUECw1MlfzZHZ8uVG/TxZhDcjsug+PVa7RzA8hBRWmL
Ds3x8/FB2LYwKQ+U4dxo5J46DS0EBqIqMB39SR0Qpb1VSg2fNWh6Z/RPOADXMa/LB316XcLN3/bW
ki4b4ObBg3bHaKYV1kJv1U45s/kV5uaMI4mh1i+E2c1mwDVSr+Q4H9CW3/Si6oHxfhzq+ph9q9qx
9kt/n8h6gHrSopp4Mloc4lChTnSXtnQOnxcWyFlW5D8/0s7wAIcT0EpIA37WQKiPNawZ/wVPHG1o
/yZoP00IqvGm1k3MXLAirlZCun/+ZXDTDUWQnnvnoraXaenE2Jxgsmk1IRYgPdmJ9fxkdyVs4jl9
V0aDejTkFe0cJy08ji+hzJA1wdAmeNs4nDxUHMSytF4MZqRVEkVxTUpNPvJI44k8NIfnNnyCgXyl
MVclX9eQJZsdBuM+rSE4aBW8s2ZYmq0rsrIWB5tFOdsXEpkBZDXqyuYRhIJ8oHea6AyQc7UdanOz
fGjb8jsKTO+oJoFMNAlWHtYQkPy29YJKlicc3yQXXeuqzkkn7IXiBIbpB8fFFbZDbB+qkaMBzVJY
SJHrJr+pmCc2Rta22IP0ZIQxFZb8ghVmkQcJB52Ald3O2YoFysN1Mz4cr4MDj+U2pEyQ+FvdyEgt
gw/4zixL+DODcoyxP35x/zAFRWe68culVhwm7dXXrf83TCWz8aQ+fAA7GAEZRaLGCIMLjJNDvsJI
BKj7LDfLdSc+2EV0pwDkG8xiJuhzzfvJszHYlMTNNYu/gXCI1asIQwRr5Q+rR90hF6CZg4axN1Ou
R1NmoDOs3IFIZKgdlLaU+DFLDFzGDovgU02aIGS03/YiGH6F7972I3jlkkvRz+kRpXC9aFVXUZoC
mcb6kPqBXtIMxZC+qoG+vjI1L6uBw1CDWJCEUq+sWiH146mGVJDUw2lTYwNo0I6/NyBx4+iM2XBH
IcrjD8gCKMIW4HARcgr6plaYq0gBmParPhWQdW07oOQbHctUu/YkFyBTU3o2G4qxi5mvn2hoX7mA
NMGIsSDjtLT16sTYoXPg9dAKH6h7MRf9SFaeYbzL+gxjM/arZ7oI51jsKBdxkdXY35VFar+cz50x
fcP9OO8UJ83wo4wwg1e/yhPxrJ2sbgfAWJnYloncW+HQpx0cqXFkwLuQXfgbV1J1ZdJeKpT4TCDX
AZjJhE5zD4pg8BnbZ6bnBn/Bi5wAuFsXrbaEICB1xJvX0qHr0OoA9Pz8gt1kGyvIZeyFTQ7+P2zx
w7ch/qBTv7f1lT40qwzsx14GmQnayP2kyL6mHOUKqfTxtnhpZOSb+2Ay/P3TnXl6nK8aXkTdYIPl
iIGBJqCrt7TnQoUnTd41k/fP+CTcmXSVt736hhLfnPRLpkLZw26a3MjOFl/BJHCr8WqJUAsf7cA0
xMK5fK5RXNHpIK6aqieOeo8cRZ6RKeLsFXsFarCvSOhTXBdNFiSACsyWl89LQSdAi9eemQrnsUON
fZyFeSFhVo9W0irieNQaSv81qKGwzglqPMGnockd4xBENhLbGIcNYlHxL8mBxbk3yTVrT0gN8JF9
BjUYj0PrnpXhQ+Y9E2eezmcqIvV3Oqsq5dkE62rbPKc0NmVbaF/aLxdG/vgq8uDjb/0eYDN1yAxQ
ZKbH+4OZOZGx2uPFDC2pyd66Jw6zl/czejRXptMJ5sv7My4WnstQOGmxsM+urXCPjuM+hZd1I38S
xfa4JnA4wz5AnFlX1u1r58C8dHJQjD70v1vFoLNCCBVULe6MJs/EAIBWjP0hm/TCUj6xa1vel8YF
jWehxXlYG8HKEHnr0r+jGYp+97xFvLikVEz7nHN7+En91BzuS8NCC5O5eVZ+xutZyigeSX1EgDid
FSaEkG7RyFlbUSvpSbEtaEaFVKvfipWao8dyQmy1A+JjGYqPnnUWFNkXeWeI1XrEX7ctwasZstDf
Fk3SLyV6HdWudA/pRao1rYp/M2Rr8llycaosYQVEEjgsH2xcuG6TMY30j9+Hp7pqNvW/vKB77rtA
PbqC6g8h2tvg1h5XK4gXd+NlA2yoeS4bOhGLlk5RUCR/xa9PqpXfF5qXvqDyDc8QTxwXSJgWpjlA
3G1fJO2k0xOAkGqmRST9+Pcoz4s8WrolJsjX0zvzPfF8ApBv+I3X4NY3/x44UwsfjI/xHavkaHlJ
q77qcrAwZg4nYfSPXWXjlCmgUZ3rCwc0hwa/duRvZffLYhyj5Lz6svFvXfRGxFVDhAqcZRaP4q0a
vuW0N9qBJe27mCU0qdsmNfOfWC1JglIKAubJtEdsftLTD+azyrx7NANiuSTS4h7OXFujX6WoC8Pd
2NA9WLOp/vt3cWz35huUuoCq+1IDTbFHakkol6jZhq6mN1I4rG0vaoi+Xu0p8XZ2faXTNcNu6lQ6
Th4/d4lGMFh88iEFbQsZ+qT2l2EqVnpZdcsUF8ekqz+wZICnmPooqb3GCnhvourepUiUGasVse9w
tB6oE7hyJDqnrB3I5kPK2NoSaWvfYe7PZV1LKNW0Vt/aJ48Iqrpqy/L3CHTp5x5Fv9wiejHLz1A4
OLclK+R3ir/mbVHeSGew+1SuBSGrJg3qsNz60mVq/H9gYJ+49F4q9C7Mo++zHOi07q1ej/x9t/Wc
Lj/wk+BXGg4incVcH9HSp17ys1FcsB4bW3XXtJi9W0VN5zXiePJnVbcFK6sgYSltnp1S3LTmrJzN
S8hMLr9pf1J9KoP5OGb/kcFmI37MD+fZdbzCssmPkdRQx+ZRxRT4TQ6xJG7f953b7uufUy4K+AAl
bwQAvZMMjW2eXs8yd4kVEjH0uoMKlGyjxYDZFeuJ1OVGboFxkMB4vHHLVW1z66Ki1jqh6x1fPK0O
VFrr7aEddBYtkEjHoCHrGnbjpKdXBNKQqArhxzMbaDuJjyhjZtgI/4n32+WknqVEQj2Zrw8GgRxA
+tehAyC1OXgKqKjWmHvh09kCI81WVjPsM/9z0tcVHQU4LGTTqfERUFPXPPWq+6bhoAPYaJ5KzsS6
iSIJh8Mv3Isz7NWcszFiPGgeIiXg/bn/q+d3aIzUa46NLlwtR6LoImm3rqtLbWJH88TLCsuho7Vo
qKm2zit4+QBKzPXLlUyGgS5NUEqMIxtUSAH6d7ARQN596IA3Sj3RXgx807iBChJcupQtNHLFsL4v
8GXoTrEz5hW/a1/H2oY7Uhj0xUfjGLoq4CCvKwQqwYpg0Ky61rZcfFxftGQDB//QPz5Ijsme+pMd
tg+LP53/2OjNxZZv8q/ZVXtILBjGeZeFJvyhvqK0nf9xgCaj3rw4epwBdJnxEjwA2iXqLe32bihk
9QusWBY3wI048RlowVx7gLTdXe2QpJbeUDmnZK/od7f/1BcztXJgrz972B9Wu3qWMQkuT5PDMS8X
qd8CHgJASf2f3Ace21kDVM95oaKe2mKi43yBTHQeGtnajlLMHiFnTwG3mAX15GNOVG1auk/fr6kh
R6739WJf1pZbG7Zs1lWV03ySxZVrDrZUlGIHJPIpCCRKWvKFH30PPwrCk3U9n2lWi63MA/GyNek0
28gloNRiByxsec66y0izpAjv2bQCNxdPLP64AS94QFdT4pv4fEbWhxiHW6RBG0MJFHiw35Z6+4JD
b/yKgcP81mg3QWa4hOMBkDYLA+OXgBl70etOLIVl+ptmbXvzcjRCSzIleCBEkYuQjP6Pq30W0872
Urh9GxdNO/sn2TmMq97Gz1LYTJ/QsLiwZf95wLSBEUgisTsvwAh3TUvYK5paCIf3A1T+WoLbTIe4
ZRQ9iZ30mUEzbtbjiZHsxR4KR86nsCfctDT6nwX1nHgogH+zkXaXHU20eeR0UlmL6hBvmxNE0r9F
Y9+GgW/m8hhiOsuIy3L6ovzdfVTq4mvBOeaAGblhjofnjVLL+QxLbaVbaE47D5x3K2Oztm7WlGII
E/Fkey44rGaCgMZOk8pn/P4cfCzASvPuaJVB/A7hjGEFhr5jHDUbm2VulyomIluPwy3GK5KQwnbN
7wBcOdYAZerpLiJM+qSk6Ng4nRUUOCCpSH7jEAMtf/HZo6pOHasPjqTCDPPPkeTL7FUdskSEqgQE
2gen91TFolxE1viq8kBG+WimgWwuQtYN4ozvb3EyNVeRDw/eBnNjV1mEvJUxbP0T7qdKnc95fhGe
Nzzdq4GqapVLeSMrOqfjGoQjdPtKJYMonBbPQQ/RQOVJUJI1sysY/8RYyJMJvsD0qkv8GLHXARXs
19X/fM4qxw7mQ7V69c3vgQ/Z/gTByamAdH5yTHXB3IAlJsPW7euiN84K1IQOTf2t2G+nIfoWRr/c
9jdUxR9xYAj/raRRMtsOdEnwptzPmtCQtIK2cHT8U4EsPj9oj4V8Y9KvMQ5d3okw53HRzm+AU3No
+8SN1G6t+5coJ5pkEi+Zsm5SoL3tBKnz0ZWPxBitu+8eSrYeBjGTMfpl+srftIQP4HUdKknp9oiE
PPnHEKcQ8aAbGpmQGFPqbLwgQvEiv+l8lOeZ0tIZ2sZW4ZBGO/h2BvcDZI9NTWL0bnmg0DXWDsNC
4cG5NFvJlBP6mTOYUHuo0WzS1FrxW7DHP2QxRLOPOF05ISC8nVfME0N935inP7rj3U3up9e1/Cxv
3ydvYzEWoU2zdXlO22x5jobWP8IoSSkRTtuUKwmX+kCurvS/1V5M1aP5ggUCm9VIjtEq1afHH5E8
Dorq7VkCHXA1+dOGGsxPyYO/w7qsmOtasmXqVKhp1Bv82ECqH2lChTPBi5lKGozUP6SgDuF+f8z8
0P/OR6F0EVa3kvSkpyJfH7V7xdTbmQ35aZ0drVaH/4GfWuIwO3gOmDNK/uhGHBZljYWr+YGjAyKx
iLuMOEIdoCdwZ4I7ae4DIads4B5sw70FUgWrCcDaANqyWcyTWimDnE43m1tsoW5AETgzrKPu13zB
48dPktIqzH46MmxvjbUFn0mqREgaXXukYPwQJ6fm2ZrI8zsCVDzpjFwidgnH05cZPlAUB1TZryRI
pRQ70EDONj2Pb+U2tnXcDyXTeYj9oGtvBfTuwJBMzY98nniTcMrEcZL3YWF9MWk7sfhXSSHTy96l
AfVPcGmK0IF8ff04BbOGOlE2rRumIi5vp+Fmf+RckRejJPB4alccgYoflcSdziA4S9yY7SkDodDz
KJ8/b5x4TJ/+bmuVD6TyvHRA+7tpW1ZZJTpU7WseswO3gT69Y8+VGsWNke3PMXrFvXg4vRsSQ+T7
LCi/ZeZLSQxoX4P6Iz2S5Cve8cYzhvqwg7fAWE6ao21te73SKlMAM1aPXfoLt5ZeplF5HIRXt6Td
lEP+4hjS0oLfKA5ZNul6bOGF4HFQX2EE9yAA4YlAiv12cK4KZvsPAddvpLv4vSdycRgqClBH3R0B
AQr5e891twgff0Xwh3ROiMHd5cMmsThPebGR8zPpufp6EHH6Ul0yKiWwDYcghjAwOTOzI2Y8gFQD
WYEitT4wwwcfd8nAONf+8pEKBJLPHdJGWn/R2Apg3BezP6l8ir1nNFTDD2W8p4UZpoPBlPxHir9T
gJtsf2oA+zmt9SPwZPE5+vm/gEFwcaV3RCOo7FlUzWWeClKozMZPK4b3s3sP5Ja2CoQMOAEUnroX
opSjzRr94EdAqfl6wkJ5kzBUIHiO/APAbx8In9u/7qFsXCxsWVJlJZOKWhgHA1iC/1vAo3y+O/64
r26k8ysoEHdtGQmPAj0N+jyQBdYxcvhc6orwOIFl/gz2gyTmdI9nPhrwlZuscBNkv3vEwtJ+kk9m
guF7i4E6QNild2HkBsukFmEUjxiOhvOEsOkW4SEabzWXIt/cZYTlM6sbS0swuadDGfjijUdghgW6
3HzT8fzdMmC2Qup/OxavzFgr8sNQ8gboEeAUBXw7pya5P6k+sHGjCj3I75jcHae3Jm4R/Yow34YY
mpp7rnyLYNsKfdOVY9PNKexw91GWvI69Z0KaUic3iCK4ubhbHi52c5dKxL7Gx4qJQ60nqMIdot+r
KcjEGFCQke7SPMlVUKMxvTcDHTMfI2XR8Wftys3mXM5YWcaa2lq3+wN9RCX8RMs8PmZwfDSozvmn
fFa/zBgSxZhCX5ttkjFCuf/JdMoT7snXdSRl5aTFTJQSy6hDk+CNnrchEXz+i0OM9pUNlGwb6JFQ
JISKqoume8SxlsikqSPxDOAENK+zf5dWJuAM3/LnY+FN8yzmJX4oigTt9qZrWaXQRdzeLikV4uJf
9dH5gNGWemTXCrXGVOzDX8tV3FtxKuQIjZBWCShkPKh7EnhxGO3Vr2D4f7Ua7T38nH4mSviFYG9k
5x5FEqhTe3TjfzGttlKW3W9FCHZGnj1gxn//TsxTjHfMFv2PipFoBUn7/x0TPG/Zw74niK/nmupL
F9wID3U3iRxqyGRyAdkPVEY6mcq3C1BtcEcaZfcLrzfgGhY8yVwnzbMciI5p506us0gb24iSGCGL
ygmqi9sc4+fwcV4RpHNUIYfCiGi0JbiQUHZf6YjpSB0MQRjtCGtY49qlbT2P+RIDg7HYEqEOMw2X
kLH6VmFMKYECYN4XURDXoXVrrqohZT0AHtKpKaWB5CLEi8fNEtBhDURxB9EM20r3CepSb/S9p8Kn
GW4yuSckHX52OeWt2JwFS8VSssoq/6pH9EYocfuEu+POt0hAIslK0mahlbMNu9bfbUq7N/v/Cy6A
Cy+eL9w0w8tlHIUMqaYd9JcYcqqlDv4lOYCggED+vOqcWT7New/kL0gvfgw9/RHjdOocfY++FJi7
iRkDLbVcAR3Dz8WuRnLO/b5lGgCDIyVR6XhZxj1AQ1uk1OKs9M9/uK6MddqspA9fN1JdNrwCgyif
EPtxZwVwLrs0nJoSMb0C/pROMXn04B6yv2crFEj/AvoflXCIRpQsciRXqYdySQhx3riosDVXv7uj
2JLFKPTE0tm95SUHEaqP4YZLgWvGcyTSqLvzjQ9byIwfdlc4uU5JLUJwkOG35PE7XIoMRZyROAsf
Oi581Vmy+hF5QgucH8p6OvIIxdUxbV2sixqX60Szlp75m+1qHcjQNLoE0Jpdeu32mUiGaYr0lZwB
L2Z4wyTHhnU5xoGFlhYTW8O45ZcBhqu1wR9JBWDYqBd21BhLv5DgHBpjfOzY5TXbZJllv5NT3sOd
UyfK/r6Ks+M945xWwN5/S63XY5v4IVpMRQ4v80rjk/xmW1yVsWroZ3MD99Pm9vLgyJnQqwD/ifoY
3uZ8jkG2O/5mOBSrvgIxei4ygQwbGUHWtPLZSoFEG511XRry7l4jehCcjd8aCkdgknvUZ91dnyh2
du0A67Ycg07PzQcjP0f5jEtM7OICeSDypzuHjpSLjKCGdOwG5xf5oHIHynCpKhl105CQPuu6UUNC
Uo5LmsLt/fNkvULsUOqOPqaV7Q+drwlBJpFzirV42JfjhGqmT3kqRz2YEjNwWwHVua9qzBgB2zeb
2YePVwV36vVzWHIfo1nOR6Dbnn9G8a/XwY8+8bCJwRHYLyEuMZ/OlpioDlomIqfIvcn53Jy3ojAs
ftXbxVxsZWbJxu7D6uX+ex5iaUnAF4dJcW2/z0gsmBjNHnyLUscZmltQWzX04LQ3Ba2W+tpwkRMQ
nhxaq9rq6YILzUS/uAOjsEjG6GZdObSSZRLtwJ7C3jFvmzUisETmUfDR53xBe9FR0dj3NMivn5kQ
qt1r+Tpy38bWgYpRhEw4bX0TCNUB0YqmFhao81dmmGhbr8QOR9asd44ZwZhIHQ3EsfP2TVDGRhTB
5eRgtiCGcjiaO+y2NwCYkaZ/3uuLjwkQ3o1gaMhQz08K7QT3BWsn6o/ADI8GYngoukrfPJNihnQJ
X01UyKWGiNUZ9xrdDMpsCInyZq7g9CEd/Av8xwfwXLe5TK24ZlxMlNlIpuY3cBmtw3qCHLA+jwwP
nstAkrvuJ3STmVl6YCUODAqi22HczKqR/YYdvgg4RwHl8iGyWL2+yQe5l7x6oXmDMdD7FdH5u6Nq
vOIMl75YEH4U/hL8/7bXqLmD4x/0M5mslF8Ql8KAOHtmQg7GdbmEk7n3WQntQSjTMsaEcNhE80O5
/3TJ640s+d9Q/kGys+6AfHATVtW9xoleBqqd5F+oDx8Y8lQ/S3lb0/tIAOjeUNUrKtulQ9VYiktF
vDp397S876L0Xu5nzKGRqDhPPm6WNIkp7rb69Cl95K01gLeVo3I5kXYtbfQdGwtwc4kLWHzWO6Qi
yAWjtxSkgcop3AK+H2GAAEvbzirPCOgIjpxN3s/tYU+FVUsWGbRIlLriN7aub9vsSrNd7+OGwS9+
gX7zTgQiNFEXKJni2j9RCKiZ0/qxfOv0I5N6o4YkT3Ivy3ZA9oJeAE402S4lVQXfpI4FJRZ9ciiH
NHiwWW+7dknrxfOOOP94gWQHzbrtpsuUUSB1eMsYz1f8wFgWYzxGPP0MgKAm5RyiPd/ThUMNT98z
Cqbh0aPsw5bSC4lcXe7XwOx096ZGXo4GwZKijtQMmGF9BfCP2fdegZNLNb0HAYQO9XV1zLU2sxTO
o3BV8Kz2gNKUO+SziI8QKX/biPRa54RZJtneyDrykcImeuGKbgRoRUJVH72atyhN14t3TLJFACPw
YJ96jJAQfcFPhkdyMm0O9x9uCqzA+EEqkhs+b4Oetuh/4JPiHf1HfJoW8Jk9Ht+8NQtc03JXy3Z0
KKSg3HwuMTJ/85BVKU8WBMl/QLOF8uIY62B6EDkyfYFfKW7bMzKsJ8fYBPipe88PTA6eA7C810Uy
7Gz5Qd6imiUSMofEX5qHyD/uj+CPtP5h7IfEpOpOFmYdudoAmZbQFg3sCVsx9N5AMBpmVNvxnneo
R2MR9pDHBW0JgQQwqCQOm/SLHmkpB1/Y5OvDQcEQ0TdEN5bnLFzHgCzQjkpNvcJ6M9FPvGl+c34V
CWi7ZjexsMjpOdJnpaZWmGX7fkiqB1po2PKOhvBsr308GCHACvszX4Y/tAkkvFq3hIA8zZi33foF
dL1EgZ1GOsBrkjICDgEKOjTWfPdrgQ9UOmx3PrrJUKlBX28fJNyhysJZsZa6vRw2z5rK6g27dcBv
1YuHoFbEcKS4A6+r+pyNUXmrGGW70KRp8xYhfuZHNtysia53ROvgBxxhHb68ixF3wPSUz08TqXIM
WJurpXlkXcqHvoCv06+j7qp27R0V3xb0Wiee/2VZxHS+e7fmXnhbMxeAId1nXWGoawx0B9B8sPRn
lX10cy1x1UrmsKLFUPrKCnecFK5GOFmgy9SdRkiiUFRXOx+6v97V0FVQ37TYLf1FxdY7j9r3tqEd
M7GiLucSuzOR86KpNKUmaXU3K4l4Xmiqrk61nb6GbwbnykHlp6cXf7Jqd9IbTMCPitioVBfv0Sn5
UnctW9WfIu6vvxuYMDt0UKenji2qXmVQ1YEHdVagpEirZJdkYhDAygwg/OPUjinuCxggRBRfqFAt
/K+EGaNz6m4XJ5FbgGP1GWNbaJ7WNVAeqN2QxKPdX82AjECCSmQAEESgl8tLdQxwJiZZG8i8ftpr
CzvH6G4NckdfD6M2Y9CChry/XjzxoAc2L3Z5SAv+rfhL29aCnECC9vZAaHvhNVNwIsP+psSbvUJs
a/gfDurpf2vEJQ1SP1NaljBBQEp9uiM+CA0r38KfoOYNHeRcYc1F1O8yEHhJygVEaHCGXrXGMlcF
619duZuanyYPRilDE2IctqsR69aXQqmd0RxDAhFW1ESDJkTQcbVTR6vmGtFsqf8zFA8utXk7KYKC
kdhchepiYODVtDx8oJA/82O/T/mSuuv6sZ0kO92pt6eHMNu+cUdHa5vuZKiisoyXjHyoUj30/RBQ
6ltVOl9DzcJhOOAjCqi/i0t8a73QuPtQ3qOWhWjgNaKvFUi0tA15hm5ILybu4ELhVr7eXBGOjAAQ
rYGsaAK4L555D0sTA0/PT9QCS1zVrY7Gc+SNksAebFbzpl2qA0JrK5QFqdmaw4kBVKwWVlmGC5pj
HbWdsB5BSeyAZ7twN7yhSo40hse1I3hXPMuh3qi0SYepgwxyG55alj0VVps8h4eaGr+AxIRF/ypS
8gi5DACvdLlQ0W26vmJt6/j1Uf1VNoPvvlyqCf82sfQ8sddKQonC7yWLGH+gdLILqv1UumQqI711
BGYfsz99H1Zok6CIANESfKEVDI/cOmzA7CiSAUirPKYzB9tQ/QEdvfloTfFhbJcONSsLCHfU0dsI
PgW++fjSKHFPGAUhl4qCKeghJnTaLSaZO1DUArN8AROHK62ktjUrAIR/ftTMRLMhzlXts0+l5GWO
RK2JUHxFYS0ULxZo2DBbFHMrTnuL+EiPP1tyKOSlFigkviuII7JvFbB2ur8bIuT/9Lyr9G6teFc7
UwGx0LyHnq3n6hOmev+9FyK49AlU1P0H0vWz5eQwGuS23CU6u+/juoFNNVGQ6QMkOzqus6wezb1C
yFRlgmfdCv8qTfXhDisSW4P+SLs844xrUUscfi/fAphD8NDMOBP7ogefhxMEJDOErMgYNp4GWtSn
ElAbNKhTj5wFHNMk7DrUDMktl1ixjj1BJJ5/CdTt+SvPxRjtwwMUn+amB8Oz9r1IL9MwMKCkKkST
iNbfE2tWZU07M8spnHnI7WgVIHMfHyV2MT2vqI4OAx76jUVbliaDS/YPprH0zy1blhGQtEFFC8KT
dBUFHXlnaumcTe41Br/d3Hl12ue39NKXQigPgQ+62EOWIW+BfOf83HNwXgQ64OF5hNHnuJ73bIBb
B38Qci60QYnMDNQ6SdeVGHr+urp/SrMOvbrZxt1i+CFb7Y2ZYOMPjL2Zv4vG2f7C/g/1+A2fC/Ns
vZjG3o6t6RJHaIVMZbHkvdYtrdmxhFyfbwcfaAUDyxg2hUuhn/Uk5Oi2blsCldpXJ8ByaIwSLr/6
rGc88UtXlPuoSRvkbhR/UBUGVrEuNicSWd4YKvDGM9ye0VdWHWmpk5dRRF5AhdMq5Knyq7hcEIhH
Klbr4KZ9zNEQlluVy3TdhFAZEoxn1b30H4r8SqJ8KMQB2NQkRWyO9hF5PwIy4763tJbnJRewANA1
3y7C1nNSEh8nwDVGHmnPE8iI8I3pMuyyBaHEbaAJppinYSZ3R50QdUPOSRWy8PRqfS4h9fhjN30E
cNYYfPiVBtjxpTgvYLG4QQSKbZYVQ5SayoWjfe7DxIJ1/X7npcoDgda7hxtCKTz674cK07IoPvDr
39vpQXnUn5IwedPUes9o12wOv5+kzsa57OMCQ1Dd7954T2dlMMkLmDN7uTc44BmdkCNPl2slzx2h
lsqkY+XNaP73TxFlm4Q8GuvQGs73AniOLVDLs3SwzOHSoYuPT88OcOclTwuIKQTPmKTgZpKxUSek
3XgpAYnIV15eZb8SnE/PmSMMZjFpDV4ekgk4+eZjyiHD5n0TAGpymUnu7TEEVmLTvD0lboujOG5Y
zwqiAOsetLo021/51GbwVzaMRULb5RvxgCfJoudQ/CzfiuOM3EXjjtnTEM2pUjk8YXp3FHnP3Qp7
tYyQ9E7uZqxDFWiTFUfod5kzwmSw/BFwIV9MijjQPxhO14xo0zOgZncKS4ddwW7Mh63JoqT5OJsS
30VSRszrNQn8yXbF1p8gME7HPhyCmEwvIyAEXGwkhWf/NJhk/62wg7nfws1X5uY5GJUAb3748wyX
+npnXhChUFCEFV/8nWtG6+xvECDW+IoEIdavewl6oS7rsV/imJ3gXMysvg8zosuwF9GqrYJpvJ4w
Y7Vf645u9Oc53NdYQToD8zKqBBHRaBSFNKb8sLHHnkT+ctA3WoP7Uy+nBi6Ur8yWsR8mSh+mUSue
b3SLqqkdwEAhFDl/39BoUuTP6JRoTOOrlqSFXfLTkhbkfCQ+tDJHEHxYmmYlHnZhQFfxLZi7AY6M
d69/N/n3xudz8Acpau8WNKrgGGDdUw4bccGTrmuY7zLtOWGKtNLlfmv3Vv1RPjWCe9NPgQYNVBTT
CudVUTrmozNOeyI6UCCErAONFEQfrAbFH5OeBpdaE9ADHZUDrn4JpsxXDq6nuJQj0XNEFDktJpXS
8DKxqsu8GYOfyCjwfI++3Ohqf/gdwu3PWChXXvvQEWArLwX2vJ1B5of3dMI96ZUxgTv2UtCWsXIW
Z8E1TKxoH1GT6HmtfEdQ7kJpxRLzOGtCNYevZBBvJwqH6SBk/dY5cu/5CRXixL5fytadsgws8XcN
g4ncSW6Y2oJHzIDznqBgNUynAHxRy+ojauA9ke+LT8ZIxQK+M6FO/m/sLrLBVOiGmfcCaAT9M3Js
obnH+931XSlq400wS08NUlibk8x7zrOKXb/4oPocwW308udWzI3FPmLNGiVxNAsZxrWXP/CPr6gl
AuxzYDsm7BGXCISPpW5oG0tyXGqh8Wes+BE9GnEqQGEe9g6fYRURsCn4+YSpL/JfEVDGU+oVvNgu
fU9N/63E9pPvNv+ngz/Ph9iblTpViS4LyY3drgk+IH+JuiIp248O4hynUoAZkyBeigziQnYc1wdi
MlNqF8Fbp8aj3bIjSL4DfcC0eOkfeFJs58qAG2K3xtT7il8fvrKc9cn2KdLEvFLHhWNoK2DYW7RD
7falnrFtGqvrA5I+2L4ZgOVxYI4y4p7FC+SM0nCCMWydtqpGFMA1uNmxsNmCWptRnU4v6cqJZ25M
Euvdd93orzm5IOJ5g+jnDywDKWHSZtsrjY4dUdQ1DGh+zn8HT/aos6av0AiAHIlu+VJ9tHR4HVyb
3jOWnAufj0gkwJjMWoDbtiUkYQG6yuHr5H4Oxk8+7VQBQAhlK6mMNH2538ScEZ176Vvsbqo8JLS0
V4fbByCySwogDPgy459IfkrOoBzzz81dKw8wjGjaomsBXc6lpwwHfi+/bnCzqlJdyE49AaRe+dLF
2S0DHKNX2mVk2+Cc3DIIKBnl7ASus3caUSJIMp4ZEnZdgqLgZPAUTHcisyUdIK0etZbstslz1aSm
l8WGaimap5LGWrIcaHittAMD3s3vdNNJz2WIwblOsX+oCO09spMdw6KzA7m/GksE844mntGt3ISn
sM3sWdxYBQeFQEycmSrqQGt0iz20ys+lN1IdyCQYbTicFqHLUQJmmE2686JiyTyU9SpCnzAnB/AR
dn+k0KZ+8n+sSW74/Vvvr+5cJcAMMRbsYFa68ORMHx2oDx8BZQFNzOYTVOEmFgLTTez3YvACVlow
wxFppHL0PCNUXvkM8pefchw2Eu8oMQFHNjdUle5ITbi3w+uKvNUNgq3hc3sJkoaCFxJpnUIhLsQT
Z/LogwXMrAH5Nq2gmFwc1KILxAorALCNbFNqGCdMBeCUmc3jEH34xB0L0YbkCCR6MyCdY3qEgcvX
eZu1PZCzrVNqXYP96bcVE9KJhod1Ens2Maq1W8AhHWMZYYt9gwekDfYVX9aotmCuHINmyF6XnE85
5iB7atkiOpNJeu59UsnMsRETTNuztv/zh5oTLUgKjAOxH+wl+wboAKCCG6pB6Y23v7cU1wLxApP5
FQtmJ5Rn07haBDBsvSQ2Gwg4rXVZoQW3L74T4NvM7oLkb+1p8/t3YCHPb+GO0uiriGW8igZYhgr4
xC0BOb8FRZ6LqgGlB8ID29P3BL5WKV9iEWLe5Ehb5+3Dmn4VLayfTyMggjLifMSiqRnl08swt9CB
OgSZVHqwi7fnfF1jWRoLSbmNd5qYpdSG1VLrpGaiN0u77ezkVE/J9Szbv3sJjqGMLQhVkOTM6+DP
wkT2B1IGw7UKC/EdUtR9ZIbhxKTr3N93gXXJ2/wQ46ktNp6RcNtoz31eQQBAe/y2X/yLJb7flTwz
gXesl49Cff9SofhdumPzesPa6qC8L8k8M14Lmro2vhlJaDcDMn2AbhhmXuuWFbIqQY8iAy+NxHMp
Qysu+MiALG32Nlxt6VLv4sY/CBj4sOwxAGZphakA/8nj6x/atCQFqgJ6EAddRzwjCQJHuR82p17p
Kfv0DLvfsQZ5mltl1jBEHghGTvi4884BTJ/njAmci0YxbqUBm11Em7PY3YNyxdmS64K9nZ+BOy78
b1DioNx99pET57WWYb8O2LJQEnERWZw5EHbjWDvSDvb25kmkOU4hj9qg71wDIU15fFTZ2goy2Ilx
Yv/uP4kffkoqk8r/qsURkGX2+IwyKrWCHCg2tQmJHIEw6Ww/tkMVvguYcu1djsZdfBaPFzZkOB6H
/Pjvy3nQvuljmAPLLS84I1sJVZaFgF330Cn6Au1uviCrjkCT+XUK6pYoC7G4p7WcIhHT6Mu5skI4
4uLjjK9FAc+6qLaST5ycnjyl4DTUyxcgfrIYTi8uF02RcAjWnGe+mzMqwMGe+hXOixeL3/OOkbxO
aB3a/iKN4g/3kzOLDgIF5+Ac+jhX14lin9/8YDo+aPmEPTlotSE0QbcVWLi7Plgn1BxG737aep3/
2ZjY9kYTJ/NPt9u2upBXVl2OgJ9LfIxCo/vX8ofvrpxMaRTxSF5Ojf8HAjPVvxfquT2EkPmB8Jbv
gSsYjlbqqkad5yP1W3HQawfqmG3j+ozh0kqRUCrXLgRdIcnJpIqc7SXp8qIWLhG4QT4Q7SzVaIJ6
TAcBe7cP56cI2IvsJIu6my2nPUW0A8LtUQJbd/FC3sT8tusnoZt2WwqtnTeOEWfg6M2PGLpe5NEj
HDBVXzs1uHxInWN/EOZYgvchjCLE8KB2nHbBIWVtNzezR+1fHkrxjGYX3wF9/6hWNrPtI/JLtWfl
73HMKE+OPVJbfzlTWxiLPlOC+/FW+f9HS2CbszPFqkN8AsrkBmnPRty0n7Pz6OCW5sgF1MHVUqqE
fgv2nJ8xu4JhthVH1TAyaoDlGylC2zAhEOxjiKMhcQojxhD1pupij1FtB6rug5Ve8JMzhHilIpfY
J5VFDReW72McPa1Xjvf1rjsXHCkp0ySnco8OujCmRaZ7sEU4SIgKrZ/xcRMPdM8Ktp1P7prbqYVW
vXzwLGm8SWMdm0fe1nDnfMz1g7V2du20gkOpnKu5RXPOPF0LUxNMcJRty+vGaHQojAVWAucDM3Ye
moHei8DaBZBJPmKB59x7k1DLa4p3pHYy4uuJxNMlQ0En+mmNyMBJ3kF93iXi34kgM4mfwiKGsKdg
rXMWEuq300Pv0AXpN7aR0vu/SD7ik2vQe1/mMiK7V5NL+V5TzbM9AvshDSMh6hfHCWh7IRZp2dJv
ksHO/D26RW107Gp5P6Uh6+ITx7Fq2MjMtsLMVNDA4eEBmUjnMscnqrif7d0v2AA/tZHI7Pd5I7LM
EK6nuiK+8Ufd5K9P9MKwEbh6IcDNlPwdeNr6nPNBhSKqk9I+qRVeHu92tRZkDL3rlDksxdWlf7Yp
0qrnxwpYq2RZLsNT6IMT9VogdZnPd0jpi3KZDHT4AFQpV8LnNm/t3BmBlANiGD2mdnfVBQ33fnzT
WOaVvnfCKvUbdLkdQjJunqJwDdT89JqMvFbPHE2JmMld0VUET82YL3ArT4xsbMsBiMGQGSlfjEcX
xFC811ciGk40kl/yQZEURF7Hc4L1P2hD6ro4KtFI+6pmYzXqpNkdvTV9gWbaCfSXy+7zPux5C9G6
aewSp7ELqPsnyr69Nbuu3QDjgVUjMT6djsVJf/E7noVLEIMZ52g2OUdlzCgSCYu3gIl47H/PQM5F
PScN4S+Qi01NIPs+L/Y59F7ei5ppW9WdHQgrpU/pr8e3ok4ZWWgTBi0xTfIpDzsfYZua10E3NI3e
gFwoJenX7pw9U/o1SVMCr/wrZHFSot7/rn4WofGLqgmNLhAHAWhKtpXV6Mgt8jmKb4nJMTMyXaxA
wi1QnpKGFew+XlLip7ptSuWyc5QI3igbleAwsvTKo+VJ5RDOIAhYd3HbWmlJfc+nLrgmqytG6NB2
+re/6nblnuALzUS8ek5p0tjXvyhj0kg65S9PZV8PiK2J5RR9aexIP2sB7Q2BL+FNQetZbZdEftIw
uOOf1QbT/3fEYhTyxJz2SgldRFBcQLOJyhaL/dQikLJu+Nh55fjjt9I3Hh4bFlMLVNHcVW7wUvka
oEmQuhfloc2ThgmiaHNPVDMfktowPdV0/QE//NEs4w3s6/cX/lDsY9KBJ+NzyFBW88hhNRIX8GNZ
ybdQkWGdnsm5H3PW/E5v3HrenqX0+oEIhHGSVV7kjnTz7wtoNQ3NJJZIWZV4HT7GEChR1OFCXrKl
DLJli6wz5F/LyfnxdMCDs3j1F9VfkwQKGp+P1+o51IeQEqbj2lUQMR9cRN483DKrbA46DTt0liwo
zydRLvYapKkO17mgmE0Lt3U/m0d5HA/FteG2ulcAKhD+spebpKfZqFxqWbhyu4OumQLyH3hd3FSt
LNoRbYfEbCLwDbfeqAGjvnX1wKp36L/D1WdaDaT6NGcy8p4kQ3wXGYY+vSiEZ3wBuBx/65sv9LDL
BuOzs5r0AEa+3VecXl66N/e8uDzMC3GRyic0y4Wsz5r00uU7jCxWKN1FNZD0skRwlWzoIj20V0bu
Zggdt1avZXf1CKTfHReuK/v/nuZBJ8/mmPVvC4DW+1Ms8/sWfjz9rZ6on5RdBhifsBWNXiJtCLsz
y4S8ThcjdPGpBWDKS29pP+lGhLrp0zdgrdD0bAK52oZq7Uh2y3EljjLA9THD8BbmfR4YCL8R6gIY
P89PYZjeGIDwKBh/B5aztRt5STL4EA0ZYU3GoVcisbVoIzzl+XDReEMXzv0gGv4OFVf59XwngyTv
CGhb6YVShGFx1b66tQilhPS9dL4Xyau2SRm5fqT71TUngINdxisdLncg0iM7aO4qrbcCxrpt71ud
OsNl6WS69hKA/3WFp5k4ZjVHYnQ0LzLpm2/LwBvzNcluwKClVq1QdCtgG07XZEUwBgn+z786bk3c
DkYnUghEUjULLhZw8YQ1BPVJ3W+/76TedHTATQJSdoA6bcfZ9B5ReWya7Nuz78kr52LC/P1dKjM+
x8zt0uFAjhTJUbH48SpSZ4UmnLe21LeePH+62vqbYtN+dwWqMger+O/Ko63B72IRMAQjDggzqyJG
DELbFer9OzTgnMYalnaN7SPDSzOQ1wrNGF0wqmxvRvybwmyz6wNotsT9pVf5ku1ZDGt65XQrHMH2
W1KIMvrdMRkW7dSN/6rIeVXXb0ptmEHdd40drLNNVmsTzdUuB0v0jVlLMMRHkttVzVXCDNd20ngO
RyuAj+OufccuLlN3SrVkBuRw0njb9sTwXjHtqro++16RnRwz+Y08kx923yZPTCIkjJ9J83inwoAb
Dz8zLg/igjOYQrs8otL0h7o+QeRax+ylcju2mM9M9PLEhyvKRFBgHdU8OVLrpXdUqcP307G6B4Fh
nbghlwtuf/pE2+zNU826fONolxBVNmeMQJ+Yopo87o4ogYXle0gxMBQh6QADyqtbt9/Luq8JbHnj
y9NxX/+EcNvuiGjebIo9gSHOgpFY/pxgNglzdKZ3NgE+cYA+6ev1mt87LhK8P+mLR4J+CNjKX5m7
XuV10STpyMoZBPxzUbQe2bS+EtmmcrjXEc8DLRUqLPrrwHpvcAZ1liB3uypcvtZRVoa8gZEIgWMz
Bh2RwNFU1Z8q2I7VhR0T7kQqdxEWlX8rTMkBmOwugN2MUXNAg+p5swGKjK+uTtotGdi+meQSrdpS
yADaGDbhOtboEd2BmiWVVEitXRO+HWJ9xdTU2/xJ3xPm8wC90EAAqFgkESrhdoU6C45E0Jr9N4j4
SsNPvrSZVm1uVVtIRS19AdZUy4kFjeoBXNS3W/4DjWsSaJIsHBSpKhLGl8pyxko1k5GOM/TSOzEI
G5Eg0e05Z+IR37vG+ST7+ftIHjbxPXIvygzMp0HRjtDbjjK8QkY2cyY3kjv8A259GEABVBEjp3Qx
RV9PwMvbomZMPsif3Ne2rdMcuYFFJlD0N/zznoIxCmLvKxI7UehYegcQNnl0IW0iEE6Zo35GXXRI
QVFRWfGgZhO+VdJ+xs5o3PWkF4QfKu+cnG9uMWVLAq2hMxGQC3Fk9XQej1AzM7JeGpOA+/Hi/104
Wq7sXscQ0SglIcmwSLanS+tcovxNaL9uizhbz0W8IuRspxiY9cH/WTM0BpcV/6ZqzaB9Fx0oTJtp
zQZfINBoDnPF7IbwzuYttonRx6kyyo421wpMU/l96fK4rjM3U9G9CGJdbgotP39hNjHLVLSL90ZA
lbAl3Xa4jnErQwNhulbWDsdbKwE2SOtbkDIXXLBk+ttMfAnmKjqjWO+Brm+4IPU77zDQnqidIu+8
Ao17GM4nG869U1ohZVjzOqmPvcsoh4PekoYcEfKaLLbPuVfD+TrEy55tnY+Buu7n/Ba9lVwI7igA
XrztFKsH53pzxD46WMzCU69ykzUi73KH54aPYNUmAF/MnyOAXaW05CWquSNCHbvyWMYYa8LCOgLx
wRXOgMN1CtEalNVyI7MeoP5sADGRKBKBZdV5CDLUtvYi9RQbf411hgw8wQJI10g85F23gjS6Ehlj
S1sA0AIZ4W41vHhsstueb9w+wYiyfHn39RBNvAxjxifldr0SSR5CsKtfygyXUuGsmFA5lsnsEa49
+SC7ulrZfca8+7bNhXT1wvFO06h2osrMk/C/IY/TXXXUwmyysgVFEOk2WbdGXnu13YWJlJgzukq7
GtDE3xvRSTv2UVDwzWSDnaREk8HZeiXTBT6iiZOBctam1kII0EiJt3sYUdRQnFtaqCHZbGWirA+O
obvUEu0dE/xwmVF6jR1nBukBouFbc4BsqA8MEALShTZx/ollPIwZckMP3u4NYuvJMXbTAdaDcre0
2h0KZ9nhn4UCVPTQANPRCjOTR5v8t6GTP2DcXundzsJ6lzu8bcHWYDZpZ9ymW9YldemqLfNLGatr
2ePafOrXqCJgCWE0P+mbkoyTnw4wsz/gZIq65MzaTLHsN6tqGM5d7hnfbMLMsRyEwqKA5N0bvQzs
1OdOaxCY9ZkYiQSSOzXrTBegQILpJO7nJfKhS0LEBvJKi6xgcCQKX8+SNRn76v9mQoTkQo7pYOEr
gmvBcQjDc3yd7Fm6D5OpEng7ZK4nMG1WJCrSvUCz1ekrR593tvv+VmSBmH2BKCuylGV6BQw/mpP1
sXVtHv/H16QxgrqXkHltKOtaAHm4+I4HbtvSgWyjLtLsI8IBK3p9ytthCgCWvtErFKSLdWov/Fu3
gfn4aOZReSQpOgzcpNiy5e3QFISzYrlVkxVD9Vs6MJzxuKGzpEeB34Ulf9wfwPy1d36RUHiEA9ig
FYFXX3qW3MwVnlXHonIl4kD4n9jsyXq4Rd2cZPQtz1vGZ2gMKHmKKymvKMGlr3lz8EQBXQI5nOEk
R3OctgMxsj8iOMqc8grPNzkystQ+2aD5RW5jU31Qj4Buk71jyvHInHCz6Ljr1DQnVwx5jwA1u5IJ
LfnpoUl/eUyx08y5hhS/fe2UCGSQbWQKUZJqIFuFXDz4CugzpXUnolWK4NBRHJFNiJNsVpGPhzK/
Pu7HrVYqjGaaXsFx5+Jo7PFJMLfuMoNRW604uSz66AMpiKKVtG1IXbmvoPSvvlvZ440DCo8RZAJA
0GytF0DUzgBLGSJvsIGbaY5EPNs+8j7XndIXJjTOtiFjRkTiF4DoVpbwdd9ZJWWQhzxu1khxhQAI
bLUl02ImqKVflt6ca5Lkso2+bYFTF4fiBEDSaW3u6S+B9NJF+oXfeFN6ugQ/kw0DkR13CII5nf6x
r6NJt8NEMXnSUG1dH0my/cZi4PpovNhJLA8PQBeinREPVhrkBBvka/3qukc+a9DuJSd/dw+65XBb
09wEbj/6L6+uaSvM92ZVC7iUPAYy2n2XnHI1rOMj7SjOZIRlYTPM+zl7F2qb+DR55m5l3kUquu8e
OT94IoQ4D8rlLqTNXzvZLwiKJsHLcdrV/yyLvSJzvlC6aFQVZrhjMQ4NLCa15ZQ23WANSS7lnkC9
mKsFH8mAcF8mwih9eKxsV37OHexr87h6mpL7Pd3iMG/P2izgQqH/9zm/O58UkrzQVs0+mkXSl1mL
ZVpnN6WP1PLu7f406oKVoo+sBTImLGY31GZqKWbg4Q1+rbqcm02+OrlHqN+gDDU0DuGjCrxoECW6
zmx1NjOu7ueJWmK+h3988tySkRHTOrsKfCMD3ZRu5tIKXEe5JKUNwiDa7JKPBm2J29YHJY1spf9M
J0cPdJ9X8E4Rdd+lz/PMFQdTDlxm7tgCz7RYa95H9w/qE0zH0y9JCGbPklpTxIALcGju3thAfCu6
1TCGns5WZ/MfifDKHc44jmd/j9vDwBxHsoBmhaq1FgWe+1LUbL9AJNt/N1I5QexZ2LiPZNQuQ9Jr
SAyFWB31n42rKcBy00djIIdCQxaMspEepIExsKn71jjzrzmCEVZfKkGLp1NgZXhhCTYKMvoSP9/Q
Y/MOc2zpMkUwMJO1YRfvpSfWKtp+klf3uhUhcWQFAg2LE2nfOT2XCfshfWvGtbSbbQ87n1+DcFDf
brTqVgbD3kOcaDiWnQMEhOmfFjT+63PKQhYNnhG8bF9G6HgTaqCLvI0JgM7X+KJ59tUWPuv7JdQF
gmR1QDxbEhknPYKaaCT1oGYxhtoH8nqipnoITHf+QGBZXrc2TUlpC2ofYk0samn62YLQVen91k32
hdySWhxvmTcyfDdN65oGkRVYSgoQPYUpnsLmYijb7tMI2VAsvRwtw3xIJNjNU6r0wBPyDZq/vfOW
HodKrD43QE+LiK2LvqCXqiDhpiplLa1TI6AGlZGvE+a3i5m+XGhp40vGgo3UQVdgIE3ab16fQ8mj
KN01qOPyWwZ1xnZS5xt6bidLBr++eHqygJpVgKO2rf+d6841ti1ZyLLPy4DcSvLBu4aKHfF26Ywq
caLfI5/ORIakP7W4c+Ip1CnPN0wNQrCFTDtALlQUZbW/cISopDvSbB5fd2NGCOMLeLElzDEmwYHS
Iqg2mUtMOl60OdE2ZGYtKWMYGCYEo/pvjEsD+lAyTHKNef3u1ioeI96EAULJ5xEPxtVt1a+VbX/O
r9YK/QiWan9vn64w5Sn3tEuG9Psy/cgnoICJUDYfW6qe3x5s4g0a01ouZPGKokgxPzBh/A/Rfx5G
iacrotYV9ovaF5bybUCu5hzL64HxW7QxTmT1ul15PdWzkmwxJqTE33q0qn+iyRJfGJ3yDCalXdV8
ki1R6UeTSqxenFZD33/pULm9otdg7L4+O6Fe3pLBkyojV2Prrb2ZCW0KABk+B+MQFdiIZG8R9b99
au33zGClgJeYGaT9sg+Mjf/MkuryWuhpaZJxW9dU7TUkpS6UfFdSq7XPyDoCZ4yO5SZysJF3klTC
z5T0nyKVzjfcLE/1Zsrsr0uci0bvOQlgMPZ/I8lU2QZ6DeSMxafbyEKvuJSEf1lDYwko8tJZjdas
jLHP4F4MWXfLbfjC3x8+hux1i+UNCNV2UAIv5YGz6kDHme/EdnWECqjc2N/kl662o6OWrQA0fvzn
RFAgf5i57K2bvROM/uOL6Up9hstXUQrbEEXgGeUk7jZQKBVIpX6bhQKZXBG3w2b//8H0aIqHc3i8
HDiXZKy6Lv1TNJVg9CXArOUttckYMkpp/7H2S0o1odjNN4ebtu5scVoJcrr+Mgapj7j2Sa9n9TGx
p3f5ht6YXF+bJnJd/BYrefxBujfIP70RMSPDBAPj1X+9awsz9PivpiQbzejTlr6z42SOcKp8KkBf
sLm7Kripci3KE8LQnpVmA9JfKF1NTc/1mQAT03L3C4NQUtx8ih7EJiJeHHpj9FN6Nvh3mT/k8tuD
+gm14IvBcecECcniXOqJyFB/RCHn4IWWNygABzf7yiOo2uEl6u8NKeSBzCQ6SfSvv1s+LWM5MJSn
Iqvv8HssaFNGVE/o485Vfrb1bdgV+nik3KAIu1vrAerWX9tn49UtLfTtr9Ib4YKXu2dIRfwKLz15
z0qC44gvTBkOcUe7IC5g20vbQSE9gj4a8J0EAEn7aXPlt0Ep1awwACKH0nl9gHoBpJ/Gc9sZWzO2
Yh3ydmi6qfezn5XgrfSy7X96qxKbIWYNIVOmJmUpknFhmMJyQOOyjGIlBd9cXr1+ZwHQPC531Wt4
4sV9UllRU0PYO2Fi2jXkZZv2r1I2IQqmr0FuMKR/9SfarRtivsK1AqHH1UTJJxlkTVcNo1Y3Bao0
NI/JelExyMD7LRZl41I8+LokQMyIv3saS7XyE9zvHq/DtI2w0EeGByGTcFqNmR1ozBwZvcCl9po1
8hZqSjCfD2983zDBDrMljUJDkOg+DN+uvoRbYlamhS+EE3Bg38oqvwxWr23+YU6zxXoCrfz/Iy2V
kuCv/SHJ3mOq2qN4aEuCgilEK0e6MxJpmiNejQ9RlxOMl7stUZl5OrRmo53pijy88sDV615g9Jev
dPXHmy7mueXG9HbtqOoSpiR69La180aKXGI3iIdgLIb80l7LYZ9NDvrZDW0s92ywo1cpMy4qavRB
l2RoEBHRgWVuDJ08Wp4iB8+lIXJWYv063yAwZ51V8mFmu0WYvbq+tH9xaB9Wx1fq4VmWmvtYF70B
MsEvTZmupTNHkfQMANnreOjqARBYPa/HB1bKolUjTG7puPPqsOq1Bg5JaQvizFAbn5B7mP8vys7O
xfoAaMFWsee/pOOjlPhMNXerf6WlujA2Z0gq1bTn3CUTNNTaZtkqu4sbfuD0fw7GZCoXGswUv5Bd
Z6kkuiW4UeaM+Vkvk9pLNpCja4CjLDNWVkWKF/aLrw5/Heb9SPQ/dQ9MeEQS4HF4mOrGlfL8kAB9
vyCSzBODjR0tpOIW8OcU8zJQRN1ISUONZPhgZnfGKyJKyrbKKx5LCvoqJ5SVd/UWSNpTfJUIENid
otUJfiF468nOaWGxfjJWW1W4GRDwhc60GU9oiG5cX6CWepMvsPGDE8eD3w/3FxZxortasOdgf8lB
469FneFxP1wqhEwhZRXZMBCWg1WNQV9FJxIPvK7CbQrfv3LCchLIRwjlkvB/FBrONlDVqXSSvhpB
K1lc+XvbR5F3s8GPupQ+J/kqpfC4/ib3XcrYNZeexcI+1TtCRpX2di6Cv+8SNLukTyMNzpOt3MFs
PSsyB7ePIBHhmXbZ+vEYZTYUiE2bgmJyowe0dMGEu674rG+MMkd5vppon77s0KR+P7f9E2GUT559
nLb4mK2PH7VnN0gZ66RnSlIDVVGoy1WTX8cL9sFSJILrtBmzC/wirE+Q0RzbDNtlxxEAApHwld93
6uigJ9ju0armr21djzLWiJaz6jb3Cb1vc+Aq0OBinsz3a8g8y6rD0Cudy8j9uf6j89xrNXrvop6K
rXohxs3aZ9LBQ2ejxvZnSeaRpwui1fuk02JJoFXhmDlafhiOdoEgO3+S/LOJPqIVPghAzc4p5fnN
nly8q1X8SgW5OlYmOGiT6e/EjQCvcD/q5B4oPfwHHLmdqVShJAh3AXm6kA/mC4hrU4fv0Sz9iEAU
db0Evfc4yAaEYsXpOQBS6Pebx6J1TISGa9PJhkmc0sDxlbQY9C0tqHElrJocRAfwYDSo8bs/pHBR
YO3FBMKyPONInamJEMGoGQubUy4Lx3Vk35CK7BfcsFafTLBqQ4P2kFBU3xu/F72nR0z89aAeCfG0
ziKvb0B7A9JOdtzMQ46ftjluSnUDwZHdTUAMGzasWPtulcKFzyJHYzl3F+tD4h5pNXj7wZ5xHWsA
ER0PrG3vXAmYcPdl6GfejN6Ip90em3yahUq6o3hxitMBZnK0j1IIRNrzwzBIxJoHd3//9otv+wzW
f9kIUwLrCupnQRJs+jt/OsdGStneQZT1dD72Y5EYjPMtyRjUOSnHi1jn98qJjPik1N77btQGxXGn
+HTq2fDwlE9vmRv+xuVobX/gz2SwY618txbzjvC+c33DnebgwdKx7SHh+xfAGf0IM1XMeABdRXh0
JEnCkk1hGdf2kbhjEkj2FB2pBP9WEQPr6SjR+7/iXWMoFP09X5Mbx4C24bIICBoPHb3oKkzu1q9s
bzvBdBANEwS9Tc+w+Na7/IY+liY3IxIryBetCbMHMqN1EEqGLrPfg85AYasX8nogXAjMY+uwp0W3
KBAq/eO9TVC6Fr/1nnBzZSqRwfCtC6om2qypEFCNtK+XOTSChLhCIPMzB6ttN2dLmY6U71TXKjMD
si2zxt03BsNopb9s1V/91R4NVxpMNT7LBU6u7qwVefcff652ICKwi5bMetGTLrOokmFIJvKPErmH
r424kAsJLBgRM13fPgzEwf0T2rSZoYYPHytmT9PgmOmFiQj68MXQ9xI7ry8dayOfjqcl74sQelAX
tQgu9hjzZViAGskVDcBNzbIx2OCGNFBJOzxjrXmGZz48d2DzndSfNmcAygUQGIZmX7jvb4E11UFA
BK0gXBgG0l4tLbRAPMDWS7CHylUNJE6eS6AvwgZWGzZKHd4DZS0A1ODzHy02eEHoFsGvZgay34nR
EJpFNMYmhu+AisV1vKauaGEqS0Mcyo8auQxdzdkb12lpXqcrR5aRJSBpV97xMLqN9N4CxjrgkWp8
KwvD+ZKcQmO7EzxDSPKF9sZPdAi1gTqEzT/ExLnDU+Vv2w/r5xWQdOJ/qbPl5KdaWXwwpoMxnRy7
ATgVF5IxyY1b0MIoZhSHA9Sw5tnijwiiFcdhn06W2XGPwsmskIp4XsBKwp3oWiZcXaENjXiPgNEX
Meqp2/k9lSUh99omYICPU9D370MFVSbQfSKLYfM0PNEJXrxggJPTmx1M1Ge+UHzfGhCkorSUWcUh
mpE8Ser0nPhRGToNPIZ4N6Pskkw7JgchivKPQNxS0OgtyMZrBDn6fgnujX0vRTk25Jq6CIJGyhXt
36BGiwETeUeQwfNxgsBQ91uTDG5aGkf9H4wE2iF81pXHg2KPsdaamuDH3rv+Sx3QZuQ64olCOhBn
gXZvcMDozf2vLhJRAELPMuJVpu8nNFWI6HKsfdSwl8zsdZ6WXkKTR/c/IHLXmMzntZ0RH1yqiqxP
pMMkUsoFZplh6oQHhmmfxG47WkgZupqXbNbcnOgfbq05bRUJf+In5yOn4tSFNU9+dVuUOyeRsy0u
hQxjtpcXZFsWg43TNGUUc1YZgyNf2TLdKoV1pS8++gU+zWsNHSyVmdNSp6oU+Bylm0N8S4dOX+wy
Bf28W33CxbHvcxxJDFZ/kq6oAl79BmXsLkRT+SMYKwVOEkyUVZETW3XuOscBPIvpaBhw3ff2ukHr
8TJnnKE5IkXCaYZYpIGZ7j3qIsDPZenxdoC19ZRyVxjMVzbWe14hCIAYAUKmRmg4KiFXenf4JWrd
pHCTHYBgCPpUG42eaa/Yet3yKzlInLHJaYnKZq0BMapANQoKzzdrLQwFXPSFEt7crLQlBBs5ERgj
Pg0GWQ4/ymAWWMjJV9DHUMJxWC0pbf7bhriNsW4PhjtBpGEmw8BpRflIVx0rDFxmzJwM/87XaaSL
yoyNZyvo4oSFIHXrY6rzxj9IbodIibX26h6yoat0jahF91fd9IGbniDXza2L6mzcwQh3R0Luyjp1
n8WR2uyVD1TeCAAid2Wfrcofrz5rKZKz53rTsjsgOnIpcpnCnK3MzEo0I/sna7w01r2+yFaLjhol
dpj4X4HR0GROPoPR/6l+u00GrpDSSk/jWqRHUX4pOz6XLeuO1WbDnV0F3Pi3J3WbkahSiz99ylYX
fwtIAaGNrSOBDF7yg0jkGWGmqNs+4lD9IdzkQc6zbnJY7/07wXSGh1pzqckeq76qhOnfrtef93vW
ggdMP0x7nlIpNZh0Zs7PFzdy4k/m76DJkSHkjlGHdaFwrfTUnr2wGRM2xCxQB2aWiMUCSN425Dde
75jUwtyXPoUg12D00K85fiJ18nuyrGIZo94CmZ442npDXxn+iPd9BYT39r42Id0+R5gkyVQvgTPe
AYeZRfRht7E+ci6JE9Pj9IMaNjQO11fHparelrVto4sbbMA4jrx7132LLrH+GTBEtvmwJE2osOUG
BBu6clv+Yc2hW/RBUFQbbwvjLv57JjdYm7c9lUqiXu3ARwCuELjVX1Cm+CbSoKn5h55snJBHeiUo
UbXV2drgP71MSjY/phJbbLJDdtUCtlcwE/ZO1UYR4SG4GkxtTG5y4ot4AmKU0RanFpsYpDTh19+K
pczpeT09iDOzM0gUGumrH1hBho3s8rZ0ZYHzVpqbbktgJa/v9kUDbp13Xh384O0UY6PKj8YEuP+G
y3W4N9pFX2QHnerfWOVd4fHpLNC89c0EtV23sfPVucS9Sx1WUyzJS6vRx7C0mxKtjbllgTi29Jpm
LuPERlR5cRcfo5AnlSDV0WgMcm42F3FgRofCc5BeBVFKDeB9GTqF2tOVuVgy1pa0Y9JfzRRQsAkT
jIaN6Ap2aoPr7zmlhUBheEC3Wxt/9q6Wady4kpM9K0g5vn/fxnsLiBdWB7AzWJ9HJUnKmtfekN/u
nAQKM2XlgygcUKk9WPwrcpVb2ernWnvmVauWXO5jVpG8mNTtLhXxGN0T/1ByHKj7S6/DV0xQ68xW
9/WKRCqRepgEbInfKAYizd9nE2Ioqy0oE6uOQqui+Hbub8rPysXtA2+2Ps8QiNZryEa2GJWvJS+U
un+Qn/kDW0Acn+waTnJjB5j4nsyxPTdO7y9oT9LtewxpXAUkXKWocMNuquoQUWXxOnn0XcLGbP0k
/MtU0Oufm89gqYOVXH5fu2eAM17TvrSnqQ+KuONulDruZQr4XY3i60Gu9OUCsd5FnFWf3TzFfL0w
B5HqtfFm5wJ7SmqTgjDEqXrXJReh2xSDF45otQgtJcXhLkjXRg7WoDal/uCBC0ztnoGMugzvJ3kG
ViZcrFaU2LuDxsAoSpU6Up3g0vBIcB/3mbnLn80SQocwzE3jOybcq1iL3iYU3JXnR7HbXeowmCEY
ITnxf9PMJkKOT64YYsaeZWFlQEExSbrjds1ce/qg/lw0OQjkQ9+qVCHjaSLvrUvsesqaV2cz1++I
8RokDWb78rjXm6fJxlGY0HwSf/bqJPonYp2SehrgwjAkNJwp6Fr06WCVo43jX5eNVslD3RTwEy7i
S/2YK0XikT601enQCeGAh4IXV8iQALOlZslm7rG8w6x9nzpPShBoVcNCcPQqr09w465eKCvoaecn
ZA6PVKAhvq8W3KK2DwKs/1Ca4ypwopbP3i7fB2UbOyFH9UOs/v+xNOdgpgty6ZwRCnnlb0hHbYO/
8Q7qH3RNK767xjoCmPtS7+44Kh4Uy7JsB7Ty42kEGMYJ3p3q0MT9/UCk/SJ2sjprY+BHP+tZYN8L
bYxbU057t4z2moF2d2s716H7CBTZMjutHftKxgVq7Y1QPG3ArIIMWeaR3Z/se6Chl1G0bw11/1uB
QCgsm5Lu5XV6Fa5cn8FhvraW5a4MEBqwiRQ8LJDoboMwTDfprYiw6ns2/6QIuz4eIzhDiFDjW/Zp
IbsJq2i/dznJvMpeNYnZncUeXkwpqzQlnh9FLoJUCj9SmzaEIvJ628pCmHyc6napTE7Efakg/z+x
S+nikdujr7u0lHVv6XcTSpB7/99EmlfA3NY/2CBLO6X4iFzx2HZ14nXU9TOWnV0oZiJWDuAjq8Ch
/2h07iYoorTF8AX2VmS+tBVkqLnVbmejQUTrw5P1Ujmx+JEFbQO88QlCNSy9awvfCOPMw+1LSWMG
uG/QUEkTNjQJaacYGywudscytSOitY/r5b9JcR+JgGNcNKqiDkyTnZfE5G2FRzkpPKSyR/jFAZvI
HP7Mz/ylRH8PGQGEghJ+Lhtv5goAA1bTRd1Ymj+vfT1sVXKUXO1inKhGbxMJkezBq+TyIad6oCss
81ARML+y6EWC3X+jAs/IlKFRoe9VNpS5AtAYsCx/ImA92v23v5Ycqi4LQIGv/rQoqX6OVfmCLQ6N
hZ5sNBGQkxMHnnfmnHX3jzJcMnx4iip9WFu2vPY0PrCvb3cTuZ582BT3n5Xc4qyZ6SGBRShXp6H1
JJogPtvkK4Nj8JcJEr3LYk7AhQsyGv6T66W8yW7Y+1Gkb21ZF83gVYiiKOblKpzVByxkFon6ivSC
cxaHPvpgC5cy0IDKPW8dQ/H44XHN2md3KHnNuUuHLJ7X66Za4MOMTeaiIMHpY9PPLVLjhN1jwweT
k4xxVdum7z6LynZnbPjBC8lP4mf247izpQYjWaNU6mbdREELO4XRGIPDrOLSaSN9VEanvUJSHsQU
63fb33Bzv6BIrK2xFd4DopZdcqY/hl1abcZSksMntM14PnA9D/x3YQ5Yl0CD5gcr2IbjVvx1GTle
w4XFZ1y18ZCg8ksq1l4i6FuKVZ2cygWsofZcH24P8sndOgc/GoJ7Dz1oVOfUmFrniu8U480T2SAw
TvdOjHajgdCTUEvVq9qy+bAMvLmhv+5ChO8Hk41dE9aUZN7KRdwscsST2OGWDuy97hGJ45ISNlT2
A+gz+//wqQ3AjDAhBxICOYk4yGt2xSj1RicsvgiMkG8o/b62t5rKcdDGjXvwfxraHLt4kk52pape
huZ8ydCWJD6yCSMa0W9iP3XtZCuKbK7Zpnf809Fw8rwO9xOyaVq+oOQvQhm+X/E3qs1LMtVmr5+P
tDJ3FiK6TTqQd9q38ncvPDi1TV7v3bBP2g9kWnWFHOUrV+BQHOgXP7upwrcVSHlrDkI/lRur/tIk
2THKxhJT40KophSXfpE3tbI3S+nOZAE1NEhSWS70XKfTbv2sj5OgOOk7s+tAU9XfnqylwE14xnRs
yXvwj/Bnbe94UkWVIOooLOvUOLvYOzNkMSNkIpjm5CYohfIM3qKq+f5Lp0BBeWMvPBvBjaX5B/Ka
nfGIT8tsOQbaSdJyweku09QbOtTISr1mIessG8GXMKywVthXq2uofkCCJShhPmL1xhGM/VhnHFdK
+WqaefaW/ymvN8fc6S1f3HFpGhPASRTxQ5o9DwReyADr2u17AXqMejrPn5ZWSa/UK+wL5w16F3LJ
wevxi7J66YNagcHQe98pqvR20+7UB6V+HdoQ/0W4ZFix9cfqOlwWvx80410/36YlZ92hBnnqMk1e
i7avvPtYQSOZgZsaSPYeppLKBzHMH4+pYihvX3LA9C3vcyFye60ozQkk6Bts0REmTtr6u12Fqrma
lCEzbFY5ZoGeEF/7v0xLEif/HdOAr2CkneaVATdZe+m0yG5oBOuMb1GWdmszXJYbhV01WljJjWkO
6CQS0cd87WC0nxQFXZd0IgHOLsml7NZxSKDm0nvQIgf4rT6H8kkM6TO6qs/uC8AvtpqUacV5XzYw
LdCILzFiR6Tx7T9+XVtbgVsJJz1eUmpoTYL9wGufVtP7cCE4iVr3VYEkV6kTubvWbUwPSzsrFM5m
Bw0SlN2taES39UbROuYdO/TkRXi7u1hVN5JkFMRcaO7A3m10iabmJlf3SCr//dMi7aLYaEdGaFBP
bZRqHeagdpMbgzrd7k5c/WEOudfpJFus8aOyDChqRXe2TOlKbYS1xBWDox5aZk1DPL5AQ51gsbFP
Z/oL+jOoQecxovT4EhsmuG4zCfyPOuZ+bChvzqBWoX7VSurrTjq2B0KdWifQBbG4823p5FW57jZP
SlfCkdrZVZ+RuZ1VLFHkKsmBPo/NoCAEXzjYkvu5+GIOnzhaxXBpUObNA+ksNohK8e1l2HcQotLt
SpKHAvGBNhOhDFed0d9xbBZS/2aga2aaN6TjcgjjCXBRhscLDD5OJuzyU1ms168o1oFyNVBI2BrC
TgGdZE2R2w05SoVPc+TsYjuqIMlaXO+drYSgmlEsByHJ7516NuQTgmRrtwQFK5xh9eAD7RXK3m5H
r9Yjf2cJeIsR9bWF34bd8BZEb5/apOAvRT8GCd4kB5+GMkeDP4OimRpwje4tANDLTaiLWkFy4k3+
A3iOrkh3GFvVtgrTDmzZY0tOzQTBZt5iRJCDAym3ZNyKTsRjcXuEFNmc/4emFX8kniA9oh/kZpWJ
apbob82FoiJb8TVVfuNhKjISytBYydimnrNP0r6niyukaK120uFK0jHF1mvTVzbYP5KrjsxQKl3C
WnoTOvrrA0klyhrZFyNaPc9xhN9gjxvqzqVn00Hh/+6bKcj0tGjXVi2qZmyOM1PQQIu0CWA4jQw2
qWCDHYhNS4Rj3caCNeyIvcWgmNqDMGoPxw2SzklJccwTL78nLw0UgdPDwVtAYxbwZbLJDU8Y6kcQ
WCsXir87hAw+zgZMGA6uifxtPwa542WNtQ/kXLHjOVgPWOb4dnG6NHfivyy3fG2JmzYFJaDvLtAD
Ig/xap3Pryg5/LGswwRHNbTUAkeNSbrP7dbYezlH+HdJun/bF3k1q07nhv+hPQc2qxw4xjckEGPE
cGhciyNX5xP+oXalqaL0rEAqN0AGXpAgtCRWl8F5bPFQao3WG3jYoJ+zXIFe16WAwDOY9Pgx9GzE
LnMvS5cuytjBCqLTragnJFF8+W/PeE+Eb74KV1Q9BDlVDjFZWqHyRvcaYvlA5Kezp1R4ytRLzsW4
geePx4cygn6B3UfE3bgl4c0alodFncjWljMauvfSWi6e604vh0a6M0rIDqeKQrMqAW8h2JUIWuSg
G66q/wAqGsV3spQszXRbbbfVslzU+YEr8vP+1jajmQZ5iFb45htiPoFbxVehhQVpl338sBUbq2Y8
JrX80S5RZaAH6/NoVoKUzDCHDznr2kCw/iVfZcfmVFLwjQvQEpBHU/lkPMsSiRhrENuJ2AFRu94/
zIPcieGjEAeF9cc+LE8SCjoZ7PlIkKdZ4frBtmdCV5AmhXxvK9plQMDQXGuBzhnZpYs4C2qzJ4G9
0cSLNYh8sw3eGtZMgNcuIxv/PZDuHgb6nJjgeJQXP59NqZCu80EA9ZKVqQNVI5RkCxe8O5zcy3/J
6Pq3g2CQ7LrwytDffbcrMt8NPQcAc03UTs8FITLq/ypvFWu+PlSGRIbuWu/WaX8SPmXggiAmX/V8
IRSHslzInvcL1xdc7T9CmFtwyK/WwGsqatFNtlGDP4N3+o6KF6G/6spgZlyUnQd5L5vkG+T94zqq
VSHsGqND7HEHBTACn/Wq79JoDMExovXIOhdNuJYbeyhBCITD/m3kFe4g1IP4UUib1B/KUKx+uPqi
JZuCQ4y6IlTFX1ZZNKqXriU7uvX8ZoVXXJHmwQ30g26O3LcRk3Dn0BIeL2F4cjzxmnZGSDHIWH/S
suKZCWW/ueWuk+sBvaXxcCNuGMNyOHRDWJjlazYeFsqDIwVEQcQjhl2XCuP0DB7JsrudSIYiFwGp
dGQmfkY6JHwmdVrqhiC+TiGRTcjUcW41C+jmHr7KOWi4Sd0eFcvYmvaKrqpNjnP3f1wcieFB5Et1
bgXz7xRz/BY4N0hHd4ES2wle5LSC4TBmOhUGkkvX4m1f2EFPtdA0GTa2EVyyFvAcTYROnVRlyAVI
2U9xOPUvyrICYJpQ5/e82OizgQG79/8gy/HqKez09z6sXbEN7t45dcDnNi7maFFtEEqaDHCi3MnN
HdHSbRDKzvd8QpYrmd5/iY0j98QN2skHdiGeT9GeJHd+JEv8GVXoStzoIXSmYRsfimhi6wHFPasB
TttqOWos+VKqrYr377F1ZE6jgfsaA37YZpdHwdEkdtDESqhBKbRaLPQf4vAabUNSQMzwhOnCEche
yyR9l+Bg5BJgT/jItaO+xF7zQOAZiK29wq7lMlX3j1iWnc1fu33pIs//giB3mpsjxmzk2pETUjot
8BCwzLAIDylicTnsakAf6wQjau0N39DePsNjhKTWUN9eE3WurcC2y8jSuYxBXmj68eLjpBaC1axi
XgIMaJLZNDFTgR483pcEWTuHfexrQE0CzBAoEYxqoVCxOgtPZ6TCa25ycC02U0Pf2qkgAEOKXqFt
qrpjYr19rpSbLUvR7VakfOVcENz3EQyEzU1DuHKkoYkR0291i8lFVoio7VQ27kV9KE6WfKbPahsS
bCIDqCvEaNZSF1Bw3wTZnXrMEc1OD5pjR2Ir/XD6hZDjFAgq8NGo/KGhIh+GGIG15Ky5dmsxpvlI
NwTmJsWKklJzaroDgJSyuzqOMQVUHk2w8C9+UMOlWCy5GhfZRB6dUelX0dK53UM1dLdW8+QkFV5c
kYseaDaTTsVg0rlFBh2YObq6Wf1tjwwpCgsHdWIsBSZGfgptScMeQDwVoG0j2xN7scbQ4wPXFCdO
VBfjxYtv8b3bK//IU76Jkeo3JqRRxra2T9HrHq3nMN7CL8EWXJET8MtwV4DRw5ZHUbBWS0S2tdTL
YxxFr/WYqhLa2jTjm4XLihy6mqFtPYiCAiBoE4v54jtmB6Ea8Ub/c617bmlTNKc8ZIYYp6W0gDGi
3V6VZp2sCfI0GgmI1xzCqBBJRXcZxDcM0SjOhJ0hgBaPe9N3gRyAvDbZnDWGHFFIk+Z1wMql3PVI
BmgNnLzR64bjpE7A4mQOyjbPvLH7wi/kpCnMKOPHa+KSEm5+4DrAuIJFqwbx4VFRzEvL/mmys0dF
BNMG+T/AUlToSuv0Aar6hBgJrpY6RqVZ1o0M1M0TARqfhP5BAnZvXp9jn9/wJQE+I8fmAfqpltrb
xDu7cSxNBPLs3yLaAwhoIBzhKO2MK/4+f9nD2L0M7KhK3sX+2/S18UPKPmqoNdKRiO2whPC/R/QL
PCDca7Sak4M73VUWQ29p+E3BVg6GkhFL4/36hO4sUM5U0EqFyhuLLKIhOlk6miROywNzXwQkVBtF
QEaRwuKHrCXUNoVgmg1Z89aiHet25/ZipzHW23dvhheIBxrsl6ySw4hAwSRFc/65X8P1FpuL6gRe
8ujIEWPPA/PbGAjz7uGaSGAwdviFbhzb6gk0upjJNacaEFK+Od7F/BBY4AgjhFwhofoGQduKTVdF
vlPFfKSOJjsvwVVpW8bDhf2kvhxOKGZa9WN96ic6AMgzcLFlr6oB/A1J/BCUFrEqU4HrcCpYZoIS
tP0HYhNF38KlYNmzSEOYATcl8l9L/L4wjsv93x8rpE2mXtTWlKZwqBcWicVScxe4IS4SYDgZ2H8W
0GS/0XsGznryI7SGZioy+zCvO5IQr71OBET3JUwQt8kJ6VPx0CudMkIj2+NyY0JnoZhFskZr4eAU
8RollNzjd/2GfMHW96WvJ5aIRPm1xjy2goIC9iCPfJ4dq59qRZTN+p0mCDmb4DGF8zu09o50BjmO
LIC+b8MiV7rFLN7DABpqP8cWUTM6h/WL20mw9lMgGBu5o0FWOzXIr2Djwvk+1HWDQw3wEC98EG6K
FYlAOhLSb4jRpT4pe8DH3+ox60zEYyoVw52+SSrhRrAbhmH4k1yxZTvwp2DKF7b8MVpuyxl9B1/x
KXI523oinMghjYm1PMxZzLjeUKslVzv8ltKPzeHnO6JzYWVm8l/v4DnR8CzPppLeUGumyQ5D7RxU
Isr4+Bte+K57J5T6CuqxfAJ+Cx4uAj2eWWHZiQTk11U/ohr++2sZ7x3h6Zhl4z4LY0BMAuAPtDhI
mRJKynCYkgqP3G+3t5eqTkVXT9mI7G7KoEWoiQ5UQCOd6rj5lTm+WGwjy2Q7Cct/nw/UoERlvsMM
r4ycOZAe4JcwLFklrNTd/Lx2wEwoXbqBPuN+zaDndBumRONxkyB/wk0K3hREbFhfx8PuorshOeEt
PL3L2hjq8Iml++uucvsvAWdVs6Iet5jHjRqzmi51teuzf1fnEPDgR/61bFB/AJYA8k+dq5FSjcA+
jYersWJnUqXCz0R8QS6UEh6Wr/aYO9TAKSKA2oj9WEdofOw8/KRupthQUjoZ3BN/o+lBx20D3wPl
Jm/vqoVoTfJcNKKbHukHOpQD9oUX6Lj0s8tx7r3xPI4k7CDQamxr8GyVt5ZofzEYm06CDA+etazn
+hAH+vETjiW/4YFmkURoAkCDYny/Ye6gwp3n6aj6Fn4hUKi+HB8AyirmTcLEUbd0ZVqU4NnuQ4Bg
VeX5qcIUMPGJKougfHVmZTYXKM6FyMaZq9o+O0j2URVzgsjpgGP+FqleGYtV2YOD4CFE+vhlEG+b
WrIB/KCztvx1rkLUBNJ8VVzbZHs0qrnjsog8IwNt3FuW3mU7Qd8aguysRFJCOCWQF4EEwDDnEI6A
iTDUFjpECTaOrhUCWWhnndWNsbnDxll1llcRygX0wtM6iMpFCC8ClM9EoyPalmb3+5vxArsCYxYq
mO9Vh/sIFjwhWv6PyR7Uvdgbo2QyRSZDqriYyV8QPyEqsci3+SE0yStfMMSGQylanQREaLIqS1Zz
v4Z3VV4zRSOhY/7rF/nhNQSXLRYTMAXl1N2XeUzUX1Fw0/viyDghGEHUKUe7bRgifPgocTkAvDWW
wqm7YOSKSfRONHyVXIkix90bOqWdkr3RAmjLgs462nLXnRmR+hOLlQnGVTF//J1q/BJNsxb+OHdJ
LFAkoDdOM65tvGHkFme9Iasep8SqCScOC6sCnd2cwfQM+27zG/dK00FPSeNyKWkfQSXO6ymsOyUF
Qm5WeGLqhgyImuLxw7MJRzCb5NOzf8tBr9/kCV3uzZBA1UCRsAUzAwgD0eMVZwcg7nf5oPXvgU5J
CnWsou8X91MtyVvqO/cWNLO61DFPmXbobKSwO4+mpr3GVJ7uz0g3nuxYoRcTBgDvsN65NxmymSeh
w/1lAfg5fimSlGlvcTaL77KqwcfxRdLs4gO4QgNP2hNgiDMOfEGjMGIADy0GCVScqlO32ewpEBfT
JGOMLk3ClN7mTC/WF0puQyPtvYU1FvgrbjQy5RMDEJx9uQEuSCzpq8PyD/j9imhIb+TRgA/+Nd9a
BCb2JzcoY3gZFX/tzCIuXYJlJtfYzDRrlZuiP5MekGUbNK7NTAl2eissKHlwssqJPit66m9z8qrV
6uM3MnD5Q6x0eOrldZCCeTx5BXdhjuYYLaBAKU++TmraeMRQ//iQSZ1PoZ2U84mrPKSASdy/JUz+
Xgt1g2ONrZbFRbfZKo7nFsyvxuezD246LFg+sXzL8kN93aVxw4Tp0d5iu/XdBHSmolLSQ0E+GgDQ
lHDSd0j4nvC6mFd17KdRZh5Pua3L17fqzfvy4yIL8zRncfF4Um4NrRDXs9yTikW/Cvt0Oe4Cck6m
H/OYS6INW6Z9bxYpG0najdQJZs0UVlRsKTTyIZHPKbcaVV/007zvoEnjpBvAHqiPyawomGkk52kk
88Cc+w7rBfjuekDlLm5wVbEzDV4lAm2mJAMLWCyVCBq95VuK45EVBDgYLsbWTWicSetnXqXZKxEN
//G91jlVOGsZ7XH4bABU2S9CiVszyqyy2zlDSQeDah8XGhQfTnJXeR0K9ZdDwoueeZea87HCuhMj
t8Hr0AjERt3c2uAIFqCVZwVGGzbBN8MQxTkIXS9+7HTmmx9Kl+P5xhfgnLEaQoUzRZC365fLBlVN
vqZd8GmYOtt0TcUH2FKy+pZVC7dWfjc6FYcx7FAzFkmuy5Z2LgZGUD6eAjLU1pVTVOD2Lbtwcvh0
IeZSunq0Ep1kfu4rhzkHwY3gy8pIxydSJRM0bERPV0OhIyVKUvRctCMAv1TtcyJCjEt29T9nxUw8
0ixNtS0k2I9uQaKwjcasxIkP+GrwdaLfqgqF74Gn5jVZt/fVa6GVVLpqNC/uCuD+DQL4YXdFb3PU
qiHxaD+Wn8mUr2q7Tde09CUAYopIgBnYfMM4LDgznzZ5h2H2zU7L2iXQjXm1UahUYiFom5vZelRj
f4+l2aOd5AiLQX1e+KDVMd7d63hcUxSsHT47xkDcMGoLqti1ivodNgbmbQwOxV1BdWYaMKEfE3sC
z6yRnf+o+FWlU0XTUX1RzNayUu6z7BMm/aM5loeHJNdBeJCXXmjxmgyUg4+4joqMtHnWJeXcRvF7
AYnI2IJ01xMSGbB0Swz9RbaBAfKFvMZp901cnn6Xzhs6gsUYAVVyTDCHuG0i3f5iY1yLfteZEoUr
aMmDM7h5QeFp20uQqbQlgUm+qLEOt4ed3vEA81OYQ+jrAyA0LUu2a5zvI+bgD6l/z8ncHHYbY/5E
M4E3zdEqBS4fSlS9ZxT3gWrSg/5KOQq8DVa1GdeqgZ/xoUrjdwtUm67i3q3Q/4+bU2sK579MfEmn
aenUQ+g1AH8xVAVuxVtI37W/OHBDPyoWBmXDf+1KEQ2F4/rGJ9gcQUhJ1axJlabir6KW4qDsUTd5
ENyasMUj+ydLuGWwQ0RtVJC/u2YXYzUVqVCS/0TZX229RTz8pe4R9YifRMb0Hx7dsgLbZUVgqwsa
vYDD2lZlv2pKipWtvq6ZZknrvaCLyY0FGs3MO+sK0DKgWCQlg2itmNKLqVLeeoIX5fxp6Od/y1Mf
mFh9nA6Au25Q9Sh2+4lqoxJ9e16VPQ0fRhgrz0FtIr4snJ7XHT2C/nTEL8VVmbBl1xoe9898jHOo
SULvLAx/FEj/ombyyaY2zNek0Q+34MR0gfSQRclLxxi2hrjHJbMFSR+O+wrX3Ey8rF6Klvrk34/7
OTgxhtPfXmtVSGfNJDLo3YsFXBE+lIOAU0eId0A9U4OIEvK8CsdGWLL4z+wQpHotu+lI5t45/YqZ
BMdhsV4Jy5HC9WGq6NyIAfU7aPS8za2FhKIk9s+C9TUnCsM5gjKVjJeU/xEYMlvuCdR75JkBrwAG
KnlYsQkzsDnOdLvvje3YtXOnvT0i1FZy6jJHM0gWzScUEoOASEt3FivIbB9LKuzRbeaRthHKEa23
PlIvN8wl+c28lnURIegd8SRXvRxyhfqBAyRgyu2aWTWAE4thLqq1A6diY60+fdAXr8ogXfynY/ds
woCkzaX+WyOoJo7QeBsHAhDihdfDb9dmV92VVtfAONobkiVMQVUUusQQyysLOwGIFkSRWn5aWCWc
/Ry2h/05Qa4WUD5BEfwuHjtswVq1ZpcyjxIrbrl2rTAHEL5pKKsmyPjfQybFBOF9ZI0JBOX4QJ+v
GPpOhyopd/f7J+8K8oaWLUK39MZiWNQo5/pchwiVFtGSKtLGaR/X02miLQaH/ZF2ngEklgnJ0hzK
a4vtpF/9klIkMuPVozMWUpNhCTAzfDpT5G5amaORsGpWQANeU9dr++ER+L70Or9wXmjQvACxnof2
x8N7ci/5MCruUEJGaOd1K7Ljnv/b3NlJFFACI5bNgN0KcvLH30I0OfbKE2egvTM3ONuBq48IAOJW
YkqjhYG7r8gzJP73PyPE8MD6dzQMsL5v2ANt50etqRAfxdXzPgwJnRdnbMnFQI3S2wc2Dq9Ya8/X
emCVdHWuROr7ngB1aDEcqRUcTuLQUqddb2/UyIoH11+Bs2gUfBoUGFfHyWjgxOOY5Vnhs7dfUO0t
rrLIk4GbAGi1nNraE/cGm6a+7xQ2Wq6H9UydpMmbNMqmtloPoSwmC/WAuRdjvCRYQNS1XYHU5f+K
XMlCyfSBsiTYgTDx1J7rC4Qa/OIdLBL3gex8MAKGbVfoVCYo5DDbRDpqUFpmhtgqUsuhUG1H4eLW
Rj5H0xezj7O+fF6jKQSIt/B10If5CPZ4kYe81GtxwMxUYDfPJ/tbxVN0KFneT8DVH52UQ7/BL45b
0CmzWxZ7Tu2a9iv1JZlqy0/YKHbs6Qovfa/aOlUbeVFHKiAqI5DBXUNuDJ5BBTizVN8I8YTQkl8c
oI5h6EKZzBE98Kf3l2NsVQGkoI9aZaLtaj8gHZWToBuAEWa+YKVSIh75H00vQsl8JGzyAHkiDTP1
LD2sjnWbuhU/h4+RAmLvpZ1gt91Or/JWJG8YBzh6ogQHoa1by1QVAUGVlZm0mnV+e8z2QhMv5F9a
PUMVZV4/jJQ3xuYDUnPK+f1XZvXvjDuMFOpe4lnx5NwiM3vQEYocS45gtdy4ij9UlNdb0BpGsw+k
ICchcFH/aqDigeC0E3mZP7bNCATnL1wrUX2p84EMZwokIOk359I8D9cvUcYlJTuHRLMlX4p3HRvD
0slUjQkkJBHGmafsePsYbC0x9+O/tTMjIogOWeveRfvEnxJ6Mabo7Bl3k/I0Ns+5aoMhQ94Y7lwL
I1iOT6aSkWY+TNT5bxqKfRM+Srmb2d5rspA0z7te3XX7FT9h19BJ+LbXMHYmbr/x4TdyZP3JJx92
0mnz1ViqAgb3o5+bA4ckZTWtkJ3SQektHmMGedBtuBW3S6q2jBlKpDMd+92FzjKoSE+LykD7dMC1
pfRxuVI7MqgVW9ovUCSL4q6Zm8Pl6KErFPI4IO5vb4EY2Fn28CTbGvroB8MEvvnb9TbHkEoDsQW9
VHP7HmlxOBq+L9bV/cMPndGyndxFmK1YkVDWqxcThuiiflp53TKuOcUsnTPc0QisNIumJ50dYiA2
Cx5S0JDYgkmS6cPtjZ5wcg7cd008Opotd35x2wPx8c3i8GALaSENBy2VTmqcnWZdGLDcfi39nnfB
0bO0cegNx26EngDsc8BZKJy8RyYo03DJtsIRX9Pi5PsdnNTsaJoRl5SV7PnE+sqLP4DrWTZ2zPmM
/PldFfFGLB7rOFfikoi4A0Y4MbHuaCoYdTuWxeyjC5VdL2EgIQ+/TUMNhEapVjiNMcE80LpReAl2
StEcwNHjwek5n8i4Er9N3j/2Eht5gll2N1+5BJX7zAvdtDP272XugHqexsvPY9d+P8aa3qgQHso1
/i1/wQO2oVsXRQtPGQN6qnJlF2uMOXkZnhKSViQ7xJrZoRL9LJ09T6ZBTMzlbLOZsF3pN1M3bm0h
iu1F/X5Laa57fkbKCs4ryrpZHo5plEzlR8veZg5TLSSeauhhCv5aL287/M3YArQ6Hm3y8qXTgpSa
OeY0NbOGsLKlea390Jd2stfjrDw4CH8EI1slDq2jb/P8EgYMLW1gLGjv3OMuB7DZa8nW22xeai4+
4GrAGDroURS0wAs7RXYXMCnHW+AoSRjvTJ2rFvcYS9gNidPyfPyFb95LCtoXWfD+35JosCb5DXmK
M85YUPIc2gVrqv6cG8/GWLGKl4K9qnAiDj9zcQMqT0MpYj82Mv1xiBv2rTcYby5W7gQyTXKYVLAo
8CnW7XZaRJkeq8SZKDXEbJwMMwnLcCEdeJ2oLhrf9jl4V0KNWoTVTbYk+PaQIzcyQAHko0HVT47R
fukK6kmTN8ZkGlu8EVer1q5Jve+GdXsWXKUoi7P0UJmKRuxCf3ad6GqSHzmMcRK6Gf/sFTR9aaRa
DkJ3mTpNJZzLIsAWm5q8FuuWvnWGaSY38wlVuiooUZ5njR/J2AnoOI5NAtpmdH7Wtr+mVVTpI7XI
jYfxpnN2X9PSoqgHOj+m/iXkIX5mLHPy7r9dJd4l/mTteq2j6cdTADn4+gJ2RRcWCCKrBpuXmcpJ
4QTfrnJK2+zQPXMDVmcpkVupyNoRCHGjbRRmb5FkhNkgCAsePF8QlsrFk+62pqjPU+MtpxUx7ODO
PqP5ZYNahiOsjSYHdUcE1/0u5zUnutSCCs3m2orDmsIPUaiZ3xv1CKJLqRmi7vV3x25yKZI1NcnP
9gUfReWGcxs29PqF3pMKJ/y5Y/x2MzGecNLXbiI0GKZa5Vk0lwMZy9M17H/MzXpley7WizS37L9g
fDHYFlhitOlcWd/F//zrtL8TJ+6qG1vj/3rnD3yWwh6PllPu1HBMAqm7kcyb9bDl0Qs+DNRhyYSh
RJmARr9uAV0koA8Q74ACbrvB9cUtzsA98CKoLnX67y4yOBDr4ENAm61kiemZtNqdycQKcZYLfso5
+HyKFVHB3UXoxjdqGBSbdAq2G0/sovwsbnTxrbJowZtQ1TwWZ+j5sM4YeQ9shGo7KSZAPoGhL3cy
ZiZMxd2ZFAKHrbNFCwE2RJ5Qg+Qt5g0Du5dyIHwnHGROPdqXPa5EHn9IZM1YcPsNzzjcFiM7wqnc
KVOJt9KdqdeCjVBW6PKlVEOo/K7vifeksobXofDZ2wo3m+xWbhIpgXqdBJh9Npu3wsaOfH3/j7fp
uvgPfy/6OV9LimOy+7cmptcoodtyDKshVPRNVaeEhPblYAQpSUslbkECn9qYTCnizFpsVJHIiKjo
1q4T31vG0N3uIDlIckzJ8I7kAZDDQuL/tuY/LekvUqS6UKbuGsGZE6IbSaN6068QkQoEENVjsVy6
Gc2ybcS9jcwgwb2R6HIBmAlpYZLa0KTyNQfHX/8OQo9up83je2+vztE42ZNsffv6bJx/NEbZ66uc
cCgbIUCxkwhr3NzVdGJVqCCMS3opSbvXVMboHq+K0TnbI1ZFivfc4f1atHpve0A2GruHeps+wBen
ZVxMJcRKXgqpE/uINk6QpjjPSBgRVuy5EbH6l9emOgbt+z1jPw9agMzhJ4FmUQzQnDFmSeJkaxjT
k1OQaXIvI2/e4ze5GB7IveaO8+vLqOa/o6/CTZk8JG8v11QlpFgeJIOlJt61k9eD0U5MRzlS3cL0
ticC7cJO3wywg2YZK3W5fK52lN0s1BeIj2woeHo9zlvjDMHts8mbNNzfsgY1QE70x5i/iNbMNhCF
SVIzW9OFtwtcIqHChYKSy9L3lIiXGxdi07RhudVjLk/0CL6VCs11y1cfKGZML4TM35jC9P8cF2tJ
MyNTqTj5oQoPhXhbeu/dR+RvETydsC4689FYrPgl65WfzYllTBZOAzhDf1L7QH1b7DcaQTjMMoP7
1zp55mPDk2qJXuA7Xx6tITTJfNnzbfbl7J1Kn4vrp85TC4USTWiZinttUWGHreM+nsW5DZM48jYn
SP3y9ByYR9DLmun/qvEi21/yxYWRt8FWDQzKMQ6raoKCw9IC8QMNcCBVsMQRjdJJEP2M9gzDSWyu
FUU8sb73sbXx/DrgCp3SHFDUZ1in0Zp6UctxoLgrdOxTAv3qeSGF1WeWBTet5ksnSaeRxXEirz+i
4FjzQcvnUHlokhnfPKh3u6ab5UgYd9S4QsTd7FoPWPYt7AXNffyyMv7MQSQh2Rfj6rXjaCO4jip5
J8c5M7aZkoliIue1sOCSampF9UKw3mTF8MR7Rq7JwDhkxtB+Hh54SsNxZ/yISjbTDu776Fmp74Nz
qwLRQmXCqTyZkbgVsFPyyqHblJeMCZWxHElVwqDlPgC5a9ZyvkJRUaGUynZnzx3ABviZGhPcfNzx
Sfq9HDcvkkYyRZSEXLJqHr+nB2Va20J/of6Y3RSTS9aWW1eaSBFtKhzKkNYlpdQa/PCgBL6g2nSc
5m1gkGxUptA8RGRJYF549cP1BH8m/d9HRd6Gv2t+i6eRv0KbhnHu08jdyIeNYy2Q9yUrs0y3b5RP
VUPy0jYHizLBZzCEgfh0o0igC1BZnm5etn/8Sqjphb37ReM3Midsm8LREp8+pcvZ/sEMYH5umSid
S2XXsh4KMWNItOHZdlT0lSsS9OBtxIOEzQdYebFntW4Tc75JuvuFPGzMKYj0HC1s72nbMlR8UkMA
BRyBG7tPmteiFYx8ZBZSJl0lk8QuqKf0EOsftP64pt9t0wQVS+K4CPGQ+NFvPicxr1nyphJAJrJ3
DbaChbbxWwFFON40Wnk5tB8YR5ygL8JXjOGPCW6VoYVeD+xRkJkDF5e9873Ljh0NSxMAiQ3FwmT4
qFKnxfPDjVCO9zgVkztOw82CFyWsQzimAVGXhzDQdOS4zTvHd/XBqblA6UlF3fWjnXEaHzTF+ZLh
etdPdxfrcqEwJ0HLoXz1ovl/vC/UXVOFF1C3BLyAOZGeeprFKsidIOYUEd1NFj1mVAt9NkH6VLBO
1sEHF2ugTIlz7i1VvSkcBCd6PxDN6XN622ugBH0NhvQPE3FOoWCYq0rN7TLRJDZiWPM6+IrW+GRQ
Ol7wrqcFPy3dEz4r6rzto/P0iA51pSKz9dXpOY5qo8l+kMOXIhFHPExCmSyd1GFB35ifSbeSv/Jb
RdaFZNvq1vS092htURvr7yNhu5fUsLu5zi/Wg0tKZv1NUwEPr2nZL+wsRc2WSv4f37LJGkLzgx0J
3u60vPozDh9cQgieul+7a9NUyNVOtd2obKSJRQ2k+x/gacLPTg4WaMp8wfwCny/Fe8OZ0i8Okcyz
5t1jz4UfQOGNjkR/jn6NYBUQ4CxCj4hwQwhG4uEzj3eGJf3iPfq6Br9r6KmwQvJmZa8Vz86AybAa
9rLcFel0HHqIwls0Gno+N7fzc/k5s9MpNkUdVD/sJ9ypa227hK47u+9eWDvnQ3BIW604G2IuOqkF
eq82QcanpdrATbAypJ7cavTALBJ4z9WIwwjOUOHZ3RGiSM8kMqB+SxrG5ns0YACi8e2p7SGr1Nfo
rAHaWIXPkgsY4x0NwwVYDpM/e1veM0J8ULFsUOcRqEOGap9MH6H3LCOe5XqhXUnF5HqVWvzY7lwe
B1B7Kv1VhkjcrcTHC7wxCZkkUwxn4UzpmQ5qSB9JpTBBwogAhHvLOt9maYbYq7A9VWwCQ2KaNybO
dOoAIo3I2J0iwnjiK3ac+YmFpPgJGIufsdcDHGj3peFzqXcH3M1Hxu/W4ilSGZurQLeUyktN5s4K
edebgMK++mWEt5sVmB+6bYx3IIigE3oZiZMF33PpeJwQDzdP8fpIWFtJXaq02XXSpKTN16SlFzlS
vzemZfvCcqiPSYuFhgNxXKCSWGq2us3kv7BpmXKw3XfI6EuZG3fJcI4jQbOXtTLzvscz3wbARiIA
578i3cwuIskKIESukWC/LeZBmfvYWTc4sf9VsgWCHBYE1uCpkpoHny/DuS9usDTkPQffVvQ7bQzg
l7tYUKL4NHo4lNU1RimMEZgkjI1hSoO1v0GI/yuKDtf26DjGB2lphj2M7bmS/iskJM23l8IQyjWN
syAeRV8kUYvLtKS+VX86xhynH5H5gNWHY76f5Iwl6/Qz3PkM8epH2Pfg2LBfaoCk77C1m4T9vzYl
5m+5APHNCUe+o7c++uVt2HM4FR7Tg2IQ9bf0DVes7JU8LaH1I8PEie4PvcNyIDKvdKn51c/QeVMm
x/LSiHhSymvlKV6zi5PZGwpU54JjHy8/KLj+CjBcVfls99E696MJrbuPHy4g8PhRVjOfu+iEzr8b
MeeS0IufKXU4UfnXIFtfA/yJ8OPEuiJygx6HADQXK/NXINELu6Rp/2JkEzI09Tej4UV+AaFZfuxE
3VHtE9cyHP6upXcQBdzMFqfxcsztT4XUyUg14rPg/qLPBkdi0QnWJ+nmu1Bm03G0+xVZlgfkKuxQ
H/kOgGl913SBMtih1yQ7btgB8qgr3J/xufmC60NuuzN6+iA6KW77aTd0QejFFNr9PDJWow9/4l14
+i+WXwFeIdo0JDZH2PTBelJt0K/tcUPCFiU0YndJZRKcxUjUoMzEktYRXH3U0CzZLEtC99SlEM8l
gATv4We7pa6NMuJe4Qo8pgjNKhJSLBLAgSIzRnX4Ftvdtau97O23iPq1U6BKi6jj3kqmgcfNC2PU
Z5mBKRM1vqcS9MXWUVNjeEaN+nCCvxePAhjxMTxi6GW+eaw7W26GJN47q/jD0DLI2WxbOgiGDluG
rNcuhMX0NV/JAxHqD8faf246xsuNMijen+5rPJeBEHo86OqgPzhh0QgRXXUsbkIjzSSCmixb9jWb
YEJcpo7vLbOuXiiEok3eDirVOBXkUm2Kkx2FUILebmTpLbwjKUj66vGAXPc3yiVbj7FZYudTpQVq
UCCEatKBi5p8RxoWR4n9I201kEk5p3icES6eV6TTQyyyX/8GoQ3lXTO7y3jOpHoNK4b+gAI9MFoh
wohjAbyshW83oMInDUYfnY7mILyvQstW34t4FE6uqoZBii0qMmcH44ObFXKCKEoOJ1NvymHgk3yR
dYQjEYGUFXf2hEo199kMaxBiA0/q5IfCRHiLwyoVrlBuYSgvgZyzP6ekeuxy5KKN3nfDMovkpg6/
M2i5rgqDgTeh2zpb2AFAHrxIhLCGiQXTEQ0E5rNFwL12b+i2LBdpgShWRKrXwxFcmdQ+vZAfX7np
cu0ay+4N5CMqv8ZXLlbk0mMpYcVuk4CO7IFm5ITNYzZNQXY1FZoZn/rNFihZiwTamT/gOTbY9ssV
lgsKHhk+jgzAYFE3EBDMC3/3K7DO6W0wdAnEVRHGJpjc/ogxYZP2t+uEN5yguZUxsbEpOY9voOqT
Vbcqw+UBSPO+Wm4NoPTRzIZz5/XDw8KM3tHWdDOdaKtwdtKjmM+mxxydZ0cWxLBvIPUSKJHFb0nN
jdKmhFsN+DYse8Cj924chwdY4ikksOtD/UyQ40WyCV9QCls4uAHIokRGaHtwnba/YLYk99aL2RcY
NXsQdTGxJkWo6IdXGgzKDR/gr7PVJ3K5iH5fCogRLbIKFfF5YgZzD4fsZtoEvEu4J6Y79Dr2bh/g
/DXVPYepNBMsKemvT8sZS8y6Qi+kuwCjfdKfkKFEMN8yR6FIG/9V54foDZVuBCVB0Kj0XyE+AgAy
3Evd3L3OJ8ga5QscAMLCRyiEF3Qb7LeYS8juK3R1wLGjaPOpqYC3bpZg1W/HEE6qPCeNMJ2r6052
a4buheLanRbNLgnb4cndWSSyGPbq3VZ2+gtTZlL2vvav2z6zQ+59sizAJURAlL8KhvAM7cRIEIvf
aO0IMjHBO8Onfjj7w+pZgvYvYsBrRyJky02YL4qJDdKduSr6ou6QT6b2MSiJkh1g05KFig/oTUSb
1911mMaEH9uZP0qvc9G/sTjZIHMx8exGkRnjHsw1WFzyjoSnvum5V78tbuvvymAjyravKv3jzBi1
exa57eXo10NbO8Vn9+5uGbgYNB5F2BB6soWlKo4TTlj+DBvITojlGIgeq0D3ZuLn572gefUDvNN7
KJ9BmuPOuMFyc+WPaBBcsP9ZoFx17GGKMh1vtsoQ6IdFn2+WoensMVGr9JYGfWpvlK6hNAjJ2E4H
KWDWyW7617uDndNy+mZHiH3BeXsWqEpca08J2+wc/a9u5NvVU9h8er0b+o/gxYIueHZMtY8nt7AL
JQlBI0p7xGV5jJtsVY/4YZ6kcNmmafTkS45bUKEKjm1huqatO9V5nSc5b5Ngix02eWjfbf5qXIm1
yxuDfIic+opUBcurWpa765k7bfSqJQO8Q3drhXQ8WL3tjDFXNWi1fDhnxM+NNYlsgdfbbgt7rLd7
8uK2cnFrv8NrnUl2sybTZ7ygGDbsS5f5pYz5zF8YmNwUpwniL9MUFrF3K6vx7HFDUuKmpWQt328n
SpVARXSNlKB2tEVpCZopnmqHRbFEwqHHP/DIrKI2qe/CKsk4Tzpcl+3n15a7uuPxbUUkMU9zZ1A8
xHoTAXoZJE56N5WOYL9iORkW/5DHZa/yQnCErYnXk53wTydjrHR+dlIuzCs+oG5s7PtGSIjTYBQF
EtLeqs6155BUJ+YHu0CWKNhJ0yTR0hhqGQ3w0AROegsUC+PyRbrJ9Ckh5aXACaEsAxcmOAqpkxph
OQls0MQ8t0GkC7LVkDoXbbcqOOwI4iRrHqzQT+sZbHasQVB57bieL9m5V/UeUVdEi1kXVlQm7chk
YtYBqdQf9190TScDR5WY1PECJvPX0wI8Az0woYYZd1/uQ19zS5rgUre5IMoGKdP3/VQZ/fSwkxsa
EJTA9v/M+tjd6zLNMVK1BTUgdormDDDYpFgXjdWvccEKsgn6tncLnl8uB2ef5c3mplV5pFLcm/ve
nesaK5Y7Ep6fGY0IFNGNRIEVBR/o6Qo1yRSVGeS9gYk0OgXxfbnKY/jg6pcZQpFw98ULYGbhfGiJ
azihTfVIM9MIhZYH84WCXrJmNvEFyH4L7JqnTadO5jSO8iF8LGCrkcX9ldXmqBpSZ6h4gvzQWsiA
w2adC/P2vc4y3ZjbJqkoSAKGw+ccTf7opfx7bg46jU8dlV3l+jYhQG5vmSPykC9fDdEc1fTOo0uo
hO7A7xjKoyaQ5KPKdMeE9z0otnCC796xheSXTyntBxi1FJK0fWMuByHCTXWmfgzdKncJYfHAhq5h
Qsx7V0ov/KI2imlGADowGSwu1rmPTvQwen/7XIXJ7qcsJL0mW1QAyBvB1GYtxIWiBqTfhKI1uY2p
90CNoheXMVR5iCdr5S0BLuh6/9hHYxdXH+wITSAolS7CJUnsNKI3lTzXH7FEEq3ri3dfTzuMhj8u
4T+BTvKQOi/wtNCu+LlnQnE2zm7cUiIG6rntfhtx5CB5SuUjJOJ2QasUJ8yVa7jBfYKFbFhRdGvG
3d//0R5GcgeK6coCWKTGkhT4ERLm/+dropLmEJnciFOMc1L7EXVMge+fzU0fYcB8s67soo/Ex12+
8WGw/b3e9sFXWWFWN4DWUcYKDgIF1qKbk/bYEBkxl+C5Ax2BN+ntqi4BXa7Ya7kg1tGlSRKFzmCl
9Hd1JUvfCIoMe9M/zjEzVnpH5/hkksiTet6qtH6+bP/h1xaiJ+XPD5KtzNw3OLdACS5cy4ZbK/tL
0bGsXAFYop00depS/NrbaDtPQx1X6lHhG2ETgldNVZ0wcb89uakfegBFXZvMiZAUZOlOM+sUl3Z/
3es2iqjuzqzSGJuyaF2uCi9YVkvsGV5U3ycBrUTdJQJUdEk8xNf/igknfJoTzNwAVcsR8hBo5+qt
zGmZ7gpJ+Trtk0spLqI3yiDuXylWMFamB+N6U+DU9WDi1+2YGwcMNyAk/8CR81ixFPcFnEWN0+D/
0InlmpI+ebReumOsES4uOCHWWCnieejO5O2W3aHSA/9kmBrU2Gyy2RUyQBtTVKUvTcf87+ZNn12g
VNzrIvNI7DB4+Dy0kBBDdGStIozOqBSam9dwY932JNF73m2BB4xi26KCaZsiA/1jmamcgZ00qSar
XhU526bdvI+45mOJJnQf9/Bfbxmy8JKFSG1ooSVNV5ECUciA/WK6kBx94j0/PqRjXhV6xSUjVO/k
6eNE+JQ66MnvcUm10EMw8kHqvwkwWP438WuaZyU8vSZ2vj/FREJ3U2330tex5rYf96Qjb47t16M2
NFoOozrjqk/rraPSPbhso0KNSn1zjO2tlj5nkXSCpOcYY1q7GkQaiUGFII8jDUUF5R/PEC4Cs6Io
32y4R5tPUPdKBxu/SAhITBm1ZaRnukaTpqpMqw1VhqHqZYEjwB6RkRhjy9wNc5MDfM00iakpfpCe
VeyyDwM4ZymivFFvtJrFFzVIThJYceUS13MA7bRvKyjHbp3kv7ubBc7XD0XCfObElh20Pun5O//w
3mrVvvOb9ai5gzvjNkTWiK9CQKB3XPWgy0TomSPcjifwIfTaXHVluoHrMbGBsTtbpyC0lz7mX2Q5
1RdmXjZRCwkiq4veH8bF4kfOc4Bx+GFWlX7YMr56Xd6XvK6BV50qikRmg1xKuZkLJpKI4EOJ5VXx
CPH0b06aXl6dN2l3l6bwFpyp7ZyNGhZxnvdPESU5uqolGBbbqsll4++DfRc+nBOor1b7WDubd9T/
AJBvZmTF0FKxWwNVefj1jStNsWYw14wIIaM/Kk7vQS5g4ustXyEhpHhL2rUG3hKGqsJvuy5vb5tu
CDXzJdXCs5kkJvJ7RqDPoBg6MyO8wsVTMmoL+fsI+U8qH6bjjmP7HhUJz8fgSj4GSM1tSrgIvxxj
ZLkwL3XddX7FYiirqz+1o0J8i9qXx+h/B32ePOFez2+PSNoC9KI4Cj05KJiKuNAqs7CtaaGlyoZr
cF9uHpkhD5jCcK3LWFuzCFFsOVpSARcPpvKAl31fkeIu1qgoA1JAIrf6mHOpAir/Mgct4HhmG+dk
+3lFtqLwjjhPhLPHlXm4NzD03a5kfHxenQygPWPnTMmfE/gHggw6376ZzUHzKcni1RhSHBC+RnUC
sTcbiLYQ9pDyTSxvao4qZQ49/kTMINE09e2oImNwZQwKvQNUoAGwe4T13NU2azZURE4s9cqfVvv5
Fva7Rggi2SvcGvT54W5RQFul64jIWrLb+HNsQ9WtqS+O5vknhs5qLMsy6EXzI68TuHX59JDa7aVt
dEkuumnkuHcKBzxLpTu43LQ00hC4+F7mRb2DD91DhkNMtIu0firlRQmO5nUXi8eSsuCplE53dbe4
ZKGzBD/sUsPugAqSA9n2xQkMZKsrGd7owMKXuOe6/Ae1KMo9eVXLqYp9Gq5kPw+6JWS27kdm4qGs
RZvo9jrBCU242HazkT10xrrtGu4wYnLkDwbVGbjlTt3EWduKsoBPkaCpjVyN+ikfE19oolN+165e
SCvZ7iEAfL0pp3sr0mHGQtowccEULUW0oDSf5sGskqmr2n7stNRxOTQA/PEvzMDmDLXUAiYj9odo
hrjJQFiiS72ANCfQueeyUb+DAV0WFsP2veP9emSR9W3CrO/6Szc/CbT9gjrsckfzy8QgI/AH7PxG
06OQSyI07TTAR/pEIbt7+Jme8+57GXTTq5N/mhX532sLPahKtYJ9ZmSTgaMR0viILVVNVI7sF+dx
8EWW/LFOrsqcuRRA8Z+EiiHGo7m4QaH/QK7zBvXgKRltUh8AuUsDn4uUBzqjL/PYSx3W0j7rgByj
kOtaBxn6CZwbLHMBzTyrYvRaGQ4ZJYvHYnAipddbBVK+d9wgcDYjuvRyrm+Q5enoSNHFkSPXRbBO
WCEqvmfsiOW3C60uUHq3fRHuETdEm8a/k3VSDHW3LoxOU17YPyNR8+BQNc8B0X+a61FnWbNY4M/6
9DQ0bZ/bPpmMBrWAkK2I1hdCuFxqEMZWPjjTCdNX6kMPvqDDyqPuwNGRo/3j8T9rAZtot1qHXm0J
ErZgHbmSzlGy4+/xd/i1aMhGYTnD0sH3P0ufvB5+73RTbAWX9QJtgMjKowxN/EweFi0cb7po4Iqm
rlpaye2U47ijSkZTq3nR4e94iJSUyQqqID49ZnfuXTsNjhyae9V+zP1vXHAMGKc9OQoj2PzIMOHR
skFWs+rfH3RLconmmARtCRcFH7dQzFupvZq591E0dcJN20MEl73yiEcfPjA+qrDcyCBXoVbp+Ebx
VyiNWb+wtM0u4pSixmwIC2AcXmUggSTXXTDkf6r7f5S4u9+sBstE66dZfKhZCJ3eAtTLlmOXZSd2
fOAuEatjgtgobGNcj+wuTIfvkIc7WeHOfb41daW2M5kXwzuz8p2VokQYpD1E5nMcDFZBNqAcHWxs
/bA6LoqvjeoT/zaci+i3UYuvyqVh2nhLvv2pjp64b9YFgnwt2PIhX03inUJopP7H76dv4I7+yJ/T
Wg9g+4PlNkdp3LKActjShwFqz3FJc8rxa36QE1CVAvJrSyy1lFRdMx876OKUwvSfReIW+/kmnB2j
FnVUFvfShI8Fv2wULGxhzMqn5KsvOXQHPyltEkKYcq+Df6ue/dRvpZSfFsrmXI4YgwFnlr3zCu+L
jJHfBNMfhgppv95KF0hnMU4WbiKFv49Im9o/rCtX2P4EdxzSJw+Vl5LgEEpFUQCMvK3vsqaccXCt
cJyc9ayAq+NcWJsxazgqd5rLly24nBBZoZBtFA7+9Bzn3Rtl9pDfbslf6HEeXuZmxHDXlmKzdg61
ekaE4AOQ2UOonRvsMxSe0r86LnAlvZ2SnP07KFn9ZtblZ42NE4D7DOP0XmqyCUnjI/mAAqzapTZh
yfnJ64cvjuTV402M51qUModrv3/qxc1O2NdDLQZ0EaUVfy7RiFrWRTa79O2tccnYEQlO3PC2K5se
bdDG2HUiqEvhY/RFBKiwCyxqAnsQfACq970CTynJ6lMIDbZ1nl08yIx+VN9EVXZ3ZVUtS6LNfV+5
Kmx3kUQC+vgVsX72qDx7LsXHXdV6Kgz4IC8uU5eu9wSV2SN3Iy36Sxl6wfSZYs09Pn1UtzHGo6zZ
+nMzmBku93ibVWyYol2ulq3dffKUr6fvXxG98jgyOI6rHiYZ7MVzpvB0Zbm6UW00RFaYgkOtzrLN
EVtYnQij0M6w6a6EX3ZiiTClVwy1hJJyKxF52fuXdAQ6hbhhCMKqni7iOqEtxfoDtiEN/rvvIUN1
6xVmtNG+1EiBv/nOVmsaQK7Hpjw26omDuevWeUMtIr4MqI2B2w8bbj7t5M2WAQbKoCZPsouKh0MF
iHBOWBeRvOzhDUFhuGhQPzuDc51e6Vp7CnYjutAaekCBcRrFsGcMuU5UWLnXIzie4U/avrq8yqX6
XWUDezXL6tpsCuIWwiPHhCuAJlw+VrxY0Z7NKE7vmsXC9hZa9ahwUBEea09j5b+ZdXMrZVlpUFwS
b6r2wJPfjRp0me9TY+jrlrw9B6cj2N59yck6/k4d9Kfyjy4h1i4Hn37eXLY3HERnyIro707NP2Vy
//qZwi2OoOXUqL6sGVZD6h/794gXbx0VilIAR6WmbKFs4woGCsWkvI60BWWu1OS7oc3FK/VF0FgZ
ado9S+TaJA9ERvZVE66zwFyK3NnwDehw3HDXJTcqN1e0HeGV7MOcw8UsBY6oVVhwJLPrKxU+nYem
3d5+d0zEngno5YfJql36SVG1LoR7as2NhXD3LhG1gov31RAjUSH5Lxd6lD5DWVmKV9Mq1T8GLMuV
yQSykFyRrla5wuVkV/DMRXGpXQYuZDf+VsvbKM04UAQbpTI02w1G2XOhUlrAW+DmqQ4zTqPjTVO3
Nn0Rf95vw1zHu8jV7V9ku9XXTUDyHRAck8Jgze0pVN+YYaMr/NHopFlq6YdlfrjnGK/kJabLB+2R
IkIphDlK7repmOpRc2pJRYMujL8ANLi8zZuwSzaH9/4q4KTiTiP/+Idbuo0YKc4Tgf6D1y1RDM9t
b6G2R1zLTqjK65La4FDBar3CQHxEqZiIPP9QSHl7Oa8DkijbPhJmQxWaae75QNBqBNR8sjvtGxPz
HeLzrtRB/eHlQf7oIjQZ4T1sNxmm078HeHiHkv8Bm7C0WaM7V+ppllzinhL7Ft6N14Yltla89sZD
JjfnIhAENv17S+5veDZUE1YhhywRcNpXPH/nbvkQo95y/2b1ef4j1ByIpqpcCTw+fQr2tMwNHcs2
xEar2oIqivFe4zgUNuPub7Bq98KNlT7O9GcGW6+jnL4mDuigM4J4maDl0xOyGw594fzqrPUTA2Ku
OVCjmFv1n8pErKtK+M5Btj8ONrQBORiUyUshI/5R8knEfctJGPM33X0WYMQAhpHPG4UAzwo8X4Pd
xPpiSpie0JSWCjsUW820w335fw8mMza874j4rngj4XAY01Ty5eZRT7P59AK01TSRNtp1Hm3O5Gcb
fWWmwC2NYh8xI2AIxfjW4VcjbsBh7PAvvPI1yjsTGMEu9CEGfybMa6z7zYM7CRqWX6mi1iOfpCsQ
vZlJJ7NUfxfEwPWDuTd4tp4S4vA1m9Y+vbFLOwEfX23x4tzNheHAne1q3MPyStqyd6TTgTSuJvsS
hXSZXvYDIm9LuvLb+H6ze1QNPSd8jO7DIGajlVeTmDmpVDvD7R+Lfj7ytFRyCF10nCtJ9rDN5+t7
WRfziGTzGJBcVGlSqPoc3rHW0UmxQEsczZEevmabQvcSNlZ6ZUDOIxv0mkNmgEt/3LXDwpRdn1Ya
NUq9WgrDo/oDWkTf9+9Jo8qkT4WojD/r0ppKwK20/SLSH477jkdz3k6w3sIgIUVpqJ8/EOX9Qt/2
/B9nAr75Vv1NxxVU76S+TjRkmaHt8BXey4rJCmP+Qx7Bg0TVJ8pfXYbZiEn3DAk1sr7CavbiGvX2
35HdTLO2Leiaqgvm+3Lg5h/HwoNuEua7JL5Y4IkhJKtzUvKxPRCdHH60dOz3tRHAxwOXa6fzgTJ7
ts/1Ty9n9LWYB0DYsSUjG3JyfIQjXAXyyUlQH+9ZP+q9P33L8e1JF+cL4WUEAzAekwEC6mi5kMBX
K2QC9M9lR8fB62af1c6awUcTrVBDpdmCsCl7kO4zStkSKGrpDZ1AqGAWCYz16OpzyOmqzbuBQ13Y
IZjbHHlQRPsYeaRHKAWLq/Sh7bfoz3teX3ZhmgbNnvF6b/mY3BUtoS1etI/MVteo6RjbSgoZM9h+
LBZq+o2BbVHVnqX77Ul2J3Om1jBGQFVfhsj2e7mc2CGKD1ExTTMVApg5D10pydOiFNFLOI0hCDN1
jh5gJZd82Z1C+RH7Q2orY138EIJOmpf6swSK9dkgaL4m4rsizUyWjVbFBcbyOxSftqoWfp/NZOaY
KE2KNo9NAoNgnIbkxvNA9kXOqGfm+Cp9cWOHgUXRkW4qrp7Rn65cF1D8STEHZ6mhMUfwiekd3EFH
2yZdKnDyg48bhZuCwWZkGbslDD+YWN2YfkWEhsYo1RIo+mBRj4V7QA4jgUcIqZi/271ampcLpixq
M3e79WxNyYsWSJ9dK0mjjCmqI66W7V5/aj5vo44stx3Bmm+cWtlo9nHKgLekBTzmrslpD8P8n+NN
XHJ0lWoknXOMam5fbZ5iQuj6BWaBJIZpxSu/oCHm4ugSbwx+sSnirgPqmrnoMpMGeyWcE5SKIvYr
C7T1PvPdeT14rryEAqfcswO17VbhoVw0dnoZbNbkPn4M1lgSZfkkODVY6LYOI9hDxjmsGAm9hAdf
0uwVamUkcFMRirioIOjVYbScvEom7Sr3jlQBSNqSv+dOMQe5ElFVa/5a7ne8DfUrdAmRBY8uLb2O
j+UWEORHwyyqeuS1auP7EnGwRaU+8D1Uo8GI40rV/KyfTl6Mb2NrM9NevFeGuLIOVIdkVpdIU9xL
7FD/K911jzb7oahZToDs9gzSUHjEsf/ewtdN9aBVY1a6ENui/r2j8umPzJV4KIS3zK9UNF/Cy8iX
FlzXTbIKG+A5HfacYhS0ua9UkjI8cgzIo/QX865NOfcpRXTOe6lE3KZfeWxCdDioyEbCo38nAf3B
c3qVU9uS1TNYwKCH0rQfB43mf6BDayp22xs49SU+Sto5WUyUMC9ei3WrZXYXRmFXpBqYt/+PH+Os
ldHB9qzqqzcFksbwTfsWeHC5HLEtb9JULqzZPVCZ0/qxeE3VLBNWCXP9XD9X0HY/mYpn7nan+UvS
5/UkqQS6T6c/hN74fyWltk4PMeFkF2ZelDCJdMiratWllBxwe0Y62Zsozngc/HKl1feuJ76/tTDg
SADAcV14DZmFwlrgT4KTm74vGdx6OyOo7ZB6HE0Z3eO6aB4t/QvYVkTuHtYMBmB+bEk84uFOPW8l
HrWvPvDaYak9t9HdZMyBqvIo5q08m2qIY0PP03UOWFhpYolodBLnYV7TWtDWd4yAgIorlTbGiroi
R8z1cf3vHQ1CLtFE1M+/FViHI3+bIPO8bQ2w+lz287lsTCuf2d9JeZG4kx575FbccQ8wiuHocAcV
ZKX+Dr1LyyL63SlOhGwmFyxkKMAyMZZDVg+6bDhRhrzRwewMyVPQZZfNy1UcrCmrgCJ8BG0jAwhY
scT3Q7AMjwsiYfcRPnFNBFwumvSbLKliM/4dsWibHEZQUZHaBFtC80EZj7Hdb2+IMCVGoDb1jejY
vmEwgrxETCRLj1t8N6jEGJKAQU2z9N6yUbm/AxHoXo/B50BFgPHKaUk7Np3K1yxcWpx1seew0fpG
2TgHvAYGghL0dvnagfmAX8Mht/56pcNe+8YRPyWt1W5IX/Alt2fxUTjwyWZgJi2F9Ue338GVcKJ8
d/+bNnTuAryAf+1Sd7m+PhlJ1lG229j8Z6jg7brIKQI4r4Vs2eiaafIkajT67vy6jr5w8eTpUV2L
XPqYVhQHpJlO2l8LcCOn0a05a+FdpVOYdnQ8Xi+Cmo9HtUkQ0xy9oFH9kSR0fvO9j/h14lR6Ykqf
878gKzTIE23cilmqOhZvxIkIn55Vi9EObm4B4i1n68cJIx4hU5abCewFTMvMZa4mzWIkRE1uYqaq
R17BoRP1PkXZCj0LPIkYxW8DMnoHWdcSlykcmADK6gU0kJ8y3bxCIsJIeOUTR1qJpBHlSCMQO8So
vUsz9GA+UvIZZv67QX+HimLFFFD28sD0Z6AwHUPBdGglAuI0NIlPTGgY8qNgF0x+80Ng3HRbXSkd
F2eGSVw0h+whpUMAcA3jVezwk5jRw2wQivDSWWe3NaWKWmvLTRRh6BswbA7X9fg544B9JpXFS01/
Ec1lHSVl4VwooM/AW6KSKCqCIJ0ypyx4BHjPwqVNOojwxq2Tj1ZRf8rwj8wsSwPQTPP4thiIXyYl
8gufCC0f0G7SGyPvifPk7Hng8ZFc/tCjrk7ZAShC7BeMU7XQwu5oK9tZkGc2VoiVrWiZ+36Hd8yZ
ASf3sy2r4FyAhDpaxEyqrwhT+AvTFeox2Gg4YQycBSIOX+ktsjONb4jyjo47W7U3sJiMPC4WmIHj
lGJhzFQZ8ELkF2sfg9aymfmy7/da1/VpCqdIdp8sgkqGJSwJwX8+nIyJXgvd98qrLm/PE/18OB9x
N9cWXPuFur3x+3cjBwKMGrzCo7k7o4UB9GOaiiT+Jh1WMuKeiOiLWvKBzFlaGJMEOFMzLeR41yvN
bBs1SYFbWZuX4cE9tz69gKuusd+2+uofeEb2vrKVi1Agtpg3j5WLP+c8RHrR7EZRTAQT/n7YVBgI
UponS0NG9v3g4JVeuKy2iI21lPKoWniEEsu10DNtgn9hkHXzFoMlVS23SMXrNHfwndGs5oys6R2G
HungOHJY01xTvvnj5jWdoPb5rOvZJy2NlmI20L1sS1YraLMpve8owZGloErKb3wEKtOMINeRCLd9
1IYPpc+Q0+Z8Sp3JN81DFhfe3CdMpZ/tyOirHYqK64hKK+IUJsnHv7nQloI1Jgbd85TVtrGtrA/U
fjVOO0fbGV9lFHxmXrSrTnYstWdBrLmb59LnwiU7h/JeF2L0P4O9HeEsi4UDSYaVHgEyqKmOHbzp
EkCEgzVimrOg6dvNyzywUC8ojCnKLPo/T8M52Sk9VCTX/F2gS7MvBO6zi0p++O9r5pQYemnX8/wn
64PTkIZ9L6LbRgKXibBDuMO/WPBoBqw09c9ts7tgQufQh9CVtLujwauKYfyHip1iYcZHWic1joqc
5uLhomFbKwMpNemcrD/BDAAt+qdhIOKHOGM5OETEMtPVFe5Zl0Tu3tLcUOOIMl2h98mm2G2ZOP3F
o/gMRln7XOKInEykLkA6FzkeMBsznFn+jqnJlpQL8XJ2qkpjGpnJzyW11prf5AW5mzQ+3zIRa9Mf
uLwW7YhYroPM/n1PTwK49g1YmsdJp6YMGAqPvY1x0zVQiJnotyPOH/RbmZW33b2L/KDPQLz05ymS
+A5aYAl3ziF22Cxro2vKaI/zS6s6jEzVBc1P1qalRBjaKXEmTpSDHLxm6o91YDExmkDuZn4t27xV
AFENlfr2KzSU/ejVS40i/0OaZTFBA7IN7SCZcSglaqwYGi2osQ14996GN0ymhnYCq4iXY1MGk+YJ
L43TgZ6Ne0BOrOe66abH++Jfc1LrGIsmTWVvxZ3+Rteu9Y11KhL1BCJdlEHAO1XYwb/EGVJow0v6
YCHkChnxyFwzf/mIlvNeRsntyAGwGZ1WNeY0bs7oJ3QKNml21DKyRB2aVr+/yj+pVvxBcFXdKxM4
fZKzuFMosingcd9Glx5Q7aHRHtTtXnbX2zxYLAl2PrT3/Bh3VtJAfCGiJLHDky30RD4a8ng/c5Z1
AR+P1w8+Mi+W5yobWijEe/WlFkGre2Egzn+4EMfgY18N2Djm0TdQyQWbYKojqvFRSNueyluBqOWC
CKqvKxpFkQdiZR3KUX/LTGZnbaNNGdheJhzMUo7iixpUok0176tyltLi77xDaVC+feCrQcPKzYyq
DHzW6LZV6b7gd8lonEPZpCa7NbrP0bSCd3dxF1mHiyaQl79iqGbM3Isc2oP7vn9h/JfCFwy3VQW2
EA4/64Mpl3/yeT9Yf3ikRnmksCut6yXlVk4z+iYLpFmQF+t2j4s9pjGKUD77/Js+F2lYMKGjxyXg
GmLzD9zQLpH4jDN8juhkOP0Cm8l2LpOD83rrmU5UX3VFWWkTYAmlcJ6ZK8p/b7k98IyOicqwwimX
+F0a2fSZF7dk+lAPsodBoXegXlN/DzplYLFf/0mW6FCbYIQCboPwocHaiwLPAWNMCR7q8qYRuM5E
XZ97RuIMVwmMOxa9VepSp//DYipso7DrpiEKK43U3BoXEV6zgbF9WB61wcqllQw68Dk5KDqaB/7S
o5eDzkaOdg8eaqrdunDPaqlsMQtU1+4VZ+shgH3NkESAn/XCwT7MoN93U86dhAOtKqDrxzj7USXX
670Y39E4fBGSkYhI5cxBITVmHWRBZbl8FByaJGPch0O43RSolH0PGi9RLMXIxWQ8vHvxlsCHZYeZ
XXazoM9F3Pnf+g81LpEciA9ZWDQLXL12U+yepzHe4EI7Z0UXT5w5OxodlhmC5BMw5DkmiU+YPNTR
nS1gDkoXJwkF52MLdLJ36Ps9OdDJuq6Bj703Nkq02TKPi5pk0c9BBTlBbqlIb9NQWqna422Na15I
1N5rOTKBetuCntrBPP86oHMo7bTnlWfUlJto3AOpSKWkU244fITwFfSfaOLF8RhWh0hXmCCfBmiK
wJ3bQPiO8i+E/eDmokXpuFEYzCIkR1ZgAx6CWAY/kF4Rk7JBbzqbSYyp9lQjKZz3hiKmF5cc+Rkm
Up+yG8vEioTtTbCVCE9vuLPrdSmrrUnNzabC70fsu2+UXI1J1JiIpTqtPw29E23boE07sgMY+s1W
mKIR3KL0UNrswCHQT1q1pPa2q1y16uLwCHRoPhTMbBbG0pOHYuaAQMwl26Z0S1aGOD/QmH7CxSzc
XQdn0Wx8nfoEQxiCRTcrmkG8DsSWdrkDJ50NAqHvpEeDgQxJWbSvR12ARSK/YrD/QDyL4hDMEaLh
izyOi8cbB/KRj0DMsrd8WYCKR8nzcUF8AKZHGz4pm4cay/o2MKOC8WZ24KUtTlEYf9mkICjBvXYh
revCU8hq1pujUHduvk2lDoEAw93HlucDjVz+TLudrU4x45eapnkjzsWYAhCu8GUFQlgb0HYpSPyd
ddS+vRaK0LpWoW3/60kBi6bE5Nafc9R8enzx8C4pkNxck+lq4XNgjcRDxiHBkBBbxULC3glVQkHr
23lezddRkWkUHIe9/WyqbCgDg2MM5v9qe9Xa8Not6ujcN15csqVo8pft7LDfLOMB3uTH9GMg5PtM
pQlAAF3ZsfC8aNqwMNDzgRP9VT0rYDXJy////zI1VZTYNWkDCNoCG+UAdFPYaT+CNglX4cEyZRfp
1zSIF8RBXtgt/TmJgzNJT1+uIlrOe9RVeTKzR94MkAGWVLWtF3ad5mQiDrEWXmJH4xvB6XjamSm7
ZmL/paMQFp2CGZQPcJK4ZqkL8Q28AaQxvGRjOntlygLyf+ZzY5VAxVvuW5onz6zuT07N35f6txSl
EHAQp2sgh514ULTtRquO5Wk0QiCa+oMx2Ld+XeyZP+ZvL/Nski313pWJ6envBXwII+DcM5ZY5j3y
ShNe8Kzj1g17Wuk3leRFAXR5mFDeOCgLjsC/aHjc5t8BxhdO4KcFzjrTPNzQc8zajsU/RMP+0cB6
DJ2qIkGxWuWmAqowDgy4p65MmYPRAJO9EsVnCo2euy4vdokYqUPhgxm+ztEg5id/cZOTDOiKAxV1
MVejpZLQGs1U6UjmDEUlj8ZVWWiEZ9O8bK/GMvHEQgBrcm0s+44W3YjkSPkQcp1tNq8qOL8aPijr
I6MZFbUpv21ibFg9M33v/INp/kazKWKHyiqyOdq372mLd2T/ZVFbSp3XcmBmeRdNnM5Gok4TmCuk
uYaeC9WLXAwHHiCNRNq/8xdoCQYCujjW1UH+/mvptSb8TvpbfrOXtg5auGAQ15WcqdPLz/bRPSa4
fYpcflGGq9O///fo7V3QLj2Ad8xu/EaDromcnhTbl4Ol2qTrA2ugYy4ICuGswl7SYI5yutgPALBm
LYCKfQ7V6r3CmhcTTCCQhcgBUrA5lN4k95YRFkBikbYP4tL0TgU8yifI5BX3o2AI396crQ+PeoC7
qp+lDucZ9DXaIZr/mjY2GqDfKZiw5qHL/dJqPip7gr0eCbZfkrsxLFJYJNfslQv7xFD3vv+2rCzX
wq9skPiPO1hLeIYObRmMiPeVGE2GKGpn9Bo6hryF5R0zSGwMpulHv3P7dueHu+xl8yrcVvsj4LPZ
J7xHGhahAxTlzwMaL7C9nuUfrMHrkcWlq5VCTAVHGFZfYFcVyUIeqHacYLbn84ywW061mdxjyZLF
NHf3BA8EtdzZIjbhaS99UUzsocoNpRVLNNMjoSrXtRpVw37RPdIsCZSeh6xfBN19/JeUJBJGTQk6
15WqblxUzWuHz9mz9xFOf+mj5fsCBTGittmdMckOkXouBLkxPz7bpMttEEs1qeltTElE1LIShffZ
rWoxzNhyEjv5Xs8VJlI0d68zYUZyxAouXMXb4G1PrHxJtGP/naLZwTUiYJMziNXHdNCvLMv00fbA
YbBREHNQZp6j+P8ZXmwJisbHZ42YYt8cDil/IgxRW6baOrGb1Sj0P1qVPsGiYv2BV+HPxVKeIneh
zYUQSP9ZQz0PK3j4OrvTUSNhQYvjn+3r5hz2cb6gkKmxcbZYsGw3EpQYiVrJiD9w8Vpcf74DDZM2
OKD73zq7bXrl2K2qLFECvqIdKfgHO0az/xeWyfJaniV5o+CsE3qoKzR+Lx/zSYMo6GnGl18xUiuY
/fbXRE3upk+gZJDNkSCi3Gzx5NBoivynAkPaJ4Fo8FH/LcjGpQ+EM2pNR9YknR/zHkD0su/RMsAh
SZOJO1cFChUMf+RJ3dMvklTeFp+TxEORykm+qeApw7ytn8egbN4TBIHYgLTkXoBdKUwFRBu3gA8q
6zvexPdd+Pd9qL1hD0S0DysWjw0+DQY4jM6l/S6PEwwwVUaNMjH+m1CDcmzD5NnWmOz4MX2lR/NA
xl9HSVh7GNC34eyDuYmrymbUaDa24PGK3fgxyYkeeo1/750hmncwl/n6Q2gnujlxp7OrthpMq609
mO7t4qBuH7UADhpUSuJBDRJgacd39yq+I9sDbGZ9GAg4UhV6hB6jvOI2dhWYilMHpett66DTapiL
xer/0kPJNERsEsCtCiRxhnW4V5+cptJC9YrNTJjgL656fiV8qITm3sztObqEqBlmJcC7ja/c8doN
njhHUTo5nG8DXXqOkCaptUuwj+Dt7rrjbeguQAQAedwH0VSHbFpfs25ia230kB0APwKO3Hygrdgq
AINmO+yrBjIWoeatUeMtQSbfk1ufghqZhEKULzvqIkO5ZQyqxiNeC1Goka9cBYB4xuIAsPma9VwJ
lmH3WOsX+hEK7ALiMC2cVstfOGVKjtQYdeKIY0c5Icybz8s+s00qenTq09m4st7WlPBAhqNowyfY
T1e0pgfa4zb6dMWWtynzn+RFjz7wUtTGRwXN7GSNPywLepzLi1Dpic5uy1XaaBXJKPXi6OEVLDml
Nn3CgJB1arLDYhA2OsUicMjdFdWhgJsn61e4hT6jMWVQvCqZF7x+5CryEvyOJSH/mUv2+w0h4QYj
0QQIAEKRcdnRlvuLdFcxpoIa5UDNAMiq/Pw1IFpeFYSwD2odoHGb1A4P8IYEIgCdtJ2jp+PDbQHf
lFFwNihvoLPxCP+SreqHCEI9YuYuRVxpmAMGbrCOygZKk5sfvgT3ZGb+iQSFs3k/911k/AiqSL8+
w5UmGxIZMwAqeJXbMu9l3a2xXW/BP+azExKkEfkElwkXpm4YZOefBq/H/GjKnwaJZiynAdSdpV7E
wWwW8KEl1S7wCyFJ322fQrxRuWLxCG6ZGI27Q6b9LUArU4pq+wyVEV3OpVQuoR05UD/MFsNSOu4D
VuJGLEUQcFMzx4x4MUZxvTIvreUU3xvSBaah19xdKIlTImDq+8V2T/gHxi+prEnapsf6uRy2nNN4
6FViEko3DkLfomD6y8EKV0Afiv070nZqJtaKMz0dRS7O7b5MrzO9RR5EEHxJQoT3rhyi3mhgz7Eo
AQsISfSkjUmtt53OPQ8cREqPgOcodyj8vBT3UPKxZJwM/pygAmRGGgAEdJvYR3MOea9M21Kr9kYP
hyuzUWKGLRSeLRx+An+HuWNBYfyHprMZtcRLVp7+9RHKrAoZqdQyS2U9ekGReriPfBs317GQpNNX
5SssjMw51qq9zofjASTmMxOsT6LU3QZIUi1pKOBOYhojSDv9JhZKpJxRGnNbe5xoV/8OhoeMQQoA
cOTHZtbEyscj8Foz932b1sGJ/mX3ni32ou9TVcFLbxTVDZjymJxbzd9xnZnDHvcZf073XXtX7ZFN
9Pce2MNXrNHOpw/PreRM1ttGywvXM+c2YpVhUkwCuXth0wh1lvUKJM0cIKw2MDfK9RhUzQhq4na4
AnwEHbeeCcrqJOs09CiyEi6OGab1qSU5EFljUDs6F/QFTCtCVvxaTrmPdfQFmPrDlp9LGBi/9Pec
LvFzMqEdqPZu6kQvGAe5M+PcCFl/sMxNpeCKNBEkSdupbBW1CK4/PbRxquSGBw0f3JVClhqxekI9
ECt5T96D2lc+j0qetI+Q6GJJAjMAtC5E+v8V/L9LN1YQCl8TjDGvp85yvu3Yeb/MhvSpYuxu5xm+
K6IEDjGXyvP/BFlnjbaBB0ZE2LrnrE2U6IcVfOfwBC+axlKqWteakWec3opsb/dBJMaln/8CEW/M
iEaBJF/EiA+rytsCuFibkfXhiTeHUSzAIhv9QagES3iWPuV8y9NkTWLKXOiOapgbjevM4wlJXza5
Y4r+noXNCu6Fe5BKzLtQWSNbnzWVFKGlL6U/4XdAcygKqWL/bTBhn401V+YcX9l+BWrRS33iju1T
V4VJZuJeh4kyypetAqQpIBl4wxGaM1DjoFx6i7WnRNXP6p8D9f59CEoH8Q0hk16gWVkV8kSt/OO1
3wNs5DxC8pGK03VX5xw7FbbFPGvWaSBa1M57qPlDcfid5zoMz7D6sxYZ/Fnp/s/6UTOQQQzrN60Y
Ozq78uaq+++L1yc/O4CI2ocdDNrlJs+wh7iusht4Wbay76iZijFT28m64JratD9WJG7Y+XhQN7iN
m5nWGAiHS9B5B71Pn3bTX32Q1/ZelBYQD11xoxph3nyMRs0L/wyBUuUEDlyA7TRiA7s5A4abpcmz
ahbB1MpJqIvw+s4kR1PbbX0n0aLbvbgg2qwAyqojA/AX8R/+k3o3n7zeoS322bzY/Lhr1eQD7F3v
XUwSHHX1iorH5UrD9MxqETLTY1vgxYh8X3q7JmeZBDHal+Tr1zxqOoUytJhSKS4EzYah8mPejhoS
fFKl0dDWORs4Qa0kGwQCCmUJl1OvHMaP/fXNttFt3YszGSDdwNrxzTO8BI/wPGsl8BuE6Ruo6v95
CboZpL3VmtYUQFUbEYVbzHTbnnvuLuifsRjwoTACanl5GGoCzL5qJHC39fi22W8y8Somwd18gUji
xglbT4wsweHhQYKZyudf5i1t2imt1FZkAIBxod/TUTtZtRDjaQJDrs7GLfhePpoboJW+wT+80Y1V
qF69h5OqDqyqUy6ER0cAwBJatknXSCHV3+YaYMalkKBiUJKJoGSpZO5RSYUfmDsgu6u8WKM+LF8G
ad3QL1fzbdsDxgUmGdYZVP+MKgkM/SBJ+2HihabumZYQeyLqoxaQpNe+f3owvgq3liSKAZgQvEPt
v9Z5xPuP5APx5XbSz76cjJDkbyU8fDVMg7FUq2JSBgdHwyKoWU/CqEPkO5JJl/Cfn/VKGro1NNnZ
Ned6Ot9x/i0E2W7AUjfK0qnGsasoyeCMP9yzG2f0GIkv/zODqz0kVbzmGwDQ0flWx00rZOQXV6b4
DXiE4DQlCCe6r49yq7+u30WWSVUlRW3FfCKmfqdVF/qqbMn957N0lP6XBlvENAiD+b7PGmdSxb24
X9cYefSF11ciO5MjWEb+pb8WG6zAezKhPk+I/qHBz4borggopTJZQMKtdB6NdTDQkjWf+9LfIw7F
mK5NCh0c3T4nmUPPen6g51f8ZWOKa3+3FmhaSERhD7++AdCdvT6pwy/2xaMJqS1VVv/Xz/De8egn
JN+OkEAH1pcouMbQR+xZRGuF+p1PYQ09NcSWjvziiLwrlSjGvODqH7p9VbDCOm4QJ6c3tDeTcLwj
79hb5Flz/oSNRmQeWEEMC1GRaM57xAutgLOynI5/zz6BmbHWSz++4qjejIu4DwUKO0wwJ2HmEtUk
FIU6S6QprdNSkc/KYSCHiM78DKkfytgeRzYcDMBC0ODqFSG77Haboh9i1dVroSmJ30aP7+58mpcT
CyXV0PFneKuwJa+7MJuxpnHqYSzzpj5NV6b/jGvgAMvM2jipJXJGBM/EdP0uex+d7NlFth7UryiJ
LVTglBtYdFKKVZkdZ6jhEkiSA52ym3jnkUIa8BarAt6SMuGx2BJI3LW6RqX4P96mEx2ICKtREP4X
OW2UDZZTx3Q+TqPx/ROjM6LdAJGbe7WOpRabaikQ/rGU/dIOFEVrozUu1nyZKlukL0swKHlhKCYV
YHUat9ihkNDJ1Qce8BZQ+tMJQJefx8BmKT26Xv1Dp0TULFwDs2j9akOcFQ2ws/bY/PkmSAbez5hh
VbRthXR8Lr8DHtytz0JvKtoHaRHTE/f/8fMmhLHoERKhecgewdO+7VhjPO2LkwzWvFib05fvIf17
XW8M1CbwH94X1iCY+k4hu/1PoremkBwGsjdR9ySLrL3RA2QsD1o1P4RIiY9gWmhSVVMJN90w/zoL
jbbqi0hWYxJD01pbHUPsurFYnKmIEfR3KJ4DwygGa8hUq+1HprtkAm1ZSdEjqMxKaSPXJMZvuBMJ
C5Mfw6gHpN2mg0mx8bs/PQPaYrB4tmk92wuRpHqrUT5ULkftOgaAJZZOgbT91+V6zqCj1IBe8ycO
9IwpzBQkyKdJ5NQ3keBxM+zeXxF0piUgZMnsJoZQZbIBdWC33mQ5S1YORLSPiV9Xx6VVJPTWTTL1
Ea426155Ws2N0trRLYJuJn+nvflPMQ71yKTVj1gkLwZRsLRV4q08MbJu0j0gpL75SADtyQOfBCgy
64ISp/0+TlO8RIV79eVvL4bbz5Lyjpnks3anxJ9k5S7BtQVrBE/ef3oz8wqkCZ8R+a8qNX+FKi7x
IAUNxIfs8b51TeGRLu6/q3XUcDWV4gBz3HbPDDp2nfDHr3bz5tAvBcoe0Pye2n4aARmuQkJZwBwO
PRKhhKdBk3gqIaUocjzmo8FI9zXWKKzv73llQGkEA0hvXz6DEhIq/pXQJwZ2Vve5ulXhYrgw1Z//
L99vi3N4zz7Ky4MjDkhlJPB8nEMJVfiFQT6pM+zzLEmKd6s5S9mn4+JmWIycYtTEZIfZj/jMlG5z
P0zAHDhwdiWPXYfdS7E2FYW+bsjYHEU0XhlfcZo5CozF46R6XDpa/CPdQ2MgGIx5ix2dqpvWcXKx
72DSMkouPS9EDBhjJbWllq3ATVN8zz85BoDFZhjeBpnURJVDT1FG/ooVi8zlwW8+KXVLwRLJe+5J
n15uWD3/fWJ7sXfpfxBozzVPt9cRSueNa7ENMC5no3J1iB+UpNF4gmvUj7EBQPHOYpWOuJqdyXS2
PEK0QdDBnkJBX4fC1BINYSiVWe7Z+4fdh7VpNalJ0cKNy0gH7T/qWtCDENWsdce+0Fm60LqOxWol
dt4mYpoWGEfVQqHelu/fQ9vd5HyfsUPAiZDpwgLJT5777daFcnjfh1IooIXJc+N+c8XSRlapZ7GE
/zIhW4mWfCW6LMfDAeX4gEK19EYIF2KsrSf8BC+G3dwYtzcyvBg8pnF69PoR7TfSzzyAE8f5yffz
aOjf5NZSh9oEB48ianI1yrFWPveZ0KQKVcMHAXnA7MQK8ENfv5WVs+tBqS4cPErpenDBnK67xdxX
rBqVPG5L7rQpF1vqZuiKu0Mv1GgsvLbeyG7maF81TlAGUcx0Ul7ndHhNedhACkcxHd04BKjqps8s
2fu6Qr6x5IVZI+n+BOTS7CbJtG6/exaBg1vMwiEE6R0jqJr4T9m5XoDnysWX4oEC3TWDqq2bvKMe
eyVDG6gxPfNPWu1tsBYUBpoeyoJdYs6lIMDCsst9qNRO8gRJknWL0WBWAIkW7bmrS4N9ZdrR3CDc
fgHtwpmcZAU2dv8lv0tHvmNQeG+5eEZmVveMBrwIbD2dx6k3ehNlX/gxIddCdj59v+n/jsuFRbAk
MakuXc7yZ56c950REGnW1U69UMWlBAuRXMoQQnlrRgxphm8R+qBlXag5O5gKMo4HgyCmsfJxF7N9
jfQeF7GnDfuElGErh2XDFhNziWdvqxaGLJZgWb59tI26W+SNCI4SUwc6aEfzVqogToQYE595vbyr
InVyLdu0+J3MA8gZrTKpgDAI+w9NEwIdf7TJ7C88F1ke8gEw2iPFD62O1e4aYpmV08GNQG/RCpCv
u6yP0idWPeIgzAooXYZsTsJP4nvJsua2o9pJOpfZ/z0oRiynJvaS+VORkeDRV16/MAruu6zV4zuG
SNT2AyU2pGm9vRX3SWIzHETxApLFwEEztNthYyXv0Z1M9jBSQVOfbxi/NRKCzoqm50IJBhzCxeGN
0ow048d8ivza6yCs9uzWX4ZmDVdpHHi/5ptK3sEXH77VlwNoJwoYmGeNvJig1rj8TfV6KOPYdUbn
DQ4obyAPTmWJrbH7hKVx2TpHMOdtM7a9vSmjtRw7FzHQ/A05PInmf5ISwPFgObLfMm9V1oEpNRyw
CkGKLNDkvXSAhZ3RpS99Nth/h5s/5W/pSKvrgZSiF08QdMfJVtRIo7VBI7vXPMi/Kjx7SgBwljtX
KggCQF77EsIeSCdFNXyNjvt/uJwFvUEGp3zsxD4z5ZbjlPdK1g5RVi8ViiuwYdoX62HggFCiJffm
EzVBAMVo+PHlROjLwTQ6eMIfJjC7GQVx1hcMCRRO+Rmt9rgRIxwgZD7cIYAIqiaKD6X/GmQGM/MZ
MzSueJbNPJ9ThLW6YslAr/sXUvsn3O2EjKJx5QzIEM3wTSQIlr8cQ4SvSBhEAbZWzcuEMVPKc2kI
b7BEOnOKmwv9WrlFUOTIoVviB2glDxFaqOuP119VU4piOd04V2g6qvh1fNfJ9zEHe58LXC+qy9dr
X0f0GlVRR6Jnjk4bkbOmH6mtngO52/0qR3QitH8ncNFMx9uIp7gcaz/xZnWRrqeyCfj2vrrQEdll
tfEHdwsCHAfqKfpxqiwYLkhGnbU0ESjKVB9AT8wq6YFTh+Q8D357Ht2I0AlhMZ/2z9uCcT8mP7SM
GNYija9Nj6Eb/GChNEf875Dd8Isa40q8qUBGqXx5bgL0KYBZOjc/ecZnCCv/LJ5e/DNuhqclKsMx
f3/tCBRv4CKMRF0CBbYDAUHreaTO7v70oQ93QXzONG3qJQ14KQL32TvF1pJyZ3uUKNTx5ynR47MD
0qv0oSuUbxADPzawe133yiMF3PF/O1TrCyzEL9UhAL6ZI6EfrSRjEES55AApt/FjIH15gXLUy61m
b1KRB0RtOPdUqHvzWl2ehcjajdNI3/WLHOT6wZ6+vUXov6giSKq+w++jaYOo2+TPLb6y9t2/H6ox
00ti/N1rxaqunImt5obRtQgFZo8tn2hTyO30yHJfLOMgMR8s8Klbv5yBPWAzNS/SPHJGu3/1AJ+i
4qX05+A37WRVFtLRtbe6ApGB98l+mqfXlBaohWVDi4/QDjLv2xRfamrRtB89+i5LCOgCgdF07G3A
Pg+LV/nTMjvueud3yrhQPcDhNyEgasMBKo84Z6IRbIstKtfrQ7gR+ajFjy5ar5ijs99ARo4yg1KL
NlR3YyI+zTr1QJ8Mhu0m6vic0MDqe1SEKF1XPQqvX9pw4Wa6aoq+PDv8TMnWuZSMPtOc0ndP4Rid
A1hy4FRK/U5UuQ4Gf/ZYeoRZaGVqY4uZQgt7PVU/dHD/fozPPiPfDcMKqOBmQahuDUS4ER5rLIgq
zQ7chtqL998a9wJp4N2uSgrfEqYibFnntW9VBA++k3NwxaH+szrEe8W4E7iruJhNnyBVaXrQAoXp
xaDfOMuzULIt78ZvMHch0tHQBZ4Igssw2XNrkbvfcXuYL8bQvp7EGh2fI8BRDpz3Nje0LlgIt5iK
Va5GSRfhRK8cbV2lbL55wDdAZk8p3ua3CD6j2vppPU9TTv90LeZZqtvlZ4U4vEc9cisukwC9YysN
4DCWeTVKa9A3A2NWhNOu3bYxdASQJc9oV3g+blJb3IbPD79qRdaYLEmxHStlSwKlrCyepF5FMS+B
utwsJMMBip8JUmOFTfJ3Dl3RCQjf/C4KZVObHZwoKYYlKz8KuYXCMbBE2tKrOEyDJ10s2aULL2p/
ImNHpGiuCu59FrfIZsI8fwPLlwY3Pa6cx99mKPxXgKtdSnSWp0kRMsnybeYjMgsOqJtwjmCB7dct
U8sn0tnI48XqzoHE9idLWRm4Ci7wNgrfpMHtR2gNIobKub966UBemOttkFb2ZXMUhiMeWpNMbilB
oEXaFMZi643EKKxesIAUIVGm+eWnwjOs9IuVwlWAz/JIO5ilbDf52KtLuJoFITqD8w46aSPkbd9O
11frVD++CF73c8q0QybO4desD7Y7/dcruztZCdQA+IJzmxYZND0/9ReDZE/4lZVKamMbb8t1gKI7
RNKvw09DgwGaEJX+PYa7apO9CGQXSF9wVRLMcMNYyUdqfgcsZv7vZwJ9uG/TpEPDlTJ+Wf1/4p3b
fdLk8vDc/IF5NnaBObVJ4xqywGwS2Q4fcF0S232dRnGVdxhQ08J1HYoYJ+7hkHXBDvyOUklCjbdk
WwxAqCW6vlw8NM9iCi9zFebyT7Jki8Vtuwx5f8OlTRPPnD+ymPK4q9/P3wT3Ta3sb9DZsTJaYd3c
B77FaNfmpscA+agZJj2LKqPWWr4BUa3KPVPvbD2iianXdAEaeoy/93uG1MRs3ORkSrUSTFUmfqXd
URhKgiS1kaaRcLRY95cYDzZGUnRbl4STucABFl5FITwp7DeB6qBEGaLcDVYlib5BD+xscCZZkI8t
cEMfBVp24zcbZn4gpZyVAPBS/Jz++4SRxMqAQ8ADbnHjX/Y1GJBMtzqOEEeImXSYfijYlQsAxjDT
kpFhr1LIFQVAExh/umgEO7hVA7sKMI4ocqPo++TO0b6EtMiPqWtxw8A27i0vZuPsiqqd6dbdK7QA
jKcOSgmVM6JeHJFODQ6GPn+eaDKMW3283AdOq3lUxwyFFOZG8Ccj+CACrMi/Ka6uh5IyPPI5RsCA
aZcr48CRofNoJQtA7AH9x24wHyN6Mn6s68pcCdqPocaOyCXNr9jTYcuYaSvyXkpIPco50JM4Vko4
99cWG82qE0W5QRUSBXBbBQscplSh7NbmIoPhPr1eHA8hYwtAtwRHY8ap1g4ebLH62m3wYBOeN6xt
KaTSce+MWHmyFpzONwQeS1QsfB1BxqqZKvIFo9y6UTb9K0Vyks5Hqe6ReNsDS6GWRfMG/ClBlnGa
E/1xoytlVCnknUqnHGMftZJtZo5FkKPIQXacVhXO+dPMz2B1hB3RUS+OpYubsVAh9msoaSjZ0MAr
9SM6gqXCgqNMdFRbn0JjK6W6hGEtk8cuPBU0fKh0G67+quCj+kL5zOlfHszfOoAG8bCSZkKeJcna
y6qtSm1lvJdnq5DPnBL6D0vN8knEoA+ZypCIBwqjG/iZpNNW7EQR8f1olVCAddOkK3YDOJLADhrl
djaRQh/FkAmiI+8dbgf6/9p6Oiqbbhuy/mLNxmpvnRElNVVgwH5UBc3CDDZHsjbVzuNpCX1H0NIs
yk3r3ZL0n4mE0bQz+N8V9sF89XProrJn9J2U8gSU2j/kDL5tIM4WPyP9Qt3q7RyiXqr1f1ku1iBy
5U8oh33bf0nd4sWGoF9CVn+4sxu9ClwTc8wv7CQkHfS50XIuFQs7KjPYnmiYyUiScPvyeDBFIj5p
wtTzCkRauaiGraeUyQYFBYk30U0+0VOgnae87WdxksyWTeXdI/VbuWqg7vBPjv+hjWmhqmN0AvFw
hLo13vE4wgyW1zXX6dVAIGycvcsqnxOtlfzHYe/yo2WLEYULv6RItfh2wavFQJXaV+56+douVyRp
7kzGiwNSyIzUFBHGU50MoL7O79i28WPQ0mwo/KdWv3gJRgEda8TY512hOHj7xoQUOx01MmX/xChB
02LveaF7naqIVeNHpruNMi/zxjqgtGP+DimfT5mqlgaeVncNHfnqGXECU9gMZ9eFckrFPF22ECa/
r5WsQtS+s60kJzV/+SwI9FGbieLDVPi6SVj0Z199vCHlzhOSlypykE/Eef4AHouEHLODkFx2D0sJ
kuPxLjiZFnDNOdUDdz018oD37qF8J8pYbk0ZWn9okhcnZZQN+oX2Tkb8u8X7Ur7hvWzRGhZiJPNi
ZFFO3L3vXfQsQTRTUSgi+yPcyaIJ8e1iKHEkJbFdgqpvVCEYep/qxWJwOjANhTKqhB/b/QGuGdmx
WCmlDCEsBOo/8xWcf/zKBsPBRnHTC7Hn2yrHUQC8aCqCQ8g51SMiq0JAPPkkF6rNqxQcL1bA3Rq2
uRIxmFUvoFA4yql9fCN6nwOEy1uxToOgx139RoM05b9SkBsMu/a2I0UWXGWPEonNWBQkDLbxjZD+
YyX0gK+eRYMJPpyb8wiFqofk27ExghV3CrQyQZ17UBv59sd/1dMZqWPfz3UO+Q766lcX11XIdMSM
LUAYnd4GBgc+OW6AMwAo9hKVAHMinyDqnMw2LTcntIYe1qaKg372GoL3n0BlMo54UgARxQkIM229
YGqp0AM9S1bNKHTL7WjFSH7dgqIk2MWXzIBzlLAqjQwLL1VUR7KwyNIsTrI6YS6ZWo5KctnpVzYv
IUn6nECfOrDNjHwN17OojWbHgDQk+PkweEY4bjY5S5rRFvDkFCacvl1gyfoWjzzvqLUvGkheR9RN
BaMY1neZbw0lQZKh+424Br+i7FTVOt8TqfbXWLBhTueuX2H3TmCJXphIu4AFiAOpTN/Vg+UyrEMz
htCjjfoo+Csziv5weskBHSoZtvTJRQMm2tK4Ue6ecIIgHLkw7FZsfHkBtjhphIa9a22n/vej3jjb
YclVbHX6ZXifTXP9qh9ButzCfG2YPVhvwfO+Kc0vmIbRe+uEUMN+nYnwqsqEk+Za14WI+B2d0MYJ
omFw6PEaeZyRKbOrM1F1MnTTurcDQDffCzoXhGu/u327nH3PS11jL7VzZZRjXluExK/gVfXSIOfP
E1aZPHxXmTMjATGYGXg8y5h47Dd1zKYZMwFiIlQrLK37SMbVqQQn31AQzAHWOv65TKCBsMz8J37F
FLmmXlgsvhxoC9+/WFVTT4yHPag8FT0jaraJkB3nm8IczZgkxBG9OwGo2wdCHdYtmLJQmaqvUTue
/Tpuah4TR27z95CahIMFAy93JnZQZGm8v0+1/zIb8U5kzAFhwnngWRnXCeBWlvatpAEcy73vtagX
Fh0K2BSKMntcw50LoiTE8GlvovTHvV6IQ1xMeMhtJUT7CvkdfQh2QIrsf9FftH/N3pxat9Hu5goc
exHKi2eLIoj3oTgDKDnjOW+DafNLWT0PfckbvIPCx3fNYmHr0qzmRl8fNC1cfyeELqUvglSYvTnb
ytyGZixJ0ebXi16EZ5J27GaKQAj4/Mm9hvejx1YdpK3BXife+PFNV+IISRowS77cJbOeli7Pf410
FPQi9Gib/4w2QBLAro0JkGVgemXHLOcl0wE9eDLNZbXLd3lLz4VlwnelYeIyQl8zE6CSjWs+x94n
TQo6a4Nta0SiXBTsBaZ2TL/HTkEGWE/xzfcj0ExA9G25DJxFbGJyz6aNoEvfUeisIulRUH2IhUDs
tgyOAvudISQ+Yksq5ntCzKVb/idNrXSwuctdhOF2he+S3+exumTESuAipz4PwkoylcOr/VE5Qpl3
vcV/CHnfClwRXwBw344ihhy6+01wtXy9WvaK6a4JC9ByDLUZRYkaTzeEt7WLeuWR4n2FW33tjFU+
0L50p//mdBQxpWVsc1hSSL7IGdeFRHhZ1nznCQljelpbznyL8eBqXecPtsJwI4a2daEr2jEHQjjg
OPMpK3jpFzwY5FQKrBq8MzQbligDvWEgK+sObVLM7UZJAhsVpOPQj5Ug20sY30HI3sj8FdcYjbgZ
vKyQGr9LLUjqbYcrzBVh2mQhbxVq6UC3a9q082u8Qiw/GQcd5rhOjkblNJFkS7Vg7SrDPHez6HwX
vDyRwnEn7x6AmKgAK3UrSwVnYR5RjkyHuHUt9I4ELNNh2yyMqMY03ow6I9tmyfsB26h4NHyUxYh9
PfzroTB2XPGCwvCVfjA7558NdoTGT9+by/J2dT3K0oZDSm21ESRiqg+ToPqSSbgoz5HMtaKtPMs0
IaAoMw/+5z6O96xaNDqdx2xDTbgOzIHloJX7ZGIIIVyJE4masT+qkufOQ+fsVe6IZJVuFXrhmsi5
gb0gVBZOpxBtcgCkWZiuSphX3fXzZeODQfMH3M4zpyj8Q2oP8THWG6J87bfI+b8S64d+rC7RSuVH
i+0rDN1MVJFfbDHr870tcqkdBjDSV3ve+e3yj+7rUWhOS9HRNDj+MBm4Fm9pVxMZDoBXlpZr9ODn
dtHEnp3jxSKrdsKMBH7UTuSwOW9SkZGiA6O+lcr6TXZ6/7eL88Uerpye//OR9XYYiLcVzT+fDLWv
p0OIRH9SI6ETw8XA+qwfXhV8D9uQaUFbKhB3ZfFjsqqXguho+6sz6YfPGMrCg2G9jPJPb88fbL8i
+gTPDkhi8NCdFcB+mHmPGO/QOnWNmTRmjEko06hbo0j/G7OuPKKm/34U+knEYd/pUtao7TNGaz36
CAzmc52cX0aApTKZRoQ8XtavncyR1IgV6Kqc2OHTLPZLe0oawwhG6WQeFJUCZ9+zgg2X/IwzXM2X
0oy4ofOLlyzBrK2dDKc2DiPpaUmKUjy1Sjfe91DxURcJQkmCCdyzFPKE99bphftNKRLdxNmM9JPh
Et889TsUaKIRgY3Nt+vz9+L9WAtmdI30oZR6oNdTHDuR83jhwHQn4hYKzca5J0Xh8ZYVasLi+6WD
7ptkNGywn82TYPZWn0hfANyACZC0YY5hnMMV4mChWOQWtk/a8ICNOH6XY4pHoZz0v1yTe89SlNAI
+mnhpfdgTJBOw8V2lkWOkpDSTqY32yAHXrlLlSR7fs0bbUuohr/wl+mQ11tVTLNJ+wmpufhF1vv2
6AFV7v7TBzVrrkMT3TAJLicI8gnfvaffrgD0qnciXkutTIuxc9+UjsDIuPeKEO3MgrYDDJ5j+H4i
VlI7Vru63fnVqReUh0CnyNwLS/sGsBJB6bIE1wgSHw5a4e5s5oO3skG1qBiO+rVpavVpbbEEV7CK
NYp6g7bHoNrH0IXxr/WYbjFSXRQi6By2DXE1noTLuUP7RyDTlKIUIcg/4IbOLtW4F+U/X5gnKveM
Cw5L+KOCj5jEO2W8P8r/bfrb7WAR4usFkry1qxjR9L9aU3WpYu2lBJBdIKdwxxT+TVy4EnCGrpDG
LvTLY30AV+cLYOFcTy4e7HRcTko5zCbIkkOkuhypAagunAKBGrw5VPnunrpE4PugTG5U+cZ6T5YD
SSn86RBUdpOeFQ+vVM/mbpneXW9P+BJRMhpju7aLo0kOHYZCkvQHh2D02Nf6w3PnyucOiB59SMOc
+s46uAMiSvg6F+WIglK1MQKBzp+vLRJl4JW6QcG7o4w/O++NmcJs6S7CI3x+XYlod5wbrqeusfHh
rLOG6Tw5HBtWwmSw7G/VQnWhqpFMDvxHz4CrJhTdw2JLfZyJ9U7XJcneqYl3CmkOe7bE1h3T+CCi
URnasAmoJzs5M0MQWPD5NcpPHiBeInirUripw9VT6zwEdJm56FShZfzfVazaTxVKmiK9B+vBMnVa
HU49X/BxRFmOpToEnhVz3qTmnBGPJr0ISGP1UVU8LFPB9JEwxY1yf4E1GPWfGFVSwsTxmCTaLtow
PGyYKngUMcykaD35lFIy7uQRwzF0BltX2S/KbxKgmYo67158GMTZqtlEebCVjxAgONxSi/tA2UnB
j0AOiRCj9DCOd1FainL7WKcTIdY70PljzbEyprwdMmj3ygRf1SwsnTefj6USZbTp9glcG3jk4bqu
G/ymokckAEzSdnis1Fl85HphcRWM+STmoFr7IawmZn5w2yUgSb2kgYh0+N7tBrt6e8lKwwNqrzw7
UOD/TV36kuH69GSmP86RsAYoD8aAHkKgohrdgMlmrmWdQBjHNM0CfRwGmgxNAYv82osw++JO9veF
0IJWUadePVLDAYLheNwcDZJv0i1va2oiOmwIUp9Z80hoo9AWyB3uk/CNZetdgMkuxHhaMqMQkydN
CI+XK0a+eaPwqCSC5V+urcuwL01Mzz41+keoupOPynvkMN0tZLItJ37aCOX/zCh4zSgOM+KMWRR+
r7A6KCJOCFbGvZ3SQiLoUdcwlDPZT/JEqfnEi79d8gscLa6bTlmxYQ2aX04PL7UIhErp75QbQnxJ
aGSnpsZT8fkS8YX3CJtWkCIoy7phOBU+IK6gt5602stTCXT579TEZyV30KRPe091U4hBlPKHQk3O
0j8OI4//Wm2aBmgtQoKo+eU+wBPnzgBFduV9hXnuqbuPPvaVVa0D7NJZ3OkFkRqBIL8iHZy6RlqY
7ZYdrU/REjirHALGPxm9yNhjOilId9NJbjnuggwRVBCcFr2aHREZog2rwdRSOHWT7+O1nNG4h5hg
qlGA2GPmmgvF6RjJm4SPnjCDKdFqtSdRSmzT3i65CseS02e7NbIUWI0WlPOxi2ITzvp2Hg79l52h
ng5CXAHr0gF9huHpDMd87jY0TEK83sA16eesCMJp4DNEEapvcvs0HB7vgkhYigC1bgpYevQcymxF
rr6oH8xh7g4NnTV7ZUk07o7yJoqkM0lXCI0bcl86KZzCfSwqk5yxd5g4ngedxbJZOFNPeEAgQ9CZ
Budd7SLUdAKHBeyXsCRnFUOb1ohnMDtK9g0Z5CMNSNcCPGGuZvJz6669BlvX4HyCpSy8j73lhV7W
/vvzuE9LzBFN97qNjGQ9Ndn+H+OzA9/9FuJXWRPi9uUmFKEO1Uoql1tAX3Hl7wsm4AzMb6ThnGnh
6pE9OeoMMnkEcJFM6i4S1EyVLvt2bmabkofOBrXijpTtLiVwOn+s+OElawLdC8IuJHBREkrw3EHM
U0+dYD1P0X5VK1Fo+gYEKzAdNddXcVOn2q0lm1IppBsfTAU38wqREre3MCQIA1PqF14shYxow8eI
YmVlWh2imtO1FWAjGSUqj1JzKbSt/rV3kLEOy+WwXhyXsxjyBJOyzWGkUKXuaGxGSgu4HDYegaR5
nCSh90toHUGLwjEttEg6YJBLQOMaZc0khZroexHb9kvruFgM1gFG0YHsucWYD5udppxIrRRE2ft9
X0ZVgyt4YTVpgLKWobq14+yvnBEQqjkFBZcOjOzp/MoUX6D6vlZVYIxPKigiIcQ3lAAqZG+Or1zy
DX8iSn1dI14JqOYMXmyuEz//gwFnmY04KfkwVFtJe9FKPxemgpzdpxkQstgztVpJjJ176vtJYOpe
FEV+D8zKkwCi1rW71+1UTee7V50u8EX2jPYmZEbrtdC9MZE6UFXhI5XmVRK4O7RjAaRLiDRbD9rA
8FZcQHZekv7WMOvEInzNg255aw8CNnnoDQmRNaVGknOo2NG3DgDKL6XGxyouuazcUfyC6lYTK3Zn
+7lnaHDWsguhJ7N50ilC0ed0HTvYy5GqCKZz7vzIvDi36sQ4eQpGUUmqWeHp21Nr3Aq23mo/ttti
FRzIWeavQUj+Vksku1kw2ud7n4HQBpwTBY++QIrl3WJ76uwsrlhXGyiGTRNBi9YX1hWAwR0hq+TQ
7qi0o55DVq8HyeUapQLp0YPNJpVMdoHQi1Bz3zBGn1CsbCgOGHy+uDTq9r1ciwqyMLjlEP2zmhOa
7hribpi7z05k/0BAECWPY+z/LixtczPpzAnmPgVC9qSoPDsr4SoYDJKWhQaclDp3dh0IJLzJZj19
lVkQeSi6U7WT51X31WKJvyEb1DXMAIyqxB2nl3WLvK3CC1M3kEomxB6iGwM1PTz0OuFUqsUZ0wxY
r0N1S6q7exqdB8Btw1LHZtsMcdFaIVqrb8rK4Pp2oxcr51vKwDbb3p5vKmDCHxeZyTYXi3O7d0N6
bkg2pUXDsTCR7RQK6sLo69gFVpO+w7PxIEzzJCsXBgK6WYMPuOrxAqY8/KGl6x0+HRG6NTjPO8Kt
B4KNLTm0+0zn7wKWqMyqPnI65KL+70gRU6CMp0xWcDiLFGpxI4aPQLHy+EBGW4scU5mAlIU9Py+c
BTXPQzfrboRNBJZQVqa6MtcRiznMDQT8erylFxmsubwT+WnTV1as7/o6ir1z+Y9HW/EalnRO+LlO
wDqeigYTrcenThLrArb5RpQRAKbrzuEZzaRX20PeAP8XSwqxzkvHoWL+ZtMvIH+12Wdo8L0ctREA
o5NGQaca6L9fpGP5XtZMpvR79kQJGDdO0zZCS2QxkfkOvEUpPbK2yMKGulfMqvhVVf374qFE/mVu
ftFaSYbaMESTCTNfeAxaNA+ao6h4iWLnnnPkJTAAl88gtrfa4DJZW1wEgwVRniNSQABSrKE8s1Ks
GZj5rvz56vMqPMEQPbMLKP6ZNRpwf0SGo4fk11d957qWxYz0DAqGNTNJ/oRjFRniCt4MZMQ95dz+
KCNy2YEVzMUZfRH6JJSbAmUWmOnpSFC2f5Q1MhP1Hc07q9L1UE3KU7x8PAUIukEZn+hdpCVJ7nZ0
Lsr7hwKvUklAhRO0k9eY+DJ8RX1fqyqIiOzBCPpMLNJXbh+sOioeCgHbTb67CdB/LOkp80UuOsLX
KOibes61GtcqjSwiD/1NM4eU2016ObJdZTMHEisNyeFJqGo4wcHUytyB58CbAE8Y4megUP21KbFp
J19MxS52xUMEl797eFHK61Fky7qh+9+KOocDWIgcI8WmwAu8fpdgvCVFaTGtqULOvG2MOaensC2D
kkz0CPi2/6tcBLFPiNsPv25h3edYPyZQ/P2HU0SKnGTDehmkOwoTzKWDPE0PiG28Se0WvFd70jE8
p6Vy6iwjYJhnu3cMhX21f0nGcgozmQviXXwx9eLQ8D9XEW0t1U/cAgGq6hHYpbyne11t0O/OmhWl
N4ugTZEjZIa3ChSN+1YPSgI+I6AFFHE/pzvOq298NKDOjlW4n/BzbFYRgflPNsgrsRmeZu+GedDi
L7rw6FdWd4rxO3F5CQ9Sp83TR2CvB89Ld2iGDel+S3Mo2p1pKVflJb4Ms78bCqt5wOZAoE7/JELn
qLVVrVUfw/kMYyOfyh9UKuxMR2s+kMYpQqKQOszimPD+QBWPjbTbxwPYDEUbP/LsMSrAVwBe9ZR6
sNvxrtcwBl9JoJw4qHRkxhzo3mvDnM8CtohLqDTb58gQnGcI8mRw3v1pJ2XTqkCL1ePnjG72mFbE
zQThrPt+0b/MwEjwrDkCabTM7NqnEfN2tYRzsFs/B3hr8or56l691eDMex8Np7o9LWK0wikOABCA
pCXAA0VfsCBzUbF1Oy5VoD1jr/h+IE/MgPZ61qh4HoGr0lyPaqVFMVElSqJADISpb/buADFi2OtD
7cRBkkvDXVk4ONJK8uooRu87jmjeMb4ooeOMmr+YyPwFY+xP3UvuinpXBPmwWjkZpPcy7mZMsTOk
f23CbVmDcJ2/oZyrZicnapVgMtcXfkk9K1SfGFpruU800m3V4jeFVAqVjFw6NZjUU3thh36WWsLt
r5Du13j0lhqDOeAj28w60kWwnqRV9mi4O5TPeV/jlnCTFnkqKeJIEG4KyIU1XY3GdGgP1E+XaqRq
1Q6v0KBNTauTz06vrQd/PCBR0AU5JKIZP4IYtn9cxaL11d59JcZbuZJZEU5wyq9MoN7Zhtr//cyX
OviUnyFVK5MQlif0vVIcKDkjgMkGm7WJsuuaqxDJaH6lyo3WxG8SjC4DVebQR6o02r3iX/CEXrUv
NzVckVeumSjMTy5AQNf4EpSlXNzIfnA97QGR9FTbpMwa6C9+GNyKW7bTFkLJpSEFTDtY+qytyJpb
WoIDKXdF3H+YJv/QtG2j7bFeTVjuErtdPSYofqJo7JBC3pJSL0zSmwDnIs3uuUvg0bou5LSb4437
ZWKMSBsKrQ7ffANCCFhGndVT0I9auFIKUmYTYn/FQXC4HCzNr099iNVlw0Nwz/n0G4cEeLjEr6ez
4DmgdVq21FDtxFl03Wn+j5FfbgeOP5nh0llLlEnviztUK1Moh0GtIdwHmr5TrkXPZRoZgecdV63x
O1SSYjqo24cexJ0xK9BjZvGK2KfpeA2yYxEvs6CVVkcTZwx6h+Y5Bj0e6A711VTLyUsqW3vcHrzR
W2y4tX7kXrg35QXQ2TOcyOTYC/3cNImqy6vPXA5yWHVYM+r1hxf7m9JtkpPfCFDK0PCcIC0JDRBc
0TWL0rhifLSIdNbexPV9Etfb9zTZ7LNLdlndEN3edZeeopBU7jpTYX1ZARah6nQyhuNpLCwk3fB1
n8e7Vfsjsb40UnHSwN3hlyicJWJOH2cFfAvyVjK07RQJ7tczY8j9s0+9n41xXnhrSMwTnEgs5rZc
cO4M+hZPFL2evyQtgY3TSKPxt5f39I6Rt+U6f3pJeRtk7A4RC8zgkH5NBh3ejbC4jG2YYkXrCcH8
aAVUsGbTNg8/O4KZfNT+6wmL7IPa0ecIpaPB0Av36VvsSS47wyRh/a6vhEoZCVcDuqUO0igBVJJr
hVDxPMDniKwbLqoCseyX/I+6+nUr6wYACCl1cm6s0phqKELmLT/IOEU6C2uVRUxhGC4K2Er9zKKA
zUIyQcINHZh15nSdkIZj8e6dCV+p4UgIsF8CHQegiht2ob1CFTH3iljNBAReJM+cPqA9EZsU4QbU
IxO2u4NRvC7seZDgarlRxEoVwcNCxjNePN13rrVANILAK+Jam6CZ3OOiPg7mAfdUAlOelefspnZ+
7/Q0vEHTMTg2EIw1Nsb7vs+rv1jBTp8RXPFd1OsEU75xu7DdwgFCKOPlwfIBCT/l6lfzo+I91g99
mi2z2UQQnPGegSa4P9muTcOLNMraDVRzxxSzF3hdqfbAo4a+VRBE+xPegxrpA9MJ463fn3PGQ2S0
tTwrObPOSReNVHz0bse1nCKbemO4JC8z8ZCmYbR2kYciKgtpv41I/UpuOFEIKoOdATOoQnkMh+j3
lf3ORjMUSYc8KZrp+LOGlBPVWDAh2B7CVZXlBwK9KM4An89Ax0wmVMaRdr/S3I0h7aEwLWAwIoB9
td4q0l4Di95SxkMAkjuBZQDGnorfrBVfSfE4+mp1sVId7MlQDkHlpjcNRHj/jZhRvH4F+nSz7wC6
75VLobgBxv2j8e1Ac+6y9anqEpsSWPqYMiUZ18xZvGyTijY0KsKJScwWryHhmbAfpzOCH5BsHugI
rRW1Rlw1pgdu+hKt3bDqBV++/sonfeM4/9Qh0CcMIjTR3vKrXRlurDtOxYSdfSbaP3KqKv32PJeD
/PG5tavDG++3+NrPr7hVTQ7UlD2qxnOtEYySl5/uDBztxZR9CSDhdHsvqkTzDqBfTIjRPKtW9CjB
udRpL6wW5A0TE+uwvGAdftR1+hGNuD3vx26IrGWf9hFZ8Za+FUvwUN/J2KKh0VbHmCBNH4JZBL16
6lOddBkTvUU//dKxSH6ag/d4vPgxTLDBtIRfWcvoGiDr6eIXp0uUooThToxLjcZivi+k13T1H7cc
VHs6dvVmz1+ZkGDm3V26NUDRsmfz6019I0AggTMwGq/9u9hp95TaaoVbQ773kmvT9KTIB98wzzif
toS9mb6da1zJwBGmcvUr134zj+HEiuHwAlUqGKQ2m8+i9hNvs1SYJsYd4shJKIYkFAXBMsPow7QV
0yjAmPJfF1XDTJOi2vHdCEOrEz4IGJ0B2I/gw02yULPXX2eXJFnQlX4cd0ulw1wG/JLsVriHmNyr
Efot3owTHOkX8vE3+q0DRo4OTJAa3d32WruqpikA+1ATDIAdjJkXrPPZrfEw5/LQzW7Z0bnWsFM2
MM8g+Wf43n3UEDZzM9mO+/pLsm7z8hYuE0TbFbCN77yXV1ExUqM0JRqgzS7oBf/5U4XEEWk91wKU
8OTuKm+u+ltsyU1aRAf9eB+4qwxsbLyArH32vcgWBzU8QBd5CScT4xRHNRoF9Zy31S2q8ehWQEFf
ZWiHJoupjeHoC5g+xXjdm9wzXFJ2IcJffxo62hliE5nxadZpr3+vMHC+yGKid/N7kwfrR0zEUR/Y
sUw7rNeEQNAEr/3kwGjlmDx15o6VqFwq5Tp6HkQi4vclQiawUN3yyhf5PypIOYBGHTS1LBBInAP/
qEOSIYvlxnN7bD0wDR0o78LLNPUJgiSSWKL5VnZQtPDn+CAEfN/SO9Ifq5L6Osb8RdIwBJqXTvyP
/4n6+40Gnt3Li2CnjaQFGO0LdYxl8T+oCwpPjxLJ/eNraQ+avW1s1/gQXz3rpVIc1C9sdu2QaGON
/YUZP6sakQmzNQfD0iD23lqWINrzd5sXAKbmPRwtK8INpSLqccerGRpKv+jlhFqtNtqPEwp3BliI
ytnYcoVxtbCXZC5nwt0Q1dRGVVI/S4bXOGkt5Q25jlxJhGW7ebDnxIHX7oVtL0zl0+Pt79PMsvj/
p3RtkTtM0BB/h4l55tCY5ZiezrOcEB+s3xLphr1Fov8unajQiJAqisTIY5BFoPzdj9NqXdYxR75I
bY4Rq8CkwkPGW0mQ4lR6AdklR53Qc7F9lFif6X1n3c7UwoW2dtolOdOXGL0dNDII9/mGjaCnFFYi
a/mbbJE8K7nfbQUBW2j05AvJcp3GZX4smN1AOnTBEylYnHhCV498dxk4KvZiz1nqvJMpRaHlSU2A
zGdPxs933nn4wNteqMO0VG/eG7s5mye5GcVT0ceq7uTCX0Un1E9BDEwo8ww5hYytFe4Ar3EhtQfD
5VZWbMsc4qiX8EOW7U3NWIYdvgw/qekVck93+TKM+97YEdbMA7CXqfd2/oMaiqubW4EZGAjucs75
hgvpNwwrttBnPS6uWGco1af/kZxEwCYHto9u1cMnnW7GLmT1H3qyY32FOM3QNNT43PgfsbBXWGgG
2JdMxkbrEbSGd0GaOCYJGPLJK++fWPsbZA1j9WoM62Q0MwcH+GCSNBNmUSQw0h8nu3q27zMwNpxk
ygJc2/7gwo1Cgs7x7eBdJ4CJ1uVTxgGiRmoAfR1kqCo+W09rqpQLdBFa+ACtT+iNBKyafN0MQEKT
oxE8bPDAitMh02HGMgTgoxmwpKszKozsDsvv680HCwSsQpwZhDHMGTF3qkodBOzEH9F14kVkcYvW
hISn/7ZslwbUmlfHBmq/dPY2psAKyyvyIKIphz4XKRcEIAtRFEjPyb+ib9VVDpJSqhaqX/zhgb++
iSOJk3UKzMGuW7ShoStwZThnLjCwwPpeDHUY2tOh4WrPXtFKADBC5Ck+a6ASVgXowyICbiT0hquk
c/C0ZqV3sN6TeFqBrLDDP8ObabeZoHQAur1HNG30sQSQUf6E02YqtmmIuOPZH1aVkhj+eZt/jUXn
AzP9RnzkXW4pfgq9TtEOAKRXerPDC2luspGcxwzHuqC1Ok2gcLA+P4P/hfchsYpKd+rm1Adj6EC0
F6w+eqrZPbSZ3XgmHebOou/NN547YAuyLZ2z0VID78Db+War/MrZSgmTbeGRXJoNY2Pe+WBiKniT
e+C2Fph0C3IOLjsyzXsiX4CBhbHtTNebDHsGy24ODZ6/c9TuxcA4tt0/ZDZpocgOWYdZ1gkV89dk
zwKEGxxtGUPRheU6fcY84X+iV2wKKUEsP7yJ+mYAUP86suuB3ZArRG2WCduJfTyrhtFnKTzewdRk
xQF4DSrHJuO5BEGWRPr+YhC8j/K9m+vvdVAN846owdEZV85jeBFRlnGPoB7lk8FxyTXuW6hOlV8h
xGU4GQ4gMZCIcA2Pef9CnZTztJT2Ptbi1rc5dbts/Rsaf9nzu8ITbhetf8Kv5lgBeDkwfnofxfiy
kYlfCIRCEHThst4Q/+gRQVc6JqtjeNfLAMXEuOrPTShHTPHuh/MHcylfoSBi/n3HjKNhVbUZMsiu
fol2hoN8whbhebIzxeoFwbPlrtBeuC1MaGLl3+o8O2XIlCh6ORJxOtU5UeaaqTMHz/NWXqP8CQvu
kgswYoiRjLVPkgQtU/Z1D7NN5QgvCDUWMQZE6snjDGL45VihrmuISdR4NxPoXz1oJb/Fdl83w7jg
24UAOrlpm1BYvshjvwwNfoFal3wTHw2kdZGq3ee2lL8jWMXeDuTi/9MKjtkDePjs/RuMRgz2xI2R
l31cyKBAJvOY/6+clFCGjw4PqtzylWm2P3+MydmELGyOFEvre2NwXDnhoZsjy0qbhC1bEY91bDg2
HvMue4ur6EHs7oE28EvNn80b149/9kRS8ysdSIpjQnwi1X4pqUV9W21sKRLfRUzfbOwGb4rDeNqX
IHUciw+jyq4kI99diBwY/j2ua0gorpRb/hSpBZfKrXebVF+MZvEmQFdz0FRkP1hRDpsNh9CfLOXG
FvLZylM9xl21mFeM4a2ZrqiU24P4UoKjTkSW3Ot9p8iSD9iHaLz3eQpHhwYRGpwspE/O5vbE/w7v
nanaj2ltyvA1I+G66wF9hZMLk2VpJHvM4gh7naNZjkVgaqmlmlilEUf6hgiPiv81zDseRFfXSx4I
ZINk9XmTE2i1lXgKqA2sB7GpzK2DW2SZ8rVaIcKRwLPUSJvEe2rDIa/9ylTF/StM/3ttZzLBFj4G
rbkmTEOtZxR7tm1YYKEeeTzjwBA6N4PERQxUShum1WGqFhmEeqXtFTSH2QrWA7RtlsowoCOpxlLZ
IwmcRMZm76dzQKpblm1Waq6WKI8ZOVDZlIae1JeE+tq5QfpE/ZiJIYCLSbdSIPkASnkAxkMEH+RT
eJEK1YiWCM3k1EVgTg2P2X48ckf0BB2Fzk7KdN7P5HK2mKm4l1P3n7N4xE9VmTGHPwc6z215MrUF
sMcKeqTHdWnh2cAdlmCtdgC0m+dy6AKEPQlkU93N1hj7riCM3Llz5FYPdd35eVJYmTI7VTDtkKa+
KiLzVc4UpYp7hU/fb5Y1q2KSb4Qbo4i0jurPUYkcPRYZmHmHdypQ22GFH+54AJchVxwMbbihz/EI
lrEHP3224fQzFyQO+VspGI21QgDSVJmGU40gb3W1gIQc6/UlTzCCR1zx8gpfhV8x/ekVmDGjofjq
KXvcVMQlDoOCIfTqW52Qhu0B6WVGqTqgcpZ9SdorM7jQ+RPqRoKqjwcMcXEVaFgl2w3EEVg/UQ92
JWsD/P8RqlGnR+dzYh9VYeZkKBACViLnktRX5AX3c4KLhNYvuCEWk33LzQkdpSV8u+Gc1UNqvgIN
WBCPIk0x1zc3rZFe7dXA1yGzUuwD/ZG5M5Bs6y/dgxbRfQp4MVdkLxTyodOKbehHj8K+dvxC1fo0
J5vuiuETpvMZ+52CC+0Dz7towGBk/SN1cEc6OUyvZ+7SVgX2YreJB/pBjVsE/V49FxIp4e9IK0/Y
+mNj47yGFboqYLESwPrIQ/x7oZMbqfyE5rECmAlzyMhxRV4WEhfLI4bovg8dOrB77bBm9RKw/3je
2RSpAKD6mmAirP9w1f+YGu7gKgfCR67aI2UWRv4D+LfhpP4NMSTB+udCfjnKoWJbQZtltbL49fkj
sqFJgm90nFMqubpRUtG3FraDvtKSgguBZYLeQ3c13DFsRx1QyCMvW/OHqweVimjwT15JueKHl0KV
sNV0tN0dn2p/iaBNX4RnqhM0j/lrtbGeK7a6YvM8nnv2MjXBDO1CFgShIhBfPlh67YHlEA+9nZzs
s3966hy13a/S5OUpovhZY+q03eyUMD6xuWgubVXJ/5BZFKgYGeTAdWMX/kGEykvNnYcrZqz0BqUS
2uAFGztNiju8JexxlvFYzoyrtJz7N2RrbqyyRaYZ3EwErsUiMHpF+GqsDc7C7s15pHYO6zPeGBMU
4W9tcw8/fu8ocizBQAvccYQ0rLewT9R+vjSsCSlTSCYwbtCR3LHn3CW0NTW+2Kl9uZH5aehtl6CS
CR881oLJ2CbWLAhp73uGLw85vzJx3D2KP1sgVAwhH/Qg8S62UKhLJtqJo56LjcHnYuz2UbhLrrgb
sPKPF/cNVELlnJelEd5a77o/SEJYpkMUcXCeGbkTLOaiw3VthGGj37RPmW/Pt6t6uDyyA4wwl93R
2h+az8LsytTa/CjXZvPt+Y9bGT6/MJWf5NOEv2SRb6oqFQmkV4ZTRaeddIyKbr8eBNFsgFUZs7YV
mCEZRfnAD4xviyoyAXf00+cIq9q/Oo1sTZFCQG6y6dXkpqJA6ORsDsj9i4rA5HCW4CcdOzZxDuTS
N3iFAPPvUJ3rxP/9cBx9HMy/AflNZqobbz/hj4BoruaNkMfO06apXMTVzYCBi95C9q9FrwulU8tT
U/mlzV4Kxo8AbBPzlXc/d8Qo7NThtf9+dLrpMBxIU+x9pfnqX3KA1FNWKmUMUod1ARvwWSr4JYTd
ybuza8XeeCqMWpj4V9y6ji3uQKeaqX/nMLhLkji9Ubxu7T2hPjuTlbz5pAtjxcFuLmxB4IKMagQ0
PEjUBKQBSkW6c3lS4RXZi0uN2HpI6YSUKIqp0uOPU/ijkHC45rLwZbYfAtNw1qfSMXBfLg3i2k50
WFEVfUvk3puqod2299I6Veu3J8LTHFzZ6YkAp/UGoiqu1JJFlgpZ3Wa1ob8FhwMoARVTn7KL9ePk
RkfwC0tEiZPxDuLiVW71Su00zZ69HICa8Pp99MyQPxMJdOsfjYIl+mvnL7f7tbUe/qMiieTawL+i
3WRA6WnJxJZuymZ23cp8kBIz9aJ4e1h8hRIJXMHZd1RCbPZQJLKm9bLWhxDIs6kl8HxOuJIRDcZ9
jAY+9YRoKDfRBm9czS0U+yN//ZUUaqVxfoug33E0kKJKF0y2J9IWuGYYWGNxW7Je8QisJOVfOE/Y
/B4yRswmMt2wnfEXQSP9pvkgaL9nJv2Ew7P0cAhy7awTkNS8AnPps1FqV0CgKtd/guSPnNM84JxU
J9x2uFYOUfLGrZTiyFj6YdMTBbeuS591gENzlUVVKIDOGn3dfAoLzjG1P0x2ud404VflQPgqyGu/
fCOWP4HZhmAdtNXrv/u+/kwMLNuteORh+6gC/67Grzy0zxrFZlDup+Bjrp3r59s7O2SxiS2C7M+X
+oI9lq/9+AqGShBNyjLtzUeEcWZOy9KBn2NHoHapnAdOIEl1cKkVbnuJbotx9y7KVICQMppxrrU3
09KbXoYxah/HP5vriaaMGyDtBAWGij0344aqbGEcoyg7iUBOG/9cK6VFAqt4Guj0boB7XJa2ocoa
zKkMcUCYMPVKjhLOusVfENSn0MxvXYO0HJXEE/l5AZNMSKYfIm40iYxzZI3nhMZyksyl1n50FFq/
9peOM56mu4bAKjrDa1brUpRbaLV97TiQ+pqINuu/dqvJ6HfYZTUpDYJrX38jSfrMR8Cgwjdsv4vt
Sqsnze69sWRxdIBSobkMuBdPczaD8ATUCZrp3+7dnGgIElCxj8omgWP3xgeqEE5/8IHkx9MRysTG
pIZMZCX+96m9CRDNjFBdubi4kHR683jElPD7FDvKOAdHxs8713SfejUJfXpRicim61bOYMAvbcfk
QmnrZEfAOcc6tR+LhZo6oAb10Py4ZHVpFhpvMkpWQGDnmRflHQ4KFC58J24ojS6FV1oaecty4oVs
AxRZNUtVwK1nb/mSXPzsYh0tu8D6ooZPzGXsUpm2j5tyfYII9b7i0GTd4Lr9g1BkTfDc2QH5QTqV
vBOoU/wqKzCA75U4+ZLfXf2jFCt+zQGchGH6EmD375tr848Qn5phqoyFpIzRrEsgJeSFMC91MZnK
V3SMNeLk86/+ARFGLpS2JJHHJHefvM6RY1FtGnSp6ggfjQNErBEXX+8FYbBn259S/YhooRTp8AIK
XmZ70uVdbLsMbvZPnb5Ua3dpHDk3+ulDWR+56aKvlFHjp0R+1MmxzM+2lVpf2vl+czhH0hx+Fn4R
sQTHsuLOcpe6ULMT+cl2lFs13msua1jzS+747DNYun6XnpCDvy24LEgdEnNwfq+hp+Otu3+uLdYk
FYVxg6BVrOdHMPkVhYcVJqaTypo2vcVNkGga/GgHwX545VoaHw3YkbAgy1WPA7Rn6zRAFZOBJ6wi
TUEE7H0FoIL2+OucJDMtpECGEZo37eIbE6+WB6APj7aId47b7B21sgIclRNlafyB71qEVt5Ktirr
iZUFoqpWEb6rbHSoxatuYAVzJP2s+9JdhxLuItP9CAYJGt63vwkBeEJDRWUp95Bg/UPqMDTG/I1D
NxWZK/UO5rykENk+gNRH5zuNwDhGKDLPvVOZuPeuEWaGDrsMPVPZxmL/WmHP9cYeBnAT6ihB1/fq
DkZk83t3mhZ1Qe1IcyJ7Swk0/HCyxS/ecbhZ+0r0+Q36e9r1oEW5NP75wPIgHaJUUF/aBpjfWyfF
wppwKSncz7FapoZk5YWqF8dak8yHo6TD3GW/8Cnt71pBRG3Uj9XKEtCedSTkWKyZH46UCGxvsWRN
dHOe1i8o52gLx6mzdD0slYnzoBeJnpvRHH7tPq8jBTDaCMetrpcGoJSxNPOLL2xN8Ew1+DqzItSg
TGPKHgVzRsd8hnyAt38D9FciuTdq2Mpynujh1h5kQs6vrCaKq7yWVDVAlX/Pk6txW5rz1j0T0PNG
QslOJcX1rT8SfT6yREZPN4XK4Xo3cWUAQDFGmyIW8Atvr4IbtoN2V1NUMF8DcEvXy92hBUZHZ1eb
qzN3kKStuJTrkew1iRMVMYB7xIfm1P9vcZkRz12SzGwHmLdGQdH+Jii0h5/Rz1PDmts0naD0pIlV
HYtib1pWQ/QkbJTqCZKIQqaQGIWHC9mixsnCGWx88fEzqq1zFYb/AYNCAREFwAiFU7Uz62Zm9Dbb
rRzS/De5zHkY/CxNE5KN3Mxctq30Wiv+dagRs+trd+VNBqTZa9DLATWXSrrwV0y/EV2+qqfbUAFf
IG4Oyl+dr1kocySsqb+6qFlN/VcFF12QPEpAAzq57O+g8bqPkLu8+lc0C5OCabE+QFNmn5pKtyc0
3F9rDsWY5pAvhXYTuasrpYYE0YbWqUdog6NPvq92ywdoQIO4JO4SA1+YH0PXpYUYCGiw2/WjFart
gJGVjH9QlKJmFCGiRSeE1r9JDnez1CeCRMk1cRFpMfaHdnWlNXZcqUwH1rfhxvVNFsg/sQlPnOCN
5aSmyVikPBKtP2U8pHAtvRCCUL+7dteC33XVai9g0YtQU0ZbzGiMrfQ2rYskh/kl3RAcnfvR9kXq
7LkKso2nhXEJmAZqfUBOsaI3i822iTFF7bW6eFz0oJdHILKyDDUC7Ycdu0yGoqToZ/QGecge0uuz
8CKCh65pEQta2ZIf48yfQVFPHFquTmC1Isx3J31UrCl+tTjvjsZinnKfKGCypE+yzK7cBAoQnAyL
oeIuzRdkmNdDFxOrSIlF3wbB8DcBC/Xe/2L2AhMNiwemkMnv+Q2ZiHZOTKvE5ReSZWoEPlJ3SqZp
G2e1ruIh2Bca9Qme/yoFVgok8i87mDPreA3Pfbhm0arIab0PW1q7K/oaqicNcxgsw6pL/ekv2w4R
ODBYWEyX3THrkGb+6aJ838ozw3pDbgNP36SANwAOG9RyutIIwpKI/UrVGOEge6/foC2dnBZbQxPT
WwWGNu+H6JrOg3snEZQ8/uInCMVfjbD+7TnlfZ9pUP1y+ibz2ndEt+IJZIlDJsMJTRwlxpd1/bg4
miwA6REsHr54Csdi9Hpu9KaXa3ch+3I6VHE6wDRGBmC1t0RE2aiIwEnKDz4CK/10SoVIZYQuVkvP
fi9N6LxgqBCQwKvcSSgt5XffVAUMZ2X69ZsnBqOsJZC7QgzoghF1hpxQrplkSQwC4fbrk0Sedluz
KL1f3gi6wteDCw2n4Zwy3sGgQF1hSaMOkFxbuKWo+DNGJE/FAVI5unJvcqtpsbentcBQ6oZ0ffVA
ZDpw0AyjW9GMXrgFgHHeCpP61fHg53vwzEBdkihlK3p8DARp/4LxxzbJRGOmP7CpbXdmzJnYmBSt
LaOI/eSJGLy6HpugSarWUMO0dYJt2eLI/SzgDKUiY47TZlzBzFiMjVcN+lyaOaCZnk23nfXp3XZk
X7Q8nLOz+EZuXOk9D5bD/zcgbiL0vaXTtQDf8efhz0AlKvguaFws5rIHYN1gBMHMeTBCNSg2NXG4
stPBF6NJdjb6HU4xktyMOJcAxccO6TGpnbcxLOpAF19QBosxcITFnv7D472ZEEGyQ/zYgQm1nexs
c7Ib/4UKOqztn9bFE3R0xmBHgjTpo6WzdnxPdigMOGy0TLuQt4L+PaV4iW4oufoPfkD0EOjYaNMY
LH/+KpodB+iMQo/lFemOlg0EDzJ62IonhgMVDBWt5V0huYmFYD0tU37q6MrUNDzzHvz+By+6HKpM
tkRN3daAJfyzSxqMUHbE4bPW46bXdCIUdNMwDYICDLrACFQU9SLZXdJwBIuLb9/FEzl+YkA0B8vf
oUfV247wCcOmyZzK2HEtMwbqs5ENrzzOXjH7xg1CEcsbPGWBO653xEZn2SpSg+TghR2nYSefv9um
5ngZ3IzHH8vJyAJHTP9UL6gxpaWqAJ3xRKcGhsvvGlaf0ekJaShdEW44nmKJFdUwOgdFX/PgeYuP
x0DH+HKafgUsmGcJ78u3xIDChZ+uMJ0Jr9QqSimmvUFlEeLGqWiSiyEDdoEpfJtJQxi20DUckRXU
9gJrG2oEZpXo+BF9PaEEizt/VUY3CgernqoYe/djxApz8WiD5OZYXCirQUDDXN1dnijx59Lj9N6d
GqZ5sqdNqHe6px4m29maT2LRifgyq0pfAIBO6G9wOELeCojMCZSHl7pcPUXr4qH/jLCMb1ymxh4O
Pj0uooXKNH7DMUidKQ5yHWBHxzfyYsUXzeg9JMny2gg2A6lcBJQRpCuPuLaItufnnWoIeDJMgMk2
QSJdlwwZ7Cfayo2A4jiLifsO+E9TzHr+hf1rgd+LGykvlxanLcTqse3k/gSSSQ12y3MVFDuBqAsC
kFRYTdJx+1gAXVuErgUK8y7vjkXPH/hxWckNjMZJdjh8p5GviRBb9DsHiqf/hMn169bD1IYOULpQ
oZ2cA2KibacG3MUEgeeJBWWEj15GXV80ExK7Mx6dw19Np4WpJP2MyFUnpMSl+a4XGt91PvyMnyxt
H2cAgDt15z1ZK++2zMi8Bic6ibiOu16yHKtPhMtYRNvRj7lTo8sl9ljy8Mz8LlpRuMs/z/mYwuFG
R15ZM6xNj8nylIxRSS1Y84NKqFe2FN9256EmdKO3paG2ivSxaIkndCiniJeoh4OaeSe52Fsd0ZwA
Bx5Ob+kPu944IYbfZqp/P3tpccrCglaVH+VD1vi0QClYR9mkXR3eKoyR8DEBdt7rlzPpe3MAkp3+
12FD8e9b+RSmSK+DneFwVLRJTHuG+BOKMgYP5XxiJA+0UGtyekEXwlxNCapkVVkAagQ1NPeOYjaQ
o0yy3ZervP+tBeAKnMXd464Dz8hTNZKodPTHxVuDekyGbWvykCfQ7P56WU4nL/JEzE5wZbAFCIyv
SW2TYDKG6n3joDdPmltShIX2YN/7a47vwKOWkBCx6h+7JoNLfSCwcb1k908v1r9R2uaSJGFI6aMD
YhfrQGrenKUOvcOH25rOqSBzs6wlWRjHuf8uoSlLs8d0sGKhvGKnWeKxS4mpHGe3rTDFI3DRAZfJ
mWsK6OGT72BpgKnXl8580uDXWwr3AtgEYl4e9UzfhvzKk7nWrXwPCPH1oSqVZ5PTOF53W9nI+qHF
ZVvIo8cC1tbV8tkau2PozUHD+GOLFLn7x1i/K730GghGRjqM89pHFBTry8pnx7SajgnAwN6Mqn1e
qqLpT7PmPXlkiktaNd7hOu8yx4o2XI4BufLh3AqT87Ve+ko2zcM66ya7epTcT+P/mctniyfTKmpg
dpqNrtoIpCJEwtIzw7XxhLrFRywiu1ClotoyNYnlff0b4zbB7NxFD2p9lHj5Y2gt6zd47NUYd/ET
cIxm82b3CMeEKLlczRs6BMcukj4rPcYWaYoHc9qZAvjgssZRLq+r4vpXzPfqq3zpbpumyM8nPIQN
V1RBq1IuWGp0b7jIaCu7dYJmJiNfsSLWwNskLhHFKq2r+kf+tQl10nBkmXY7lUm5KzMG9zafMhZ0
woUon0k9dIjIHkwkbTV2HJBnXm3WvL+NvQkjN71Xs7NJyrkXSTGvNxIKKKyiRlD79g1kZQfU6OUK
fARfMP2z6z7ZbVomI2Web/Qe+xu75JrYrzQI75cX8na14GcYX9gQpNnhoXiX5o5ZkUJUgwhalknp
GqTgTSmUKzTLFrgYhQgymctf6zHCxcQOxHQjNgOZaUFIHpWjUN9jQkZPWC4reDuGh0Xuc1N7Wx5j
UUa7PiCQu5J3g/rM6Qdagi0fxUjAUUSw1eHWmjLMSLntiYo7zTKRlw4jOJOqVfEI7nQVlBwxOKN8
Oe0brcjK1zmAnlZFVJG5O1/6+GEVGk/JnCLD/OsJB+UbEjNMki33HVAF+gzXX54DOk1dbtb86iW1
5gRRUmPdgu5QlXySSR31aI+1H+TCzpnsMuwtUWjaJfcb1mJkrtRK0JYsf6C3Pzy9WANagALnJDnP
K4CD1I6fyBXgcfSeLUZhe34wtza/EUxvUTtVAVvplgl8p6KeBcoJFxur5Oi4WjHYRKBBiAo4WukT
b+3gKKAL74VrBf+zm+WmaHHDJ7U8mB1IqQ0O7rZy2cVXV5W8YNw2ba9ipktFB/xIGDcL5uEk7QPW
U/mW/03167+A+c5N0MrWtfeZ8bLdy6B5d9J8WcE7zhUHINcKcLWid+qMkB6zZ1Fb2y9tsn8EqAY0
KdUDYo/jNlimZe4EL0dWVIFvp/F35UCrolt04YP3Sz0ZE5ucS6YWrstDKYWIjtEfxd3lVH7mUjLD
LYHVSGPZshCImmzB45tsUvaDlofG2cA8un0OkRQt/ng34bQVIUsRgT6JXzdSk0JOsTwbX52VqPoj
mzVSOsOAtPWk71cK06GPF1N2aGDIr/brAnU4bkbsZzEBwMj2TPNScnZ78ikaC6FdOjshzoP4SNqe
QH0VFSndFs0Bwu9M29UpFs+mImg3IjEw97YpJ92mkAcVR8fejoc5p8IeJanTInp15xpDnVbIQJDh
HdlElvizcdU9nSX8ctl0JQiCNf8DrzUarYhvdcYvmD7bl2L4MAQLgad+g8sdDotnZEmsr6fSVCoh
B+d8E4jHGUeWMf4PgeeA5lZXLav9QOkBJampfH2sBSJPzmSbxN0l1VuJxXy84MtAUxp6DsMXngSa
65kTP/9fmgIOXGsozSUFzetal6aVz7N95taFVMB2bdMaFHPaeytLCl0Fa5JMP+7kQMzvJoxdIiPF
4cdVDH0kf/TkgN8bQZnSP9mlLFKXzRUXsW7TJ7H+dZzP27xtXinwVihjBGQZa3Sz3wFw8ebb6Dyg
hlvg+yt8sWGHaocTBn6zKoOYIW2OGuNsImwP/dPjBK1X6EZK+aG7jwyOx487zxtoQTAHFTPLLv6n
BQDeBCMyiDXYX/WpOZDdrE9fZFMRHY4xe52Ykxwj8uF758W6C5w3TDP3jjWrAsrH7WCj+5+zBQk+
cvVuTv9B+mOnl4vZD/CvDR+CPvAQba6el53hMfgrlAhqEITZYrBy8yIjBuJyZ/CmB7w8CYM/V90B
sMdLUTfq+WAxSDAtaExaR6RsABTbadjm6DbEm683kUNt/V1OSbqoAEznZsrixODTR27gBhT2kUIy
tP0v3vIMrwsAhSZoFdhbuAgvy6SOKAO9kbF7XY91LlV7Ft+TFYPZoCbS9OQ/xjRXHLthjYaonhlv
9DLP2AoVW/OKUbg3Yr5Cft+oaaW+rNxI/pquyqcCFrxwTNq+1vthC96ik2MkRWYl6olVBK6JHCCu
IzAsJEXTo2Ul00JFNR9JIfzKWJgjLHelYWUmyK51XXhqJwcMe8R6A0/Bc/HbkHFHDuAYk1UW+hBY
WqH06vfq3Iaa8700738HA0OmfmQ+39t0kWD2/KD3eZWilSqrzKhF2S9rqO2eQDgR+UnI1YrpMrMv
huPfYGErhl/NjxiOpHdrnQjUQ7nMC4hZoyeOGy9qXkj6xGohE5bkSIfDoyfYx7GI6bmMhiDXEOBB
vWWfm1bY9XlMa+t2T3YWwt9lW813Pm5/OkI/o8FFxHKEPCfjdEU1EgiaSatpx2pXmwJIBgywcGsX
Mc4QBkslSY5RBkcEUDnoNFGcYopsQu+iLnuDUNx+O5t6rv0hPXiWscg7CxFCWF1EJZFJWKIi+wWy
+QxM7ky2egTJOJgWEvNKaNZqFODO/L9qMl6c8ypwA9xsHKzNwz62ERn3WnpilqSJ4jc/5JuaDzB3
Lt+Lye46P7BVS8gLuaFeuID9r3TI34T8g4hlIvMnZVoVS+OukaGhaFYfldTsKslVb0j3/QNv4CRh
jeKyKtLHjcgQ1Sqzwm0uu2VYftqjEcWfyA44wdp8HtwtYdtr3wU6A7K5tCSF0lrL3EMkQdGWV2Wk
Y6Z8GNarcIbzGNlyDqLaly2uFy6jysVPzI2uJ7NDONhn2fIh4GNrdQufBblfv/6dpe+XywyrdAiU
gzJg7mSmNEW3GY83pzuwI1GQNoK3evagqGlz2V3BujvjZHxv8zxLaPARm/s7yQBSVFSg7DbPK3lr
yzRsS60dpXw9gN5RHx4MCzYZGOZFmFBaVw/IYZCxt/iB+mnynJfTRvp3q0nm5W1NYVEscA8YFxXh
6SriV+1FprtcfvnLVq4y84GwiDETiqtk/DDbzSq49LP/9TQAqWrX5bOOeXFuPOm2OS085Agq1gRI
0SfWyTSetgGQV0rO7nN58+vIIZSG/CfiWF5v21SchUt78cVX9Qy4mitLhAD4kMNEWY9lXuxvR+xP
/s0J0pX+/k7cT6WUyVrJZN27krT+12Mgc7dzThMW5wWu2KTX5yXQhsglUnohBQC6InAzZcH+5l3/
RFuGaYpVKUpi7J+4M+h9jPF9HuiwxPpZOaBB7fqzGw36r8W92FdrCxsIMvx5r9FFfLqwY5ouDmJj
pyoFte5Nq1I1zws8MgCBYcWXx6ygu61vhp5Z1CPI/W0foNLtJfggk/GCtgAHR0f0v9qQBmFuAuSi
NgLoSLLB+r1AQ8APG0R8+zNiAwJ+mPSv1X4C9qi07uYzKqWHdljWjQEeTub4CvfThnTy1KiGUzJ/
UqFTB0WURSkBcDadvtwIQSaosmclzhBR6VURbsP05TF8suweNSfalS3pPbgQkoPupQ0ECS7xhNsx
IOB6v/ahiMxYW4eGI9CleytUePw5xVl8f8ngHIVxKcHxMXjvNqr4dVfkI1C6OUTH1QmXGv39Mh6n
vp1vnh5bSCJrjcYcWiiC0Okx4te9KVJn8UxKttVqJf1/M1iBlxomeDtWynvqF/ctmHe2oXr81zAv
UScGowdCLjzCdIJ2xHs1MQSAZWxU+A8d3rkC5uVRLyuRvA3KkJdr5ylFjiSmn9OU1FjpNB5ByX3L
vGq9jgeOEr+AZOkpm9GB85PE5ZlGiyjWTDt5iP+QtS7/uHcDtJTMNVzwqU8PvLiZZM1/m1aC5wmx
zLoWXInK2aKnRoIRyQPaztlu/R5bJDsPesl9TDvGd5Wd7JAWkcOSWM+q8q2K6RzQX3VO+hYY2XdR
eOSuftRq/PfvvsJgmDQSh3D3+5pbP9lYoeDGpg5NGr3gDLiv503LvDoaUYKau+LOBsctTl9pCt5e
ny3hisjAaJvsn5BtkyKZAntx3XVFDByJg8E7PI92p97HWGvdGuj1U5F3frXs5DmKi4Zb1LLHv6IV
qR5l7StYG9YTfC0PPrcXgGSiJ28M+LocoOClX4cU1wIIRtTYXzLYuB58qaN23ghiSnoma1FIQsWk
mwAyGTkzkb4SfRvMOOyzEQ/oHrligXT7m0zXR7Rec2DGFNpYwqFB2Qw5bHzZWYpOY063nrDMQaTb
FL6LlTpgx997OCPq0UwT8T5umevtrhoIJleoYPYW/zzHCJ8hSCy/QNnUXi39d9xb+OEwKRG2f5/R
yRHR1WHrzPP9jb23PS3+mz7G97mEYGA56KIWlpFQfGIku+ufje5wHTs4VN0e8XFjvr6amNMuB9sB
V1wkSsm6qLDc8jIV7UCmA0gMgG3AdUIk/iVm9dKzHgORJLCQn5DzdeqtN1g1iSuMRconrFknNtOX
4l8pm5TIt6Ys7n8FJkD25JUYHY9PInmf1WR5CXi9It18pnk1aZmEJYdqGpGyofgcUxeXoHkhHLch
HLMi0um++DXg54wzJcwEVTak9NUbrV+h8kSPtu+AwRhWztv6MSV5YnwuHTwcPU10mOEv0I69I5CB
P1ygYVHcr0wN6iuEdZYxcXNvHoO1ovAIL4Q0kTYtvZbUHllWpdoFOB04kd7LDEn9p63ApvSFP4SS
xp54cB66pt+vevmXV8P6YwYrJgvIPHG139O4UgvJSqf9gXP+P0BZar8LFNGdRTAbPAwwWnrBcu9c
VgUzrJphRoVjFJvCPOl6lbawBdMaCvAB00YxDUxxxkIcc/3Qj5bJMfZ/TarJ9lcw5peuo7iY5uEm
SeRZ9l9HqBloeVKlwJkfSmE1NQYvcd1dHlNznAZliDlK1x73zcp+qWcfRPtKy9RxTBgWRMgUY+ck
Ah3u8/V0+8MpwuP5GlFmkdVAK171zr5p9y7laBEIoeLO9LTYMROK4ic8ZvU1kSk+DCWideh7eVWX
ZacnBlwlc7qCY4PYBsqBTW09EbtTzRP4svFM65C9qnFe5yUsCZlGljazZN57/16YByFS42yg3rZR
uPIIlBrST7JPeZzk5coxeiZNb0ECK3wAkzgM12WR3fUQgsu6VvDKpEk2mkfhYl8K5ZALeC42nEKl
sK9MxW9abIfvheMgPCKEc4/UWe+kab7TymJ5YRC9A2ZQQsELxYTLmZ/K1+Ie0LlS9CwpVEgQvFiO
hQCMHN5Pzj9TkbELQyj8jdk3SbYxVyum0TFo9vf1pXiENWL4uJ4Cv3ZkewcAe87QowMrD5lKUAbG
Il7vnigTU+a1cR10ypOM0wkBXzcP/j8k4a9y+8kTVl1GmLsfXLdPJkSv6xTUnlX6Hboud9Mg61pi
IiXNbfLUsQDUXbrH3SShnHBcGSe9ppIVyg2Ep5ASwDujWPAVOQrrkXUGYDMGPSPxRMq82SsAGNV3
HWpHgcs7Rha96n7UcJb/VDunkcX5Vlor5cDgMFpPoQ6GZTDsqJ6fgPbqU7NkXst/FDTq2EygD2XK
DDISi87QuAlNKnvGYhQ3eRihInwVvFUYvxfBGo7q5hcKdKBK152ZiFVywGx/xmXVTS0eAsagC1Re
PwmKUB/EhhSdUu7Ilk1URruQL1OATvupNrbEuyU+dx8o8ftOkaqixJHjBEGZzud1MBnfd523a9Ng
c91EhMcPUCY8KZfdPMrmW0g/CHn5a7/fHnMs7bDADJ3XNEYzsgdlGQnn3BJax0pRrMv2/83BuzpU
lPhSbfvtpf0pbioRBpOXG0vAQhFaDqlssw4NQDhvJqms/NFO+TU+NEsXQv+40THRfcLcr/DPjmSi
p1A669HsEz9C60OzvH8vVXrDgYjVESoXLEAC5R+2ED4eL+yC1P1EmJI4uYp9NDUT7NQzfJfs2bci
VYs+D8dfGPgw/LUzZBj3vg+twAoG+hFi67oKDLrBHEiSrmCHl4zLkfXO02AABE87GDZK7G8L7m6p
cYMlgjcOSDZ09VLuknkn/yYWV0vVFyJ5gWzC5q/6DAPUbK0nNMlcYTabsooBJk+I7IQajaQrtvF9
DxWBifwAGDb/yWOm41m1/pcBoLc6iGV2H8DxcI7xkYhaZGgvS7WI4C2HeH0+z29Rf1W9cz4P7nGd
W5TFnXzGBI/dXZvsnbKmyRcJZ/8ND7VehFue9oKxuU0MTY1d15HbYYSiVvSHMv95r/DTt8GTGH+p
kb2dfeQMtjaTSdeZ7rjv3UrNmlMynBAloVm5+3cXe0IPaISk0sVknoLiEoTOVUcNfFH2IFEVC+ul
sek99pcFN6vtMdvD+z2h3MVO9oc0OLdZ2wrmM0rWcvG+UU9lpTneeH/ZssTZla7U4I0JqwOLN3Ia
XETrPXSzd0tuBto4oqiN0Esad5cJdV0+rnDA9LWhf7eBR7ggoOAMbo1Y68EybQlVnCrWewm2YdzA
4qVs7TQhPQxP5YPiST0uIK1I/R6Ct0oNPSCKNt1mb+65j76z8jZRmV0nEfYIWY24cQAxw4usNQx8
QAdFtwDkkBQi07bOaIDvvhEkjGSNlxXRHhfx5cHl+2XJgDTKAImeyheXiT4sZPTVXgK3d3R+gcnY
GFa6iMLPgZwwbGM0zlGTpgpwD3KE1oTz+ht7mnMVQhy4MweQTf3oKCfBM31kB2wumBGASFmrxCO4
AXnTFjBy2MQ7zcACBlFyUDw4Vj1CI9Jqh8zY1JQOqKJgee9Q2HcUNfBHZjr1qQwbGq3ajEP9vH+n
woet04kZK0dS12gFL+n299yPqdgUnhvsd//jWAOaQonqGjlTqUNc0LycIHVllF9CfNdosRgFdvya
4BYuhUF2fJzRdYfL+sr1vhhs54Pb1SF6HmGMj6ehKKRR6P4mYlAbfxcUbdmnHEee81ATcEauiWgj
xp8SggdEQnBBUzG5BtsOYs9NUPjJB8dbjEEr2cncXZfIOQIP2ILhVFM8/Yk9pdNY2q2B9bpPQoGl
Q3sUSn/V7TtJLbk1C7zuiiS01xDvalEIwvzfS8zTleiO3phu3x0H2aoPMnww3MmPk4FMC4m9krub
8uEJrqpZxTeY+tk5PKDgKV7ojTt+Q+d6MN7jfgSoCALY2mRZviKTvwZ1LGvkfz9e6b8WLYM3JIJ9
8yXq96gDKjxAYmO0SzXoYQuQ05dt7soil+CFe1GqIci3/pTRBHryzzu8bng2C8z+9lhYTDxofJ0t
Pw82uLsTwuN7q4wJxpxSNF1Z56PjdAC0ko4coT9ip/z4tbDg46C6BgXBqv+IfPIu/3oxeLKGTJDc
LL9qtCh2J8lKZGDVWUFlXctiDvUfOtnoSxs9ZXyT+HClyVbQlqFkq/Ko3ZqucJvS8HFIAggRsILT
oiAftqnQTjw/r7JAKVQH/TeRdfMJmTWGebp4R0B/EA4Rq3hShBsiLAuzgY8FXMJPUBk2JFHC9bRm
7KfO96ux0RbsTbwV1xkcT/1G0iHb67UxCLLLaFrsQT0pK9091UsB1xtCBhY9ILAMYLleKdpav6e8
xHs9Vbo9hIi1o3AjJfAK288sLSh1vdYeVwxZkkGXgahKiSYJGJuMMra7T8/GPFFeMMG+tfVaePeX
ZGO7cbHJnubPmdqhD/Z9Tws/KtiHv4mZAEqww9R/viUl8khhQZbHbqiaT6oDIr7WoavVOweIC55+
RF7jLN2v3ir4PUmYUzm+A/e9T5s7KVTKKpj96YcyZ0JCioJn6+qOfTnINCBJe0WPFOrgnQKduRc6
HhrzwYfoeXtWsGUWKZzm+mXuck89cecBTS1djo0KPNbKj5vA1Y9lGk0Ay82vgRhBcXoiopWUaz6O
IAOyt0ZzEkUlfLrmGcJT/X4FAsuDyhZ2cURkaRqbDoi7kJHc6fYCnpoHeh9fytS8nhE0Euzy1m0O
JCsTDv0bdXC1ve6NoBvNn3aRyyaEc0Zpd3S4fTz2u8+PinlqcjXoKSDpu2UOPV0znCEcxLx14GNq
/iRkccDzrwXtXX8fdXsb47fKBWLIZZCuL8MChHCIdN1oGVgDngoFvc7WPdY4+xuTo65qqvvCqSDM
awMbjcv3+jAegjXaCCK32vhZh032nbYC0rhfmNuKomqJkLgaHZQpsWAuhO6G6/JNbDaLMYPWGdV/
H2N/6fhRiUEmYBD6Ml7fX1z5GdX/xXKo1IO0NGXtXrjZTZlyeq88eDgNyw4BmhKv/9x48724l+/F
b2VV5OTbJXYydj/yu1B6XMkmgdSwsePn62RQDBLEY/Xr//+3QCgqZXo0zBKZ0XD/jv1qc9OkR0xy
pruhp/V/VNPcLLjNCe/pD0C7idwIEeJUOSabWw21nkAveCwIKSg6IgBKaWX6KLB8wdj1K+fN29Kt
knFGmXxv9i8NEkVwlM5K7Iv9myV0zR9TNspdIXxPQZdLmwCg2aW/FLCPYVDkCqytiFVfnn0NzKHh
GTvn7FpnMRYoxmSFPhu/QafklNMfX0F59WfKvbMHCu4lZCXb2AAoBM+km0vLrQDJpV/Gvtdr61od
2Di/6TogOn/bzmJ50xDjws8s7z+OyroXyDpnGs2D8QNy2J/lBz7E+nu5vr/YJfDC3qFYyOR5hW8Y
VhnIerFFpStAr+bO7LhXnW90semMw/BPU26E8dAq+8u5tLRe3eeSSBr7iVFkolBxtEbWwVQdEWW0
htgTJG2Fj5AjUOrBXlQBQJNyn+woOGilOUPf5qS5weA6iiAbIb7keti3GA7T7O/PjxjeQ4kIWnuk
Hl7M4rimAHx5RRvd2qdr6Cf1pqvPVBlrJgpDuO1ktaZWIvSUhEEmoNEjCNral5ie4BQIlegeIk+P
HG4uqEKE8LZK7/J/xwc2kzzGUsFK6EDJ74w2UPWporaHsAGcZWPYIwndDj+HtjD1O2OLIlhp4zkH
rXfu3Vi5mv7/f88khf1IPOUU5rU4zNC4jejoQrQWxu1GyrMH7tWntyi21550L/tkSghRtEToq3bK
/NIZwwOb7Un1PoRBj8d6Hy0erfcdThdsdA5zAkU6jEsZQd2vS9zRCM6PZXWmT7MAuJuRwPrtoFuc
8WfeOhyYVsB+c1ifYFil309qd9QsP5nzZzYScDlRvl4PQ+XlXzVkGxD69Qf6RdZBj8shsKskOa97
eQp9jd3co7sWGyq2lMC+qabXO33H68SSyh2o+gNJmNTISiezwKb/2NjgpxPtyue1X1ldgvE4zoCu
xoI/WTPzaNiDlxloO3Fk4w7NjNh5KKs3N7YHda7OTCsbn2Ty6QyvFNqzx4t1yD6ZZjSPjjN7VArh
SR+cE5qSth+m2/W2+7gaoHu6Z3j5rdPhkkJk9FyC2QDOxsRieH+A03ZuAHBrWXTnwxYPdtxw8Dac
PJ5ijChX41S6qoq3Dc/2VXFj/ww8Dr2qAPBq5a5FH9vrvTAUJv0zSr2CAqjYiaigvC1Iuo4RowAV
BwEQhPkSTeJ2zjgrW7hb8uOpJe6hAaZsUSUYJlsbcrhKPnJKZysaF5ai3hTibFH6mPjD2hmHV5/n
cf3bFMRWEDsgHaE89YCVxcVXzT3yaRZq+eEshOgPyGshU3fOUsc65a68cdCESZqLoazl2etcaQjx
8IvimamwvhAGsfeVvSqcqiW6MFhVc4TBY9YwLRfuSM7g2SqJUNcXMO/W4DbQhF6F6Nfe6UusuU1s
pA7qtcdlInLdsq2LqqWhb9t5k3T6SEdgmSTGOH5SrXG5zVK76muq5OqaS3svts5R57k3FDIYP4Zr
O8F5lPcCrk47xdmL/51V3hzMVZnTlOHdafMOFR4/afEB4rz0HTrKSYb8bVUdolEEITeVA/pgPnxr
F2qewixytg2AVtYL2FK/pGj5Dz2J6gIUGLXXE3gBIoHmTmxLpZ4P2WGKrQtU6UF8gz/JrSQwFt/2
vY89YIQ7o3MMI2Y0FtBQ3wP8AlHS1d2xFdyPCmGXTDolREN5lqvTYgsO3Q+SEKhFpyJQlf4TSaqd
+Cb8WchjGJgf4B9xXzjuNQ0VAFwXElFXiccrxPh4hna/DsqERrQmAid6W1c+jztJ0yFM+FisOarw
GL6no/ruxig+dmjfFl1LJr3vzi9YbktEU5Y7nFT+jiTl1ykUp9NohbT+3EhfcgNE1O0NogC1y6OH
5+70rXQK7mOcAJnhp5MQWgP0iTryXZf5ioD4Qte+MtgG4aPzQf5yT0UyeARqRwMFNghEaDZIzzST
Uuwg4jCLk9qXTBpYfJiH85jgHCOmKBkJHhGMDkh6cWPSHIhe07cmZbXTV/Hc8GVgel/WuWx9V2Jq
T5xb5u9d2prEF1JCwz7OtEyGT2wThsDbLmkI+YCZf5+1gPeAR9s1evh2h5xv+J7Ez680Z0ggk3zS
/7nmOXasZA9mh3ZvABTv9erTxZo4kaV8EH6I5YlbLbr5EHmLaGj4UwAV4Sy7TImbINboDKDtBgVy
TMtmsSiQmr1wKiuu3ndbsFFtV6Owf9SIkYTa4OkYahuNUK6GjVsPfB7E2cCe177+yrsPuDl4vKzn
ejX7EdcA+9sjm0LXGoS0hpNJ23RxXoJLhOBrtmSBUxx9WT3irnpLYfd7WLF0j1VoLpRMqNlo5wXN
lX57AWBi7FZGLa91Bkr1jyprWFimvh1sCerB+C4uQ5lxsnsjBd3AkYhH70eIUhmGi/fDOmhYmyfS
3NjP1/q/pZGlBatQy5inJSGuK8eTjvyEgiV+EhfEmtt6CRhNSo4otZTw2LYd9LqntaAwJ+bmGJx7
JYP4v4vwiad2QGc92S+YY8t+iWSxSPHFk5XExnnububXTbyYScrMTu8Nh6AMWkJ/u+9AzNyw0h0F
l2+sJRxA9+15DcQ56o2k1TP6U0dasNruajzou2cHtBhQrXNMfjsTiF4SdCF/XwAFmCljZ4yl3rs5
qPgoxlmYa6GB27oZUazSeauB355itn7XjWZxuwm32IJwLwhhEICrpqY5Zmwmp/6O3i/6XkjDaXpO
b7bhDO/Y/eU9W9CuDc6ohszsvQwmz5WFC4gu3sODXV9zg27dYauI25N8XJeyqUDA+N/Rm2+ifbtq
OGJsJ14greeXKrpg0rA7qL6HlQrOqlv+ygfCYs3lkOwAOt9wsDALOBmhuhRe3ZEzOUcCDp8E5/k+
5IbW8mI+cCXZm+u3i5L2/P3Dt3aQxkYQfujuZoxIeAe+bRFbTGgplxSdQLvggx/HRG0aajL4SylV
B7fwBznhahejgSB3+qI1rGvS4MWcbGEjuvsxbFxjalIrqguKcwUXZqQfgqZZUTC4jXiiRQ16Tbmg
Z4nIGI4dzDang1r3GP/WvAb2tLMOGKuNVtW19GWQwkK1DVWlMeOFdRUUolX808mbDIbhj+25rCZo
c+KgL2FaCo0Yqd+9FPsd23JaggaGu2PiNW7xm7YOg9YlhJkAxGGCDpPVE6ceXS5Sd3N3l6wy1NMi
bEJKgRImyl0QC/dINFtv9bR2CxoM5own8EiE/GAfB+BTxT8xmznYtw9mjIDqY5dNnIE8CfaI5mym
Ft+s+0vp8J2u8WnNhlzzYbjrqAp6/adbLZzTeFDGguQcx2letyWVmWCvP1mvWncOriu7+YtibMrU
H2BF1RaHIdmrGsvlXJVF4ZZA6YIzZawjULl4/30oABrAETjipW82USvg8QTuLizuWftQhI3/MMho
C/A6jcHI+t8lCBu9KV40JaeX8DBd6Zd9Zpf2Nl+GkZ1b3Nyz+pseoWi2/Ty7DctvV/Zsv+ClIDL8
YraFJcxBXbWFedcQnSJHxZmVuTZiHU/OcFB/CW6kc8mJC+9miLO0SVGRakEkcTS7f7s/3iRGdWuZ
J/YAV7PamPTvLPL/5Phe3SPu52miuLQY19dYjTI92HAtZqb4KtmmvGyI+f7318wJY8QIpl8B2jSv
4cNTu0WFWGYsIrmMqqauzkJeTXGS/FZRsEU+TSqDUvzmr/FJr8COf/POamGGLYmAFCyWxHh6cYri
4jSliTbD452neOfFJqOcZF1NtTBt+Rvkha8t8eS6fJw5iWEOoI7jB/mAsVlW0v+7mdHviCVT4m5h
b+9GTEBvev6Z/Yd0duBQ0mg7iD79eHZCXKJ17OqEhhD3YYoHSBdrNJelBbwh4jv6ai8QZgLkyy2m
aL+w9l77NDfLuaarOQ98vYjuHquOrJ+qtPV8/3yY6wnGJRw2LaupscxOITsPUG0hXw4HtLxNdBXn
NjixAzF/TjXpuUQDMVP3wtt72c3gx9FX3xoCBBzI33bHWUq6eY4C1xGnBRjkQB8E5OJ5RROYS+6O
9gWoccKkk0WBepnHcreLr15xQSXaZNfyHuAPd58KrUsy5iIWAhjPVgWNCiQdM20PtLGcwuxXg0g7
jiGFT/3FkD6bwmo4uOmiFEdjMjGskuSgIaufBVe4spLVIwqqhzUwGJ02f8X00l5nH7uJPq8SRa9w
dE0PKfGMz/2JbIXhQEPAgkMFs6wbjpD+Kfko+0Vv3MCwTijtuR3DySjgGQUQWf9NF9rDZmlGsmN9
etcBp9jtV3s3myDQSj6jsBPxT05nnBCfbGq76kx5UHgYtBE3u39kXBy05cyca+s3+3SvddEpjXdp
q60BEm7j/9uoH2aAo4hQguKaxZyT8zGQr+sse9dCRRJql73AuUZoTPeqrLew0KVukx+rc7PeYcDT
lHM9IgBHDP8orfAp5a87NROcPkqIkhuFavsttyZg32+tk/5MtFgSkgqzGtabeTierQtftIE3lP8n
nSIQ6qoni353ARUtiWDrhXz+pRQqf+FrxoYleZxsf5BbDOuEDLf7nLCbcDPUvxZDtWsbPF/5/R5m
/HRbiuwvCCiHPmcFxku4QY0Ke4vIrWIKnUSQ734uLsua4LejPbqQ153urxXo35hQWaRPy/dWTkEH
J27FQ8bsYu/IGl8t0roXhfLjP21KJ0BPqEPk6YNghG/+bfevCjlJYcGP0emr1SvK2upqSEC3ZYhp
6EtRBoSvN4gox8Tk40vAf6CBXfECrMdUC2IHjS8PPbiTCjQopeydOxvJGF6yQLI+Q1LrfOVY85km
CzvoYTK9XzTPE5b5S8V9dLLZDtpvzUpaG7UGx64ngikon2ByD6fsgu33y/CV05CoLiGd9vmPuFFv
8KuCkOtkhZvsScADDZjbedV5jijYtv3gcruFwMdH8MGEZ+CVEAq0aJgLQMR9vlicO/dFX69Olp+Z
g8VQQTbigCXQAbGljW1clgC/CIOLI55ngVCnbPMCCXHLdmAdljByCW4ACHKkC3yfCzjmtYdsRQ6s
KSZX2s7dg2eRw4CeQmSCW87KoXXNAgdkprHPB5hi7MTLnRpss0YmUOipoxSY2NNt02afGWyLrwM1
GZj82KmrhRn5jIEQO8J3sa9egIKsXw6pLCFmJN2zsPN3wlpPa5/7SlYzuUtN9vyuD2z4/7+DrmKQ
TJosR3tCH1qRePcRwNPlFbU1ju6xI5StFi/8jR8rGLk2jdHHQarqkfH7NTwb6HGNaGyNnTaDZn0+
3fTxZRqKgboRqpDq013jBwAzvqHRAc3f2XzHcll8/g7GuywkGl+PtDmd+QpRhP21gHoQMY7rIOTa
hUfuJwnUdBxZgI8I0u65PadxvIAOpH3MITI3cIdwhvc66T0XLgC9pqOJTEx5qyZTkCpri6/JazED
G6u0LSO6/SIYD1XCXjYOUeqg39pWudhHlVmOq90e3TlPcTV0Jg26/uMOkocE71WeMjUTFsZh9yau
fcSKZitw1HuDHTYtUESiwart4mcrwQ36MqHyyV8kDfl1KTKltaLLTPFc27vuFo4z+xiJgdE02pwR
QrmNPV+VDszLZN8ReNihlM525NC5RdiQHFZBiIWujKGAW/qMQp2fTB1kR2/6cznYXsMKfCvmmZrY
v75wb3npYPrOGF2vMV76DfO4o++IfqOjFruGytzTdAq5ADOWLDH5IAAGH6oqxQdo0JzuKKb3JL9u
01R0lk2z5ZCauceHaeyiIL26zK1Nr1hGbg+Se6zO3vjEMcwX25bEhPPV1R/h+k0v11KsbQr39suL
xJbiRhxeVeVnY3pIzxLx4gzM0BWtveKwxFT9KdozVl/FeYbqBMH/OkgmpoKX7xmUd7sFKdGwLGIe
bUes5Nbm8Jc7/EthZCEeoUl0MUodlBky5xY+YYrUha9r8n9MDevWOlzIzBIiqwfjQUHeJX6W+fsR
BL8RL4hVAJH98DVYEceRbok3Vz4hvwsf2uXyrKu/Ki8kQTbHxHN8aeXjJ6IFWnI2nTLBc8TvE5f1
Z5rPyGcQHzxf88mwxSKdScU5z4Uf9TCKRteSoLW3pRyyQeWJN1Hj2r4ScdjHHAzzxFglfUaGquoO
mjcONi8HPFBhlTCCz7t4lePHr9I2N8Wacp2LuR1qhqKkdMnY8WnmlED89+NDVKjctgK1cCNHtjeD
7DzrvMiTHGzsUdqyPOgeqxD0LN20kzbi0s9A5wcX9dFkR24WBfFj2EfHBBPBHFX4dvUMj3odyT6R
FS8b1BhA1c63LI4D51STZ6mJI/bp/iWkr9Ih+im8RjWrTF1wyD7hnCBDgo+607CilFyh3+wPTi3D
+6S8ucNKC5GMTHa9UYXz2OP1jmQYnXiqmKaf7DtXJoH+5zMEB3jWfl7+Q/ItWNFfyROkcKEnSuY1
8lOZ8C4cLH0f3lYxJNjgcnUoo5IqmXAvuW1YAl2rfoJZgGWhDi6BmSKTzObW90ejSUrDnSKgZ6S2
/tpfM7OApJVmwBmloHEasgpPy37RuitB9hLrJ9UZieb2PmC5lKWTZSbpLaKhudfzn98Cj/Js43vy
Pzh1qG7IyNLowHu8ghLGgeXvJwub5UrMV8wZfKMyuhHQhWF+p4KOW0HDh6bYimwf2khfrQHK+TJl
Sg+deg30SC2FB8jY+d+4bUZ1+7akRO3gz66c84Ws4bzu4iewuLq/bW7PhxZMTDUQG1pUVvNQY+gA
I8inieodBnXuLP/Ar8TQP+hPInvOQKdLnUo3ZII+M6H7WRWtc9R7ou1+Prz9NZf3dYmo1a63pxGC
tamesuPJ8DxBSHa/mvZYVMcRed6qDgjygRis2Sv/QczIZH2Drp7KPn6ciyb4JU1TL22GEZMRnY/Z
jAqrAGGoVsSLxiHjchcKXxOqNn+uJQaTpSVHBtO5u+pLVbHPyQoYsyQu4nD30g8rc6F2I9TQ4sYz
AWB9dT2ptRdkTtrBtHooGPWqBkDGSEz8pQeBhRrpq0CU1/7oj+DEIVI4m8uos0TAR6dRaQosPHWf
XeKewT2bvgm/ETRYCaNQEpWer+jbpflO4tRphe5CsW3zrsbsE1YgKRrqy2uTrUyVXBl52SCLyOkB
+Gs0SYevMT0qQ+U6c16t9ClYB3Nj4uest5UWkrA3gAK2gniSLAcgP1S1lD3z4kTUbNftjDn0fN2o
7b6M55v8YUZZiTQ/5CRhG59IM7XBWACwY+VJqdFTdK+j1SF4dvRRV+15agK59XHMeGga0n05Zzrg
qVIMyZx47mOoHx2o46WthwZsC/3af4Lnt+jANtcKKvdPdTDk1nzhfZROqtDVEHAqv0sAkm8CdZnQ
mE6HPXswkE7+6ZnWbWyyz9jyRCvrdDE02wJ4tqnbz8IVu7D+ch60t5WmqDtr/lS6iDfpqB7Y8TRe
s6kWisC6m/l1+JedmfaczNKxXddvEalWKlrIGJV/LjWWQ3xx9+/MTuj2UukBVmq69o/DhZu43bRQ
8Xz6awBKNaKd6q7HwYOWOMBesvEx1bEumuFGSLsTmKyFcTPFDGHIzynVii/MGGW80DYWqeMM1ITK
HwmG9HtMqxaPFLLxr96EuMsVEa0zHf9IimeFh0n8+9fCUGrgrQf7Cv9V3k/GcR56x5nlDjuT+PKK
hfpb0hwh3udRJxUZYpK1qcYZh6l7CiQIPFIR0/ec083jLjKdemfHAmkOGs8jTGS2ITadukjR+6bw
cKTKCnhPgM6LL7Wr6s+C6g9gco11FjWMetJlhIBjgIoCVrhxKm8hpOH1Ogndpy4ZlXrycLwDmFhZ
DXVVJcb/gkKUPUml+Il8fRFn6soxvt+rVNWSjRcYokn4odj2PEFcPlLBpamU0v+LzYKizLyieGQV
2K3r0XvavvhsXaQQqULAGCjUYNCG+LZocCj2WQAmPD9wlxFr8HxK5z8jT7dAY+o1CY8UutU9aZgI
n34Or3QXT+kKZkXUmsbRUpUNNaKAb1DtyGvFlunuSXdlJVHH560Kf1AZIJQEVLzF9h0MBRmnMYf7
1F2ZfQD+QGCq2Pujb0bM4rlfJEawjXnzefhIhL085iZInc5Y5ptO3pQzdGVagXpt2a4L/kzsr/+Z
pJzoICgnsVDIXeBnMMyQ2AHMqJC2LItkxSh7lmDQW/AM3FdJP0ESlW6JjkgF2Eyrmv9JyBfTR8bW
2tSeBdDklmT/K6DHMnqYkOSpZB6NMD7SbQxt6i8ae2L1JHRZoO/dh6uWLWlpYTD5ly72knE9ci5E
NLIPCcMEdXJ6X8uPTglMH0ksgRKHxde6QkRxZjpkvNCsphL4ui3R57Pym9wmXssx6ycqGZuLEmld
KM8yrW9XzuoDkA640qaFcLKS4otTV8wAh+4sYR8lnuGSmWTqfRNqjWt8Q3NuApOG+pWaru76uvtn
zTu0arhPVUuQ85VqhdArctJ0r+fUi4+sbZjD05Wfmf4yIPAhictJ6XdECZ42DVmwAsj+WwwP8RY1
Nyob6WyXHtWptQ5yPCMqzxuGN29U1oYv8cLpiSvFwbsfLQ12bX48fNXqOOZeNp/3Oq5EXfJyG4e3
WRgWB+GjikodnaCFGCGPLu3JrLnJFwU6Q0mUT21EP2+KEQ9oj8CCO37ciDNHk8uR4UVSdnHR6/m2
k11wbuFQ8q6eTTeZ4fwzTA/DGpKMXpeTETH7y6Cdj58kb1y4zkxpWrVwd7bnICw0MYgE8XUmCehM
2qz0r69gM4QzqceKq6I1CYeGhZ+JV2OwjlCxkI/JvDM9zhomo20nBLXUsvJ85o1MMdr6dbkgVNeH
Wr6pKbx6hRCxJfvjtKDpQt7/qTbSEiHHLVopzc7ReXb2nNz4U2Ba3vEDvrh2+sJFFE2UhvgGfUMj
kSk7yXxslRTytvR5vndjfxP+mL/3AdapWd2COluMJoKFgoRPN997HU5JVPaCO6efLRlEfz0nIlYc
uXurwaNqti/cppeaTOFUZ5RE5l84Uv+eA1wvtFnyVaR7INW/eb0ZsbGmI5SUkJ6+Gfnxheyh17sG
k6HEwyGcElrEoLbH9Dh7L/jzhdgWXS75+W9jprPq9WUjSnR8S1P1ke/lygzDP1vrYWopbMX0b3jk
51f0cUQxBdWNrTyRQ4z6QcKx4Z0ceCq4a0f5kxDkSHj7xApicGIHKRUQfuQeJtklO2QXSPWmytOw
12IQaQP5AsxaH79jkERnf4PneHoe7t5BhseCdMvJOJjtvck/N1o7fh+kjlIT6TJPWA5Iaaso4VL9
3NvAB42a8rXikwYWT1q0Fy3nIQH1yNfWrDRHf/hXxxdHvW8MX4jm7HTDNr75v770vW6+RM7cYn+/
EjZZ6S/NhBoAzeXHC1RM3hElL9PVsknhxSA+NfhUh/27gfLky7X8nyvKhFdRaz1pcGx+JVhgJ8gH
EEHzNk2h4tHXhlsGcFwi57yxCQjY45qEALZ21gnLDyG5TRXcI8zByY6O8kujW2hNpOxRhXKqYxdV
6A0knCANDe1M9NMduFKAyJ1IbqLZswKNnuV3NJ9Brg78f3a8EKHSqSIoL4460cWtlCb6Z6emqb+G
nX06cnzMvzdm3vnnoCA0enJsMXfcC/FI86sOaDLlLoi77BsEQwMyJ1Z1iGQFh8pG2eCcSfbTe4JP
Je1pwDHID0ZFzOnuUBtps0JI3/wUf3QewjMMWWAbmIEmd3+W+quyK5//ixpkLOnQTZ7/tUGt7tS/
5GKl6maJ5yS04v/VoLqRxCfvxFQDypC9RsJ6+uhRkBPmLG6vJaQEFY8Bv8P8rDx2h/4kiQNnd/zw
N0A86Lboqr6iG988GkyWcvCE0i0IawmfPim3YnWi0MSLveQ10ffWHhcoxQr0oLUr9DCCMgTKVrKH
zk+AAtTFGuEYsukX25Vz09rRtagG0rQ28Avl99lVZcTjbxRO1X/09PxHsH3HqePtU0E8MKKyRIy8
MjuUidhAcGDqYT4nO2jb37SzU1nyxmqes0aUqGex4sJRrJhl+G0PW3vwGJgLsK+RUWJvAUb2wQve
dskydvY5RlLThXSfZLnovGERk8C6O/lS6LyQzzIzdEBOZtjXC8WmeBUQHFJQ0qmBYxI5pmaQYXKo
LJjyVlIF9Tj7IxFoMSmNH4mr8wxEIsOq2C+8HT0wD/Iy3u4dD3X0yKV5/c5iZNvDSG8j/1WbKemv
C0NDRV9bvWjp2Zg/xe5AS/D4Vb4BuwPyhwXoWwjYfdoLPXLLwqSGNxHv9OW3aviF5Q0RMDhHVqp4
IiKO5p3Ax+kDw2FEir1X+SQYCzc+Gk5AvVKxcekm0mlVXAJqT4UGpMujX2RWAsyd55/uXRb/ScDC
PsapddpUAoM/g3Qm87ApBtQARdb22pDd5THAzPgM3aXv8IiN00/TXFhn04Vj0AJZbN1c2NvrrekL
XR3h3IMdWkIy0Y6T4GvQYJs9k921QH/KvipYyImaOAWrLJ0W73cZKSbryt1kjNXQvC5CIh2a4Qw8
1ujKZjFeL8mph2//JFlXno1YDyUS6oZfVoiUPLrOAJdyPgtSCFXd6Nfg0WlzoN53SIfCezX0IvUf
PjqdrCxKbyupWap/wOfC2TJKz80vx4Gs68SfYs/lvB0AgYqKfeGZ6Ya6pMPsVweJdFg5q/qY41in
azhibGtxAMY4NyWUsZh9C2YO7qe7xdpL9Tlpkm8yBoZUDMt86AZkTrrm5XaMjoFH+zTZ4b5FtHLs
x+F4hMftlIlFxp7V4OVzmS0zV78G3keBQvArtCYJ+exBGIxto/bd/9YPce5dBjPHLV3EdkCI1IEA
Cjut4Y9zoQaMPt0XoORsBaDE7ZA+UbiAlbAoWxRfgoNsFrCVi34VRS/LWE3nLqCb8J+odTeZORyQ
stxMAS4NtOdRTIpbQ/Q896VxkUHq8OSg6V490XjzXTCA3/4Gt1BvC83YXLhGhmWqGgoWJIc6liWS
lV0oj5c7afMSn7yTv/+NUa2Hsr2frrZmFZsVoq0bT/WeQ3NZASE33tgu6nv2tkQI9SddZgl3Nq2K
Nz9Bwgs9YpTxkWtcKy3XzFje+GsELBd9aEGRBAIiLitGvvw3AZ9T3c/JZdWJMbOEZAsMlNsuo6zp
mlJeRwpv5N/tOMwAehxLFileAih3qEo4WwzlRO6lS8LnIZxHheAtLI2GueTosw/4wYrbI1to4Pya
VkQdU5TPcUAaEmkQ6vijRwC8tnflS7xvpib6gCwTdWZkYyHgx/kt0BJbk+RfIrkXAlnmPlmDUiMw
y3OfSA0HBo12uZvoymTurHYIEfUF/Zdx/ASqiWDAssqgXS5xksp6EWvcBGQ8iVq07pn5Q3t0iB+z
Fvs4xY7omWZwtw5qaMYMO5cj4jKPUtF5ROxVI3gP3N4s8sLDSJv5AbvdAta5dE/pS9SnQvjyGqS2
XqvRuc6bf9SgSK5DSJhi+VmrEKDPrTxxi5z3gf5y15y14P+SxWrkE0VC3q+zFtdiQTTFZ1VRQ2pw
2C3mtAuoqs361wjYCCKUgiYnLgVDERMqPMnnVSw2r05Px2O9RrlSG2Yi2TbbZf7liEnlQcRAI75i
n7dYBjgRp6/gRKJIg5hdm2BzstEsuXY16MLXig71rwGQOPda4kIProb8NhKoLKnuv+uIk5JhOSXD
v8GyLFZ5Hc3eH5BpA10sBDeDxY6lh626xCOVCiLCH9y4DaLknod6qGGtF+QckozRRzQHyCFLEG3O
YeoDj++EYLMeGH4HsdeL0+6spvAsSMh8ow1hbp70oiIkNZdRspWdwZ19y9dZnjoaej+A8R3ly2Lu
QBX2Qr+z9Q093j9S3lNHANrHHx6ZZaGLx/8yKNWMnUwBYmHd9zoZeCP6GUg5VvX6C3+uWBlfCSi8
UCv6U+6b0BoChy7iKaeiyNmk/yPHBj5nNfk0Q+DNeqp78iGG1+CeYzYZZflcxMbi2xzNnR5Q5r9r
IoluKmweCLJM2EWxEvpDRgLYC2zUEHlTolErtOhj2V+ojQrREkTZV464mqGU16zvCHy9/6Utqo07
RpWGaB44cNHyT8NRNod67+WtYOzyuyuVza0eKRU5kJ5zqfkmXncwwrMnS78dlcR2PG2vcz1KW8fI
SzVshw2IdCFEzNe5rMzHbcRTBQMdbCUbi2U7jiInoB2jJiIA8D4PlKQgGFlreSN0yQzsgNAAJnss
gUDiJVqWYgVrRFnzrywvJph5ZLQ4kf00ggWGkvnEMGoIUdKp3hdhsi3+9aMFeEAByvEnLm5I8/NR
IJ3DotyQymA0aAGhhSuCe4Z3AZ8kyJj6X4unfkp/3e0YXbR01Uu+dgueZU1dmNYwXHy2VW9cXbJh
ngsSnBMI3xDwSdepgtGBCrJws2BD+95LsaqlbN3P6nAJJaD/TQF2FYYAg/AYgTFr0QPIwusf+a0C
VZ+kchh9CIdQ4Cu1OClkvBJaZ5i8C/siQc+3nYZQUzQRABkSa0NUt/p+k8y9YTo7mlpP64rAMGDv
orK3jrygK8F/NSmbZMaNYUlOcAvKNXHXmu9/vpHncf7EDrr12rrVFuXhWhcPERuWfT50uIAAxi5A
55Ezkb/QHMt1pVsYaMwiTolWlnmEnG5PiIjC4KezPpS1cBKJfYPmfHS4WsahSPiAYiPmwOhCpPsd
Eii+AsvSTw0KasVReiInXr47nzeA/HLEBGsEmVusVjcsfREIWLh16mDjJ0TqTjEstb6DNIfcU/sj
E+R4o7Ke+XbTdp3WUilSaLJCWlu//9JlraDbSbnM05N2NMsDz9KRGh5KVt8Rujw4JV/5qoJOstvw
eiFGthEQ8FutYzMUex4AUpkPGjkAPgSitPnuocKz5bKR29h0gIABqkDDtZ8OwB80SVXsY1mIYmzQ
S1ZqiXZ3/zP8Hj7FrK5NtP7/BXKGgsKTmqpIko0hKuDmhmVrBSLcvTaaM0TeGh9w0SxkGj0MpDZ1
Qj5J9nV0kH+RUoprswpEBhxRc6oaQ5D2RFBdI5s87ayYDWQu8p+MLztMFuGqT/ggOC70gH9hBuWJ
bOk01kgcY/ZpO6GO0QLyKNGKzCM0u+KhrUNuh4jTExBRg0kwGlZXGU8Jgt/ePhsB7k/MoPmhw1cD
a+Ge+WKkwShCdCGHWAnKyorve21vtsi9T24fbTJryVwYlYctiPiiUiZS7pSL2lyOHBh85xqSGnLU
k2LR+DqeuVVlOR0tzjS1IXbfAwcYyMCQUeZlp7lpg+FNpEsvnNNGtcOBmYa3VqkBSo511C2ztn77
z9QhPBpQINcU1vox9qaKZIno/PPADHLLFi4kPwqdTGtTCzooZ60O9j6xBEQ/OFlMMP1mgIBp4odu
BbyXWlR7UVfbsSXUAe39qPUtZjhTTlZgyUY0V2z+pA1Qwdmq19V8wmQXB/gkAj2g3nMcddACQqje
LtH16cXyWZ/oIZho4rufB0EXQ1Xq2bwWsjrbXSWbmbS3x+ZkHISBcFrdFo+TLrerEIw5jADLt67w
WPD52i5ybE1jBCIN8vdJrL9qbTbRrs8j7l8ibiNPQCGBJd5nBeQfi4M+qlVvtR+yMhe4R+BM2GAg
nRdC6BC9SNZiYuP8LPoY4ENSWJX/DKR4SDAqBeWurn60P8rJknNeQVu/R2fweIyS8XFHpefZd4S6
lMNnMtDPBV/qfAN5vn/PP0KX9AsDAVR6ijzMvMZt46i6njttCBitulQKZ+Ql9Udohzm0lC2JWChO
oEAIPo8zgoHWJYW5aNXIEgbIYHnUMPzWXuhUL7sgGoxdLULdcF+KClBuOyv65NIQxLNfWkYfbDz8
moQ3ipd20VO6VzFGVElClyBU9EfgiidXaIaoI4p57azzsfGp67EZ9ETBQbWxjZr2BuYDzjTmekld
us3MFZpkV8z/7c8M6Hjk55igycjw5D7hyXgo6xWbB+IInS1rQWmihatnNFz3BAR05Jp/CBwP+OXz
PjiFiZChNAP3ODLSWfsnYFb3Q1dSkj6gKJioPxVvdY771monaKqPvu+5acmLdMzbv5A592dOhmAE
8fjYG+43LoqAatMbOrblUe2DKHpnVNccQrQuoTEflnD9GeYixv1eEjRlZYIG2V/0Xfi24YEK5Ws7
IyRi6x7X9vELkUIGBl9spVZd8buUSeNMKWC29poWU3EEySF+jQJ/bsCui7jJfCAkJTDUm2fP4kEZ
fTNb8HvdCIrIZAhu14NthxcymL2SotDiWvA5HInX6ZrrYMJOq98ovV6/uBg7O8cJVx3bDGZcOrD1
cR0kmvYE6UAL1Ua6UR1Yk6qrnchKWs2xtK9GK1y2Oz5pSxYX6V6v4npnzSg5SE0BpSrn9L+ztT8q
QBiNPONamSNG2KAf/Ds/wLx34ggD4tAu+TaFYd+mtWXfmry9y55lAyHZ/IZoX6GgUY/h76q00q/2
FiJu7F7C93kim+P3bXAzYdUshobkghkVrzeUJyUDh04UZ5UGn6d9j53a/1RR3TiQsnQdXdGDsccq
e8LbyIigWC5uSYg97TtNWgTG6Kq0juSFzbpYutpiIkouzqqDt7SB2e63o+vDTzWtcr9oGp0Y26Qy
JwhadYII3TGL7C1/8QScTIp2Kujr82Ob5BAvnt3WA/QZvWmZcpTQGVSvBc8ib+RdC4NeC/lQOivl
9fZin1OSASokwY7sNeC1ZkCNGd3XEGTE0cdnMKnLZx/BfJXAo5xFV6eu51mmTkrgzJ0uEhady92q
iKY8CeKKMAxTscJhqr461hiIQkY74mhPh+e9zhqaxwqIUt2Lk4gFXdjx8TwA3I6U2sqrKxdL87Jt
7ZRqOHfZunMXBdGXlFzG3DJSL6DnyHY+0ZzxCdh803FHuyRnXBXDH94DoOzQAvXIkUGL5/KM6hgc
v4dx4iH8J5VnZYKr7g29A2jSCTM0kMrQQyByLztU27Tc2xMOMJEYiPaFsUlgd3OR09oMwtYfLV/e
DxzNPt/y/0Fug9MMgQjMKoYS2W0P6ogqm3Cr/OINI357Hb2Duq2MrbwjuxCfZ48fPG6UqUGen/7y
2Vy1ROcfBpatlQoJw0mIY1weHLGQXgtRYot8OgYogwSVxt/YUSYJJKREZP7O2KHkvtfRFwE97sqa
9BSGetnJQSynkxfrMUyQjy8I1Ew01H0eI0p1nBAUSrKJmHJFg1FrsNV5mbTr1Bt4rd/nq0f8EaPc
nntgVX5S2w7vOVQT7m4h7jMPRD6a0fiEpq+GB5ZuyBtzb8JyvpaFSTeqg0lR0y0ekFqy/vvmL6Hm
5IuEwcQQ934K6BednRry2zVgjnePl1IhC9ts8tr02z8d6p05dZWzSqjl1nbXg2T+gmYp5SdfOO51
iiOZ3rrobNtTZVXknQ8vaIxTA1JOUmz5pv4vd8wYXZ/jrK9iC4xA5i0WRnpFC3shaTwcwAW9Phwr
u/nFcKwG8SdHYPfTxXtUQDfU+yQZXzO2psg5FL+69bdUfVFXwhmcSlc+k+BRVjgtMBm0vFVRbXBI
/pn4i381dU+pOj0AXTdx/GlTOSdDPXVVasVU2NyrrhuIdXM7ALFF/y5jcBt6iXUQxj4JYi6nWFjV
2SN7SHWMczPsUzNKKFhTLUuLvnJt1mCYAzyufJwzgVg7vWMcezZgCqIGq81jR/5iUTEq/1wlQZ2O
bmeoBDwF2p6wuwUtRACKgLcK39tesDFO2+cFPYW3KjPcSfpHGjdxnxbhssGm7MkJWud+SMSCoNJa
or8o7yxOnnvZ98M6cJziDiPg9Nv/jDkx5nsNbfzRGf7WxvnE//9dfIgnwJnijTxK9uGjJ32qj8M7
GUg1cFREI2DWExy/RhHTmiLX/E74OTt5uMOC55kKeh+0KrCSxf8DcRy36VCBBkG9yscOdCViImF3
I1CViBrMp7tcbP06r2Ar3Dtv80ZN6iWM/BaWtQkf1e2cJu9Pr4/Uln69O0jvlkcDd39GlfhlPzwB
N71ZiMRUYgO2wpBXfYB7mnf0tZdZRYNnwwasFXSO2iINXce1BNQpNt9fIzBljiK7c6POGgrwq4Ff
hvQqQrGMaLVTNJCsRHT/eGmmTOGjb5n8MYBd8lrNH6D2iXnSPsl03VbZHKimLHZCRLtyqAkQ/jDc
0Gr8ROa79suVTjt7MN91pM+J+DWajicq24xpDw6dZ7PKXRKpqbLfKPOle1pAPZlcs651VS4MpfJP
YVWoPadVzjcpt+fVs/w3guctoqXx9OHGRiBGaVuQ9biW9o/B8aJ3p6U6H5thV6pY/7fjU53wdqDK
5dcoig5hRUPiWz07NuW+saxrJj9N6R1OD+Urc/xLcTRpjtxHd/3bB8S9hdVQjnHVz1DQDzExb6Qv
RtPB+owp2zSXg820Kg6y06lvgOT4hApln14wOiPeXvuAFh/H6rdMTO4MJPO15tt3GBDJe+x8r7Fc
Dd3cqZt7Bd3jMB760Mxb5btH9mLXGNKdgay0qoPD+n4KTL5WijxpE4wtbbaIuy1VnAHjJ1TEP8SZ
kbOGzFlzdat+8vzy3zUKKntdqH944NfIDT9uj/2URxhN+uUUvZS1wqRoKLyaBHvH5FxkLZC12QSn
JkgCqFiTbYXcwnS3zJX7vDf4XVOnPsB8cDWoGOGdI9d0q2WH2ZuD5OT4I2Kw5N8iSCosjRkCpkzc
zUM+eEhABNv+j5pvYpurFRcbPcveaBo/YIsvC58iroC8mjzDw8VKzuL2BrrV6P2VcwB24B28aKKC
6iu35bK3fApbSNokWRg97TdzlNywmsHuR4gizJKyaz3gRMZCXgDbeGTp4QrVWVJbTK89yUCOBWhK
+CO2R9hM378nPspt0CBBCHJmY5rbTeXtXQfmVz61MnE6kM7cVR4T/9jF+sDArdasJ7XGVmQ13D08
cq5uKmRtxl+ZG++BmPhibWjO7PXSoWppplUKo6vj2nJVszJQmUWRdjXONt/5TQjsYuN6EIuuFVNQ
p3Ngcc+8xmNJwyR7q5VjpHyBxwblg52ige/9LmTokR+D00HclbBDVX6lxnI0UGf/Hv+iQrEm43st
ZIUntPzyqddLhHLmmlQXVk3snZfXrmrRrTVEU8QbY78bLB8Xl2sTVPpJM2ZlHB30R8OWln6vDsTd
hlBpOkI6x2+q7oJpKaE6ty2Jb/xp8201OkDoJ5kyatnGyMRlgTIbjdrl/XKV2aNnNvVcFs9Ygh/W
i6g+mstk6/Q2vWAZR/rJABqqpubKxS4NhEM2f2KF/epn7ffP9ovUVdXiAiBdfMoTrCqbesoInDqx
woCHNJ1Rv00crZaP9jbDRO5PKlWnnVYLZ4MvKpjjpYaNNGOz3Q3Xg/i3Bu6iRpwQAjaRufgRyvm3
4axxoKp/qI2lia/8CINndx/f7sF+97810AkJ3/IjSZRPb/o92/nfbhQZ2lbHUTyCrmGCexTFsy0j
L+tOp7YbCEQH6f4AGH6zZfp9PqKQVEttimU5wsgRdsAohgDVkRyryxpSsXX4wbb/lZa86ODw+iPD
VnLbIZKW0kNEKQb2Z8Gy3nrj4bov+6RpxfBqEWqeJnJAwmFpXcQINRbNxMK3Fb+PPX8Xm07IICxO
ZEdwnIKuIhRF+1IpPO8kRFPiojLgP15d2s838zobxPBvtnm/SufQCyH9AxhVqjEkiIUI4C22/H9k
tZ9cma4Nzu0CYTpbI0rCF1tZ66+vRLX568HD0G0mGwHXvVtKNg/PTPDz2/GGU7qO7TU+rFxnWxZF
IiXqMHbm0P3u+qdCEFNAxusyf2F1h1LLPojxcZ5QEizloBysWUzjWzuvy2csTGR+uPzwp1zsdMRS
JWsHFHwub/pMjdcDVnZgrOM4Yibp7YPeTA8RVItCd9AlEKIR5jbof8Fkbxtv1ctlBLzawcgufUmM
ucx+jh+OF5oVrWdJ5tSntFHyrn8ENDoPR3LF2fRo9AstZo3p/meE08JEFPA4wHmv2kkOC9iAIrjp
sYljcwFYLHfeABzWXs0IeFgq2wKYcphgXxuzqt3wFNs/lRQrgSV32iIQMdphVC8CEygfCs6R+zmo
Pvp/tsscBSueJuS3fk0/qie9OjMwLznTVNUT50i9eRHgh97cTQajKSq7RT96CNDBbpUhVPuqynab
2p7BFDwDBC0nIjB4X/NIYs593etl6RbZGLnlY9GlZ/vXQegU8sCthDEVscePArtl1yxJ4hs5jVeE
oSdxJf3mkYN3YElOY7/X36HPyby2xnRFMB/unKlCLXAzYaX/Jo0qaEEh2Hh+Wen+wJk0ekLGhFyp
+T9bEW9agrlWyNf7gnRCobEmua8l9CRT4obdDKa6Gzs7txstWo6j7y3I0qk0+ZSueiD2OZ4SCLXm
tLVtgWbUQ0HR3wWi0i0RdVKLHebPBY/AtlVujra9kkSGRQFAuVl9l2M2oErjJi0e8VXKsBSNi2Lt
jYEQljhUH5ODz9Gy6l25X7d3cLvxnIU+WRQYv1cUPSc7WU4URhfF5Vuy3Flgg4+NVLE3YWyX6Ri6
MEFQFxHDw/qCd09AO+qdnyNnb6RLGkjlaC8RR35DYiDWKZbcp+oqSsQ6iZTr1riU383ZWpfNtCo2
nNHvKKVxlKaI2bJZ46b6KFtR3I81KfCukTmyilD7mbqsukP2QuvRLvkTfctBQbQxC4UbPgaf9RCW
8uZ+IlH9OVFiYjhobqlYblor+fYo+n5ksjAJWDZRGSTaDwdFZGZrmgdWyTSLZSquNOLqn3bgUBDj
4zX+plVmHrpdyhWBiFJI8ap/Dcc5kOyelc/Qjk20FvqwnDXsQUESx31pXNkkMRgJo2s6s37pgt9l
DRAJaZsdQtutH9797TDrdybed1XB7YxvOLMHObgm6doFKqmwrZovBOHpJCKIqpg6+vrKtXgHtNfm
C1t5FOpocU43Y7Agmu0PH6PYTW7PShd8qHAB2lwqqPN8IBD5xKTb8DmG7hpxP8HAtZ2j1bj8WRYU
kVxm/kFkAoiwz3+AlEI1P4L9l6+j+g5VJkIx8Ge+K1nUqVc0KzRR2xYRWsLufO0rfTl6Zey69Ra8
H0SIEO3Mv1/0YND0OsJNVKKVXOwbc+29hm6qPyTyPkyDCH07ZiHsVYHvYQX3vGi9R1Obd+TLWObz
I0Kvei/YLs5vFmp4RJWpbKIP3tA4dgK18GTYX0/AQP4eC2DUHFUG0z5Bft1AMkBzNQm3CQ8HAyJZ
WUbEF82nf+UInDm3w013mONT6EsDVphxFFG5MdeO9L1AG6SYvv4HAyyy8nbzBKg5tVRUR0c1hxUc
nGp6at9dLpsG0BoFdHDu/OzMDVXQTI0xTSRR4oMGJbWXLCvdU/sNSPhTNaUuqaerturygBMHF2Kk
2cUEQz73CfGKWT9GimkipecHz6t6vHsgbzNMsajxTlE9blAk1ezgErtuqJwB8ozoQuWltVvxHCEo
tqOSEJMkGcnrYtpIb4FTpmVX8QCetrQWazwyK/h5s0h+l3YBEghFfSW825tFZTZ2/cgFbBvxtw4/
XebvwbZehgN0iy/jDkX2HzWyWnANnDAuvqlM+dUsVvTZldbOzisGk8tRj8ypJKzzY5ghTFxNbP3v
s61+lwSceAge9xp6F4jLX6fNU7Fib34cX9ayBKZIqKm7Ir7H8ChwXgR43x9UClt4Qr7pxfNQRyu9
z2/qoZEm2gRC0cTmPIPFeNdNAAgwTBEdEIYF6OEZuwBymjbdtYV1zFqKD+KRrD6QHfQZAE/Qho7b
NFVtttYlswcnUHmrwSQaUsX4JTaHk91LjHjxYVLWEZiFLuv4sjZeNiBEB0asR/KCHaR/+mGjq19w
DtihLTgZu3E6bREEYuanK0q9jXpXsAsN6r0bo4pLT898i6FX/rfAGQCLDg1kJxzg0k2yZdJanvhF
StyoVhzV7qkGI7IX9ylV82QDk5RE81LR7xSggm7HkehrO+hDQt1L3d3sYN7Pr7hjRHYjjSqZ2RTh
JACXmiDg3VcJKMdpEi4t//QrXAsa71Uakv7alv2hZ1sIedvkauk0Zr0YE2xIV76rOspdf+pa9xyu
70b3e9/+pa7pT/p7A7tX83h/qQhjksGJuXBER6cCPOxgItkcg2NHHtrhXWTnQ51nduGJJxTvkLH7
1hD89aQYDCW0uNwLzfSBD/mfl16BR4EP5zUVoIdxsWnlKg6uXCD6/4X+XK/D9oOqErErmgfTaGmH
XZJDoNyq4tpvm/hlaKULdOHqVPMey18wrj+QatubiANO8b5wjOL5KzljWTWK15lXbiCvsL0U9JBi
ZSk3G2g5ETWTGLLwozH7urN0Y/QbnteBr1xLH5wIyivanp9CcXVhd8jYt0hcbuco5ccwjQtBKQzS
MRxd+T9tU0rMtnuWQ/lAm74Fx3GkIO4GlQtQybukijJhRvgUoRmj4Us9z744jWLwTh4J3nlyZ1AO
aPfqubsVxYYK5Una+WfnCiw3SqVVoUTmSub1G41qsRH6F6mu4CkgPeINK68AJeimOrAufV9t5TdW
v5K3fgfSg+SVYrrQ+xkzi59KaT0To8bd9Ag1iOjhqmfO42JEuaIdONNl63RIq03duVixJhFWAsDo
gHkrIBDBnME/jH4Rhx6IEN4RqOTdMU7csKKq7yc22h10nE6xkeGoSfyRZPCo0IP0MgufLnGDMRem
14pzAuYiMLD24ybxNKB+TfPaDx3PTQGKbT+fnkAJNkg0hv9k4UX5dP/hE3fRDsT/h2rJuwhQfWF8
D6geOMC6BMU3x2ODu9MX0GN00ggvLByDaWBuo+kNybQPIGIKP9Iq6JgaECdoVgplgoLZIVuTixIU
g12lFzedCd3q3pjkLydL9twjXHdrHzdHF6poX1qHlKgRfL0HPVnxcj7SgZCbPBwEfBHdxUfIF1eI
/FCJBnEzyqdwMNUHnfhHFIzDi3xklgpRmnVDo0pgkrNJw9K0a7EsjPfqENgmyztBHyACpQvQzn6G
mYSmSjuK3G8K2wlqtXe1e6c/1tyuGpN3+EHBCLuSZXf2FleDpFX7LKPkwFOgGE+0/PCOXHeNPWC+
S4Gc4ut7/Fm6C8Gl0Lrj/8uuDkGm1QR36ctrqtu5hsGJJZRJjzWqVRXcpPZ4Ee9657tnnfIauIKZ
OmUNiZAFEtMES7ctSPLw5fvA6GQSiWUGVqkJWuuVL9AQJnZhIiSr1C3C4UEREsnYrwklFqy0cIyq
VtWWj+5M2HmA/U7zMaDSBn7uAAowom3jZAR+w+ZK6teFalPtYkEpwbAf6DyhCgbLuZVLTepWjAUx
CwTp4FSEWWjU/xULqIPOrgvYo1x/dj6I9srkCiuGKcaMYBQTPLfePSXiNSU+SpqMscjGAZqvF6gG
YOD5Pvmd5Z6jA9uHID0CT7ntCJ6PdGQEongvd84xWe318AGVvOii5qS3CH8BE+oN6NksBCDLpuWv
Ivi8YIQ5r3VpotKSamgGkxDMfPGoMeLRrFxUbhxRLOhS+UBQ3QfTUXHO09drtq6P5cMyS6AOlx/v
wAkusbOseGyH55nHknpvIwG/oQFi1FIvyL1g6WbQZ/4VT38rsonIQ184oUtIfUhNbG8W95G20w6f
20gMfWhi09J5WgvU1BsN9Ed5OiZido5XnGuIJJ99OUv7jw22coJsJj3ERSGFsyXr4Ihz6nVcza9W
q9AypFCpcuPSYn0e8yFoa8SlNZB7AS4w84tmJNb22HU0oM1KVV/mPqR7cpVGcVovB6t/WMePjSZJ
1grBC1MgoBI2Je1WaastL1PRAhezZ4iKB3tcWTsERI5CusKGi6lM1Ny+oRMaWRpXIZYZafiP9wJm
VOob7hwbAWdCx5fdmO2XMsKFrNmQd80DS4CSg13uwFJmFkL0w/t2wFxkGuA2Q1kR6qzOnmIhM01O
v1/6JXyd4XCXazN/yPrSWJ6o/Ic2bARc8V0UUcUK6oEEsnj15cDr2/GLCFgg5u7TIXU4hNpIp0wb
hyohRFZS1dJWW4qi1azda+I21zhDQjW5QQhO9NkMk6g1FS66imTmqG+Fq7fJpDvfLoWzwcL4Sq17
SO24cQi3Wlv/WQlYul1Q9I56cpUIcsZHBTZswvmEpQm8E6697e9PMvEc2pL/3gzrBgu2msFwMgKK
9rY43C9ltbDfdJ/faQg895HeDmfXEWvqsAyYOGUwAUk4OIFxr3wQmHB0ITPSjfJe6yFrfaWHh6cQ
8ekVU4E47cNcyP1HFKwz9GER2KKiCxtsht3yiE4nQ/rFoiYAC2RR4E9LkzSEFueiJjCqmHbNbIFZ
Ev1T3LgampVt/sndtEGxaDE7h+hVe7g8GGfZy96C1vMDTrFOVXiqytZ34Avk/AER/YFV+cr4EBx5
SwqrtfqZQALo9ac4eLyHegydvqacaVg1CTlpyXJo9w2FND7EjLfBAmNbipMDE0bhVw9DZfKUGGLJ
wlPcyhxw1Qouy0dn2sntpYfEwHBaJP7vAfBSTIl6HzsYoIgZIN9AHGff4XnI3t7ltEkptffuFxNP
S21SopnFu6dIo3Ami1z7h6GQFJAy0ts8Qt2CYIYpJI/R6v8r0ulPPh+DalUK2KmM0/DJ7qqDly7d
1N3tHg3GddWFd01ctD/K4zimZPmjvDuybo9PJDa1vgCPE9mG4Rqw7RxS/jZAD3AseWGh+KYU8Nyc
tfqpTPWLdM3oLcrd1lly01O5St1+hGzOObeDiVaAKOpvxARD4P1suYFR4a5Dh44wMMM+Y+X9bJcI
yO4/ObP0CwYYC12o5kwf5NGolZk0QnrwMFMJ+nvlceDMCSJ4Tjbk0js3EXXBzd3amHQYQxIjxkN+
Qe/MWJEgYs1LzaezponDKNJZfHxhRwa7fTr8H0SlLz3bMGp/BXcdYUwkdwQ2RUootQ4p2hZenYx7
ejHiIm4/t+uJGIvnRCt1+prgLY3qwZax/G2rXO9ZG94bbtEiRH8B7+5XMpR29Z0DMYNjPvM+BevA
uA7M/H5+BEUoKl07hpNqOfUJ/AZWQoJGf4Q87Z151SKd8Z8flTag9NiWhIDwrOyL5xp7ppWszIIz
qiVF6Soxv8+bMm2fzGognaODScOsRWwuyK15B1/C3/VINh1J/bSeY9by0e2gQ80Mjp7po2zQoo7T
4wqUHTHZVkn1o04aRKhhSw/nbQbWEOHsJO8Avm3LuZeovx9uw2GCAiS3bVLjhzNrZ2EQ8qOFVASC
idM/8qy17pE1y2UdLcBGOEfQbz/KryoR9yfHLafrPRPaXC44smeCBcG5I/kjqXcZ5CGEbv76C7+G
wIzaTYDL3E6cRXr4EkyzKh7YRp2ArStjHQzPcnAdn5Eu8Iv1Bj8lfA3iAwxlzCRWjEJ5Gc9WG278
y1KbIHrsFbw9Aj87HM6EMdL4wyEcbft+ngCGX/jKASIb2fKBxwvcqPqkWBHdImF6LSqwltui0Jgv
H06ZbhFxm0Y0NwvLkOQftZuP6cme/DyW1nye/UYSCCWDxCREezRU/UbzSlgUegS8f9IK3bGPpeE3
e9jRcG5ZcuY2AW48dvo1H7I04A2p55tWdbwC7BgQzXi3H6ljuLk2Q6UsffH83PvJPHsXp+i6zN54
DLhI9iRX1+ThA+m5NLkCkoctO7YLs001kqUovNJox7zeZJ5nPio3YF5GIkkR9hPEizfHIVI8nb9H
JEexST9mUlY8xpqJMIhu53FdpSXK9178ZwTH1tWKiOVDf1JVbRc+7mt5Kzh7/z+4WQ2GRqAnJNMs
IURXAuulU30GlbGMbtnJjtUQ6vQEuU2VGBV33J+fuWMvv3BdRkWQwlJp6WMSk8zoAdXuTauBKMBP
66DCfMqNI/WF5dgnOYWZqMyPsUS+6RvhpmDiHdl/mgPYqZH4bJ0mIdbAUQqa6Oq9bm8d3qOpNQJ8
m8PYjRDUhYByyLpk8LQbpJDuk+P7nAeFtxdJ+hFlLIM24inD3qEkafk/r+8MDsDW6589KP/sb58M
AoExLbpEMI0dFp2iIxQH7RgIMsq7mPw6nNOOIYH+7aereMX8iXHfERIiF5h9In2h+4bM1+wxF7cU
zwHJWWuvWRe4HJyul8CZ2fk+oWH5qwg6VzaPJN+glZWUnANR1S5hzpoKBxzInNBgC1lLJqpnyvO9
bnBePM4I8DLVrTVNjmonccy4RUsE+JwtGWzUHE/v5dsugn+S1RIeHVGOMEL3W1nXz+0c/dXVudDt
uZtiOQsA3hQ6P2s+xFSLud5EHe2Vi/Xs0tp1XzIN8FQacXULHw12izfCGN4KRWaGoqxOa1Ll5ltR
74dmohxdX8qWHKZj8d1BPVG2nPueMZjrv6buu7T9vWM3pC4r1erTlQptCKcOTTWOpSyDiT0BHUdY
II+sn8M8Gaa130PxOODDFwNiEh0bLoPWFLS6j1TDw/GFxze8rtE+FlnpunfBSPW73cPQ8ECscaHa
xycoZima/54HHMbNq875ZOpGPK1q1e2V/8QGZuIXXTureURfThp0GRJzVed4Yp0AkxbxwjH7H0Bv
uRi0mK4LLvioJwOaCK/kQdUREfzYmPFBKgND4HjWecsDhFyPoU/X2yKbKzW3O0JwHJMpXzy2Unz7
m6f3yKD3tKYlJq3atEL9HXwLngkArNy0k8xeEpcxSDW0J1iYayiE/3wa+DYiDEgO988H0URNUwL3
mvPZJ+HDLaUj+r1Ez7tXEEpR57LFJMnXEICj7nS+DGK1mH38HeV6/nZMjkG3bIXOr3TPL3T8hYbT
/bp/v0GV3wjwz4sywelPQj1bkoAJ3IZdBvFG57gazfm+CXKyaR7jTN9AxBn7KVDoH0OGrOXJW1cK
rxx2ngQLMgH77VcrSxRBG0jDUd9NPid6SSHfa+bLik8j3Jy4/XElChxrf1rvBaFsTmF80v9HYm85
oFyyPK+HFFhl3RQIBdAffgGEIVoEbbv4h8W9NvLnKzZDtoM5PqocGeIo+rJHPlq+8hzBjnzlheZQ
LGV2+TnNDTs7MVl9AWmSolcnn5VWrij+TP9j7aIMRwruijGKRudV003kJ6hKrW79GPSsX2H0rNcU
lPxuA8IHSnC4P64hYHtmesF23iy9Msv3STbbb2HxlXH9u+vV3OaiqD6j2TDi5P71F8WRB5SqFy09
iXL5xN8GC1Tlg27kra4W9T4ucy0bIoB3l9tjTvLwxZhow0iYKQQe0aNEQMHxmlzzdjwQ9FuQe9Cy
yhBlif2GqKY9CpZHEcHg4GCYlFror/GjmYehqyBePnaZGPNKW1H7rv5TpZsKvok+qC69nF0M4NZU
zVUEPGHzz/tiDRUgsgUIAooQDwvWdqRZ4D2sLcc0CmE8SMo+RNSJLeFAOzE/xs2NVEOtVwK/PN6M
m/kNn6RmAZC/cwaM3RgVdaUNao8DDwsGpO02Xd57FCR4lke7XJ5jYoWuYdIUGPwtdVtiFXWmILhA
5VmxFiPrm0No3CVUcWHC9BWoCIRk/jXOv9P0q/CkTOUI7nYIlM+JyXTA7PunQQ/rNOaG+1dCUrSo
0fmhDNS6eWkQlDaWuxZRazoRKPMmLldV1FAX6Ils5bcjZ/DcUI+0lYgFShpNgo5Ylaa/F8S8K1dv
1XQhk8LJhSBwM3+D9r0I6n+qXQpQ5SrXgotSsKXK7l4/0BqbhC6Wc66wvFQsYDVvzKJ5o8AwycPh
+lm09dnuKBIEIEZeno9iXl74sU58ULhG8dHABGeEMF5ops+XeS7IyA3gQinBv5WsjH4jC//9dIMk
H4eHPSs6TJi3fZ6J+6QGCxsMgPy0JAgWTA26QsywIY9PBvq4FdcuxqYx8lh/kLd98cui8a7XPnPI
VIMo76QjNs/5Ooydc3Gj1EpkrXdhIaQcsxMv5S9NWxEduOOp2AbNEDC9cNSIMT3LJkAFTY2mIeGL
8XveAZ1GMuQzXBlq3q40Iw2y/lUYoCwU1CbkOys1tI6SHb7HOhsX55/9o3iYN5q8ArnPR+oEzL39
8TEbSy7OXSm/ukktztK7LZkAOe1iDUdNDnOSOEA81T8oMpEKFMOzjFwsUCXcxIul5N3X+7bz1OtH
nWATNcBadCp24dUg1M/I4A6CvWNOlI+EtnvV/c9nzL8Lqq6v2BaaTpUqEvWUbUSCtRYX0y+1xPDH
O9pt9nQ2PiVaaE9dDD3njy1yPLMwZsNbd1Nd84A+idzIc5ItsgqCGKsc8T5cFVzs1L8vDvnGq8wL
0cYLz3ny4hn47ckO/WP+5dxquTVeylEHYDBlBa3a8vTqlGvR2lnU1k0WPpmoAz72Awi8Rci3NAMJ
9oPAZJKGBvFGmC6XEen7jIUx4B770GYsevhacxBpvY+wxyGVUf79rUyjAHkd4P6zH9+jWjuJtiIL
4T485kPQziK7iiM7i9sqc7pozqGLuzv+k8Dto+Qu+MqbJwTbZQk638IFIHZeWzQX7iCL9Zdf7+Fm
VY8eIFqShMCpJnFrXieRGuXKV/wLGg4IGI3G4lY1BprySS3L+TSJ3YXRTvjddR58arZ+HHXxJrxA
UmX6CA3fpu6lifYQcN17KjJ7or29K3Cdma91qr06nOEFIRvD3aqwR2yoh+sPnCTRO104MKeNjift
MR6VOF7HVuOmJUei4ZdFSPQYKgrxUX5P510Oj9R3Q/hMKAJvM28KrF6ESGSDMPRzyFFgr03OFA0k
JK7VGwYK81NKzEMkyl89BWCNR/MCMo5h0PJkg8G/p0fyX2/r7DdIJKzsJL6HtkVpXYWmmvLI5GZc
yfX3kDmlyfDDg4m02I1RSfFFhbxO3ryUuaR/DeFy/hMDtFTICZy2vvR7zDxqDORj5PxKyua9Hcud
KFdRkYHMbx3H1oOLsBE9ohpwDJozkCNz1tDXZiVeqIzMh9X21kKaxQA9Bin+iApM97NFNURpbeNg
ftJ2eeB2q2Mqk9xJJyccE10RgQOrBM/hj3p+AsEW6JlVaCKebPHdBmR03+rDGmniseZa0CxV2p+P
dzgL4ChN7819Axoj1+afhi6OzHp6ZP5oG0USKkN0M19a5DK5oyKfG7AAHfjQdKmHdqOZ5aL9Ep9w
G7De64VymxeSRSNxjdAEUv8e4lMeJsootOJ/LMjcGbKJDhEWWGhfs2nQIfOyFPjACsdl5pYVUkKR
aXg07r/TBgL3XQcrNf6YBwbwUxmYcmr+YcNBYwccpSTjnZwouzfgkSyfmg4cNzT6wW4C/cyWBZKV
nTskmmMP3/keBQXj5TFP3NFm7dw6Z0kMcDu7Poh0itcCjCdAm6P2t0t4wWVHeAI9FUbuyFHPjUsf
G8uZzarJ2zq/JeCTER7mRRKEr3mqIPVbijTQ59zTC2RKIQ1rMw3dmjDA/bp4oCmmWzyJ7x//JQ6I
HMriH+HrAIZcXr9svRXuMNSJmbDiWvtk9h44rl0ortVqWIy0k3WGSrqXaMmDdV1X56vG6cbPoEJL
L8qHN+zTLmrwJUNmHwG/Yv1ZsjdISR69/9oSz6mZl1Bm0oKamQ4CG6uegoBFRGh/O3JShrMc4iWu
Xo7APAe37n+IpZLbmEWnXkLHgjZjIXHRVIBqzdDaKEJENtCGSV389SpOiF35+fa77E3Sl8ks5eOT
Mde+qk9d6qcxulgZrU0p7NGXuHpVlylVMqVEEaGiYckoPJuSkLu2vRstai9TZp4LpQcwnmzB6Cw0
90fsyeTgUHCauk2ZlGLzruUUoiF1lhAG+G3aOsIH1V6VHTkvdKVEaAcirqwV1aIw/Fj46Kv6j+VY
WeLHMDkYFQ7aaA8Jtemt4C6IJ6usWBZuhcsvhXWtethPQL1fJw15qt80KZbONk1otJS085owvI9z
DWTRAexsKFhiE9qa5P3aHIMANxC/Jfz2qozMzHsgTmj7K593ajhF6rn3XaRMyYBUGnBKMpQXZkum
IV6d/507BZuuDlvrWJ12igXHYHMLPSGHYOU2BFM5kWmWvqsSNFR4DvvrcktMzQnIevJxl0BbdJw5
lb9kK9+m1h4Ko5hMtJHBKTbDdx/nLW4yF2pbeIoBRbDBRuPlrcB5ouD7qu2H3gbsSLx5wuxVL+XR
UgVNTlFJQsqpXSlXj4kWJRDZ0kyJBqJZXPyoDmM/a/9JAU1/gRrgTeOBq40p3R9ksE6bhJ0RTIR+
WpEolm4t03m4gQB0lUb1gogjajJnJtpQ0WH2qZ1P09I/Q4oDd0gh+nrF99H1ynAgjWA+XjeB1o5L
8B7Gba2h9zvPd+8JsZHVj/Uvm5EhMSIfJPZhl/TVdqrCt7c4h07kXypBejvDm+KrMIK2mNOtOePK
zTBAQolChxPptTg37f9A1rXDCOe7j/n1BWDRxaCh7xWmV5/U81Q28HWlq193nxzObyUlnb3icrom
5M77idwEmz0nXT6H1uJjnWy115Rl0doyn5uhvPpLgJ0FgECDa8Fte6v1CWttr2Ngi6vbchsd1U3X
39ZBIJy5UMacJ7LMoxnjVYtR2M+Fm/ivURPeWO3RvL2HJcg5pv/zZVvY3ZpcAZbf1aaDQwCnM5hV
KrOFeGyY6OuF0wFRtiYaYWhdvddEZindAlXVtAjzGMwevKUFBKrvFwcjbPakVxlLDsvtRaW++qA6
oXnwP1qIIgh05pm/qD3eLlUKiaaOaT8fJ8+hrFY3CzLCeAtYHBeRG1RNTa7MfCBM0gc3JKdkl0r+
kwz//rdqtwtaFvHBMdDSqEYE7YJF7Oa1iAefTvDJeYs0OrGEH5d82kwWWWZGDK+0zkK0Beac8RPO
mjycZhvk/UXxFrFKrS88qUJEsU9/avPxKt3rv7D6FkKNy+FOxskFGRigXvJlRmkumxKhjUnlkw/a
3riODnyshGO3Gj/rmrYeykmi7+hyBs0q6xfVQCuJvoT+oTl58/11RbVz5jq/LF0x0alSjc4cpy6n
gRv/7fotAJ+icc3SOs2l9VyFpJaqD3CEzgV4Er1Qjd87zx5v2yjHuA8Gkq50JJ0nnQtv/mJMeRDD
hNL4xeiCRU59ZOStWm2FC/A42QGotBbDHVUy2swWWkK+6RLWNEBX61VPq4tPoqQqUCKJFVmUeG2a
K5RkQlZ2QRs0DT7NEc2dL2BjQM3MIuBreSO0xn6XxGH1N/Svk6fWm/iRY0+oOxQsmUFN+7pIE2RV
gx7XsHh2mnTgkTD2FrKul0ExCj9wXSrR6EnadtTK0OGPtmFfBtMXJvtCOkJz3k9ypMn+qXKVI+KZ
O3+lGrhgeTWhabmUQDFaRs8McnqYIO4ePuwtL+qYIHKI5fzqWiiZ1yY13OCTvhw+xBgHQ4IfJmYf
wt+97BY8826tNMvh+1DajoDkwmLDYpCh99+eXbz2eMoVXQyun25f1bPr0/oC8NwB6KJjd7xhEj04
DT5YZgYv16fg1sUoaIEGm1f3y6nyEMh0NIAlBK/T5TtycUx9MXCmEu3CfjQK/+/CwhO1TMT5Jo84
GziCMFt+Z057hcUOoJaAtcvjcJwEoq5zDgJ/YSqUbi4EGd1Qo6YmAoaHUmc9bu7DbPrW5vToE+PH
7sgp0iFf+bSPySCwlEc1f1cQeLgJLfybrJGO/k3QZoVdCrvCPSd5d1esO0TGnVbkSmLpojK4BpsJ
K4D5YUvbLiZStlv+JHlDlZY+W6mtbkiKjmz72d/3YeCqgcjidXFaNEioNxkBx0puXVvZc5WOzwLG
+91WnuOcxCEfXYduDbKQ4YcDNsZU6cSIGvQEdY58Nd81Me9h+iY5nuOTMmyjUAliAHCO68SgtpBU
8PDpDiwZv7FCiqmMyBwwKHGY5Ges+gtsn7+uEcTgxUA0Jab2SxQ0cBZ3JbNi9hmKrVzNIvXyQ8PU
ZhlVE1nBnLq80scbboOy2f6gKKLpU5FteTMCF0aMfuHmj5DfwdFEZxekcn2czFS+HwyL9Aya9zNd
3ICstxZoIVJ9yZxTmjEj9TDNzuzrlEDUM8j1JEf6gf4cZ2zWsMUhPRSUzoBoYG+CkReHs7OsaNH5
qC1BKJkLa8HIuAyysOugHByYihip13W2rtX7/il7HTs8wWWt3wbv3RY1dPtRAHj7qCotop/EiDd/
t4Ur5GJOrGcRniLj56nuWIhPLWa2et+Ti5DkxASQeKmqC0jtH0p6E906F4/c0FEi/J3GwTk7RE7+
JPkybtLriz0y/2mRVaNHZhkGIj7X1mJOGoOR7RbIn598f0YY8rgP8WZe10w5pOam1AmsTClbnZvH
cj1HOJrcLNsoZhEdfHY4M5W7lS9lixGuj1CBa1En4BH1cttWbX9zHgzyeGz62eDKmeG/HUGRB7Y6
BQ3/kloV+PbcXGogPOpfpkRTJxl+i4K3T9fCXbmCz4/avHl+LPurrpmwjkjdKjsdk2pH6i8AHxkY
q0gKSxYHqXJWRnmILQVY2fjqWOweTrjdX5IvhhAT0505ErNldmgYLf1TvNIj5KLPCeGA21JkAEgq
CRjamtKs8dfQrvcf0nBL2v8KabvUumV6bWVNtv48U1vKcr9A2U1a2BaUPWNOJSZIwoohq4bJbslE
/43oe64r28YSvbicdlBowUlyM0f35yfc6X8Rj8mDJ9BavJu+CU6tTqpIvtQ0GVsNoWD6GY7Ji6st
3XCFIW/khHHNmbI2hK/97GPbtVuIDGXuaLRV6ZVPZgZQQs0k20ygmf2fs+16ySBmj197UDLfgXAW
MTTdIOVTmM70N0UttdTwGhgOUjwjnhHQ2t6KZSqTyhgcMqB5QVwVClYtEO/wPrQiu3FEt24VSvF0
i5/Awyn5ExiSowIRPfDgv44tQ4tOR04/77aL3NoFqo+9KOspNIyyHQLxTaa2l1otbXoztGdV2S4b
dGquFVnZ3l0WUTACyQHV6KHk5pDi+HAtPbvJA4jtWJu6Vb5bm7eO5z9CTcIscsqPCs6eY1SKpnYM
7c6aLKiNJTOPh7TNLwxf9LyV60G/75WBnrIORbjEYmtCxTFEbOSzEfFLvUxyivvhg1rnbFvf0s2J
gklf4gTyvFT8/8GkeoGOtPwu2gjnG1GDjzJZXiIyr/C5lChMeVq9oZfINpmaN4CHVJnwjrvsQx/4
g/T654RdTazbpW5R86fxUrim8XYbotI250NhcsxIcgVDruTxrrr+NN94+9o68LKvqGet/EnGARcH
qFSgpdyaHiS5MdbUJ3YIm6/HhJ4MUib/AsIlu/v4Pg/50i5/boO1LFXb9oxv0gaSeYT/Lwy0i5Yw
YE8w6a97r3DY6vCbz6CTau4xFAXGl3ZcvzrQZYmsWLZxQw8CNFHttVYoxuxHFhJVvhtXmPLv5ag5
RA8PI/GWdu9t7J/fn9qZVyhgZnfYq16fBq2MoQanllMDfs+QqZUshA11cHXntoqHYYCwbvK+D1K6
UcA59gogb7lcEV2dbtwan2RT1ZHQjOOI6rQZa9aCd3p6YbO2DGFKT6+CLVz3sj+nGT+1B3s0/gdN
QLpNRfG7JMm16LXARcRuRxJOIO70PbLiGU2bDCKrJw3AOmoZxKPjgg/SDalLxEBtGo3Li8eC9jU1
MKNdej7owZGEyvFfdd7xxm9g+jSi7Ctcd03xULhs+ELlOxsYYpbhwk0bJfxjFFN7MgadFo1uK/C2
8tHeF+2oS8ed/7Bv/Ya7qkly2dHYxSz+hy0FUKPPIGWmAyhkNX1MHHPChSySC/NS7RGyt6gOmgyu
LQpDqc6Zll8xb/Ki5Tprs+DDYgti4Iv3p4eH21reWaezrx6b8hiT0bVUcSf73FdvUowAuHiPoE6M
6ydEL/ODaxyN+FEUoLaoU7tW/hwwjx3BcOFIBbMVBjacfXmFpCQHdH2zsnlNE7DQDMQvWSVljegq
fEovOyQny9CeS5P6/sZAtWwFz/AkvQu2hpObv0KkeoRkU3naHIqb2vCUmPYA9l2BOxMUgJw4uNeV
rNf2rW7nkBLOFTBI1335ShjBGj4ptgJuslKNg0fkn8+kH2zgzp4y8yR/3+vtrZeA0pM61TiUQSFW
x8tpEM8HKSm+bzhyC+nJabLI4dnSxL2P+1vmNpAQo5DLFh9hU4dgXEpyK2P4eGAHwtSH4fZB/C8X
ZvRCDIQVAejG5QCYMEyOOIzxQ/sHUVRKSC32d1hxv3aaG+5Pe8LVOBoZuuS6OooacqUeHDn9tkyy
Mx1JEAECb9pLIZnhIgKwQGrK6C71emin7i5/gwCR6tDNgx0qC2ZQqhoDi0VC2Hrd4ic1AfOUoxrR
fe0kJtLG1LfVTSjJumBy4r1FUm/PRkdxjxVrPzt9yxtagGTTztv50csSadhtpnhF8QUWpwl9Z/7N
VZf7RvTfeWcVSs6h/S303uZBd1FD9ldsJWojPqlAwS7KnqHywkObp+J89BdPU9bGotGW6cH16QQe
CyxfyFMv5ArjcRso2QjVpFEZ3olPJ7Q+HLwGFnPt/wQfWpvh6MK5Zt19qq+KghuwL+csi/WNAEvm
DR2/heORB908DT7HGISqRCawSKCOBkdxjkhO4LvyvTrn28+cB/IfQeeVSSlo/FZd+VE4oF+cDuKG
4aCRD172UHRVtnlDiYukruPtP/c2rm/DdKxWcaJZPMjvBjeGFmyHIVuKLZl3ufZt1+yPkxW2pKfc
OD2mrBsZdKYduy/Fh/gInS9YxtTy7clzTzhTfbjQkIvfsGvThx3K0mTbs0V4UY9v7MaLf2OJsiUW
fl6yeGz78GNdnThyBX06sG6IkZ6nsnAvHYRd7IXAiMEJMdX+hIp/VL/nto1zunNaHsKlB9EYYxLP
/ne9LmyrKK8rxNkNL0euDXW+u43kMhpg+gIYWmBiS9oUaATIBlMbWlID1LmdNJVZfnHrmdquFROA
MfJrn9UnAy9IR8hgzhXFr5aNY+fr1n/3mgJIXGdjokCcK4qE1e6uIuPZDPy44Ql8Pk2JYAjabSwO
3f8wmVF+ubietSUcv3Tterk2Ghf5iDlvsZEyovFNTZpr7iZBMem7lCrU0ohs3MTtwq+5Z5Gw7P0y
FjncDKzhAQ6BiSbsmbmAy4+GEDIDspotnDwV2NhZneHf4wRXHsc8AW8SkjaqDabMA3aN3P4RD+Zu
Bl3BciRmPKTRlOhSoQDcpjWZ61okGSdkdSUg6E2NplCeNgXtpjalk0Jl3DAAJa8/UlTXX1Pfsy2H
AKVhrSJCnCM2EUOgI6CQL8A1cMjIM5Zh6DXXNuNOGaXm2ivWwxrcxy48lk5hs8snXKkFyV1T3gxA
Mh7O4r8oneB3U/bJiobUo/wrvpuZqWC8MJ1TgL79coDd1LuReZVJ7dbXqhwcQV/839DyelChiVgc
X8wUKKw5KO7pZVIIi9+YNxhqYf0iWst3zAKzppMkCD9aR3Ra8doAiG7Vppya/zV0o4CBCK53PAdD
O2ytrd582JzXSjyVdxmvptR+ThJqAu1PgXIkBexB9x+tJYRnzKRz7KHFPD8vNBoxEyx30l9mzXe9
UnnAt9PxIauvfiVbVD1QB83SXduTZFhWQwxoG2Pu0BaQknrogQnb0lUso+fk0uG84eip9ZS3YRuZ
A+eQlISbRFXtLXiN69DbkJkUkGZV+JkfCNHTEBF0iVsQXPOk139qDTh36uoSYVb8eOj2Ox1tV7Iy
IHQ00bV6a/CjsVc6ia87ky2bpSWdMVitIAX9dhVuKwmfsSnonBiLNwBG1Z65mIS0kP3/Trvj74Gh
CmddFvWzttFYgTWT8v69txwTonVWLjH2mKIkmZIC69IfEz8LAX2nOdGW4JJRq5cafGL957Gy0Cfz
gTMpuV1YXsc+SZ66TYB2fYwFVtMwgMWb5cAbzWa+htwqngyJEWGdfMI7g0B50xT7SpGmkF9lYP8W
gFbs1vJFcHqKOR6uEsMIqTfKFlSZHZFQvOGVi1HDhPsq89raZHJXD2oeOhjJ57yuNHStbMNl9BVj
TewaxUouOLSQPkNprS0PHBUVG2upW4aEeqleMV3PrTYxquwUj9pLFcBN/eDCeb/BLRiEi6TYDCyT
zJpOzWCeVPOYAS161hVko5M4j5g6sIpmeuJLxu2ZFkEjjdR0EQY001YnR/ZaaFIc/uaWXcNpourk
t51ln/T9cMpx/WOHbBv43IrpC0k1ZSyaFwwDfpjvn6GQhMeWo/o8rtUB61EdLnhg6Vdoz2CupmyF
x8Sd17s6FPHXn3VgGXtNZOZP2A8COqjt3Z3KVrYpaP5lns2ua3sKqFEW4QIxsvzpxk6CPXXPzHkP
SpxUOcYFQc9lsWtlAk1GPxt45HtyES3wU6bVFctAUlif0kFTVvfUVrHYPOzC10ZBhFQgTmYMTGlp
Nd5ocjHOc2aTfOJXpFNjiwG/k1ZJyluyngNp21ZdEIS/pLK4lHvwOXLk8KNaJlzXYtcEEYcFYVVW
kjkjQkIHXyfgMBECGgnbVPNCLYAN71EPBsslB5GtOy9I0vJiu4FlHFK0M/50b66WKK6p7P+J1S4N
MH2RDDf9KqQGjheqK0CVUO87hThUx3IhJEZ1y4GL7/hVUwn7loO/RTaz/g55C/pKcDWJSElPPiHb
ntHa5pf+3tB7bCLQRp69zDTk0DrgoLv8xXAgTBenNZmjlNSz/IT8FJ2/Yy8f+xur5ogruEjttTqu
9Kd9FE/W2Kh/9Ieg81EwC1vweqkkDvuwhr/y4+fLOLZOdiqos7H3MuPj3eo4VDdMeeic+nWLaSfD
SaU914YqaE1fR96i94b2at5Xb1BYU/YSaEaac6prulrx7n7990TnvsMTlpPBabC4HuPaGUSpNsDl
dbIcDCdsfKsENdbJE+LN/XZobtfOYNGyu2c9BOpIeTSZSm5SQg+JRwH1XYyMsdDEyk5cmOaYf73M
ptYZvMcFJObs0dSJ3s77jrgw/7SFhjaS+mV33dNcfJ4/xIUKo0XqKIE3hhYlt2mv+6zkby7T2Z6l
NjVn5pc3e+tN5Gy5yqdzPMpLt2b8/vrSU69kd/kXeHSJMAPQ1kwfdC9eKoTVqGD3IYLiCbFlduf6
dYmprFJ0Lxawka+X10dA7E8wyNpmj8ic+H2oZHRozrm9NiOntV9aSFum5GuA9eMUXX8bbppkO1Z2
l5rXv2pIG2S+WUkgt2y9O6pJakaw7MN7jAmNIt1hmk5Ax+4xhiuY0Sc+dBPOuLmibBtd7tKAHN3Y
YEuapSSfSrciIa55e49vIF9odvLcd0LzKKdanR4aP9LurAfx5cPhkqxOnvSGG3E1yvUG4PmwkUQO
+3ZTEZtVcocLDMZHau9z3yN2+bc4MnAY3MfaRf+uLvWY+uis6pBMlCncCH95E+Q55+z93sIRLo/W
jVDeaN1wgb6S3EYfBIMfxcUTXIsnttsMXI8jQ/5qbHunsOCqqs3tTP5+Z8lsHi9nMkbcQNfQYADI
1dy6RX6Tqm5ISon+vzFpikF/LNCz/ewDTEkpzJU+4tqkfOjq/TK9eKSGMu9N/ZNUsVMYr0Wj37YU
81qXEqqHwhiL1b+0AqS+4IgmFmxu+BNMZG14bgVPTQX2wjgyTGhN1a58VUs00LIUgazpdeAMlIc1
Qeb3Tg9/F1PMocf4pFy9Jkai8IF5GJDoU+SxW7U48kqTOi9I6Yepvtmx3I6EwxwgJ/e1TDZgYzcD
cvfkkfxFf2NnXXrMp1Wbhcw2J9AV7jBfCKg08UDxsFn397c/R0/wL7Bi1WeH82tvv3W9rw54mkhw
Muo3Lz1JwWkyKf6yyyRtYqVfssPhls7PjxA3mT8CgNx5s/rMOSQ3gUtGBLoYuELGHCOQ+8NG9HLj
Wq4ASnfE1XAQ22CFjyISkQbOK0dP7+So3N4HYvrarCaXqLUl1dmUR8VSMd0TeKQF8VB3XEKpHNky
BsX6iUjlUjJ+RO4yWIZ5Sa7tNSK2wQI9UdE3kJ5wc0+VlXTzHzghLv4IkzlRiVpRnonV+kSenPzX
Mem9HKnzIDr4ugxICO5L9I/F7FT+OHzioLZDmtaR7fxmznq0B/UtFiOiD0qyV8KoMDWPB5Bh4PIn
WLP8MPiLjPYRHuSE8w91xK0SObDcYhO+l59fjN4/ne/FM32pWe36/JYn4gXJQvaORdWpsw8Gc+0f
rzv6WRBwvTtNakhstdIv1DqoLcoHRZjpMPDC1aR5ZR2jZfuhpQnl4hXvOpcXP4w6m8DRnkUxKS6e
e2zToY3dq256yYETTjf8OGsmxQC5IfUZmhj0+XhY1VLvZtCHzJ+7xpDV66TOTSOCtsAB/Rikus0J
9df8rZ4NeLNQkK1wLAlKJMqWlckuHYdAbcWKMZ1xeRKlDQ1BaZDLuycO38dpLxo2hkkGzdLsJaiS
2aufemWhjZFv/qBW/qwI2GM7prN5ZsryHu7EPx9JcywfxwZ0NdXBcwy504zxmiz90lll80N1cvhc
VfQ8nARRyiICsJuYk1gb8cdgZlz2lpeE8W/9Q2ELSX1nQolWt/+LQqOiiITMNJ6WLxiFZAaWrEwT
IKA/vFHGLF5xx1XuX1o9tg2NXwQNDlUauXFNhS6y3jxs8UKiwy7KqcZhF84/VuRJ339P/MHsLjVG
QImmzroD571DK+RL5e8Q2UCsMNgytDaYLLfFv5rGDjfLkOcnTXQjA2mvWrdSkUYhu7Enc3+/IHz+
yyY67eOxoD4a5YUujXZxj9wSU0KgIgAP97whPG3tAUkPbs4dM2Kws+kZwYwTS7p/C8NQoL8DtZM2
E6CVrXVfEdX1ZuBE/To5LJ43glkr40m9vzQmFZB3p6McKUpQK1bamYsVX7msSRoYMxtpf9e8mXZb
SoKoUfDJojxED5ia+hbAfozzcLvrPi14CdQqAanAZ2W2nJWJ5vU3NyPkKnwaHjd9Fu8fuuzgTq3w
R/9S3mmTkdBi44uyIya0J3edXoJg2bruFKeS1dYvtyxlM8J0obrAUl3xZeA8/Era/oJd1J5tKwbf
gmeiCQ4bLgRf9VX2QEAXYevXB8WpfMbtZc6GIB9VyvHUxp1okH7bYk/lpNr0ZCxP59tAOvnFNFIQ
xJfcRRmJHRE7qxA6YjimVLt59ffNrHHxYegOv+GeTEpBpLujHOfwrQo0Ph3W84d1K89RyLVgd8fs
iuSfP5/nMmh9ooYdse6ApXXuODRBCWau0i+CDwTmrW83O0pxpoqHgzN8MLBwLgQS9qcHdv1e6Mtn
ARmuD/7/Ah/+iqJP6GX8P4j/sE/iX/2q/zU2p3oqqqMDzUqjBrw1mw/+dZw/cOaIhvvRJhEouUW6
3xv50SGDNbbyuDzh+5vt/S6rLSs+zVZTddzwSMSQWixPuWXiO2J7qf1EaLDsQUlSi5Kk9GrdsedG
Ck1jYrYm2Hc1r7pQWNqZY7t2vggo4+FFJzVAv8UnH0R5A3Evc6pNjVKbtFtD4r73X0kVNKOemmy7
+GgBqnfysON4KpkuPmrkE1i9NeaZbnkcuuOmgBdhjSFmVeyTEX0jZLElHDgBGw3NtndnnMPUuigh
OWLMn4cpY5zTUzV50rgU6Zyql5HJ/Ss8pGoRkXO1Fpt0UxHXRjGM/CCbzMBWvKrphBWryBP7uKYQ
t8z5qa6cEIFzl+gAxSksvofFp0W5aW87hUWpAhJp3+onU1fi/Lw1g76KQzMLjv35bO/PoULh+2Pi
ms8oEywBXgLa2UGp99yyYLpg7ugP2VOcIk6YlDBeyd8Vn19nbT3aUsRztJGWDa7hrzMNHv/5qNkS
LkhBfT6echyGU9NqcTROKyaqeEGe+nySm7c8l7PgC3OJXy0c3jO77YlXezka5hWGoTkvSrk2mns+
pqfGJunrD3biE2IUM2PgauqWo08jrK7AEd3L/RrzyLvzmMS9yXsRXfHqoQ+BAB1tcru1qadc7YXQ
C9JLB8CVEYVfqrHRwxbRRnErRmr0AgM99YnAWzGTaSvbOi2+qqLH1t67zCBXusnJ0JPMYjKS0pb/
J8VY0g+wnRPKQ75adOeOyik+XZHzCPKRmjYlJA67qjRk7qaPXYlLx4lDdL660mcZUc4Le2L78Iyz
Qf+1MckafVk6F6J5gjeNbzbiUl+by7S7K16Q96SpIL8b2GqUphwag3BB2iIi2EtF3bWpJ4YBzAlt
IXbzqoqc2fhNbP2fZC1DWYvv3ywmljOHUW5Cso2d2IDekPZqnswtp9Y6kOAVkEbg3Mxm11imaG8T
ZcXNcqGmD+y+N5JPOGbWJlmx4uqL/yp1Op2Kl9QrX90NeoOwPVzOgW1g3QjOgKOALqKdAFvR18Cr
RnOv1Y00ONjS5oPyY5mkMcu7wffQYavrctgj4yqWys03Znd37KHpFlsIQvHXzbvBlZtMw+TwiKsd
+9tfZVFId4TX7N50ubljPRGAeqLfAZhIWAw/B2cBTqKdIclZlJvzb7SAEMH0xu59SkY22uCVIYZy
gcZA7ZPzLZLUBNqWj4jbExeCe8jFnfhOxTzuW2SXykoABTf8XqKmOx9JPzlS+P0+r3V1pIErh9bP
TgGF+i9dsTeNv788aWb1zxjbDxFAArJep526u313hr8SSxckJniar1QiCq96i1mKib/VTC2R7pHZ
2LLw7YScr5bB4zaZF5y43W16yVjGlT3EVgM5SIkSjKqxxIIEncN7q8Ddy1Kh7qOMgJbvRTN6eknE
tcwlvcLo5hF0Mhvz4ihTD4Gh2oUmVg3h6J7964s+yBysFFYeN1IlhbtUUSmQHuovUf6QMwR/o2fA
bZNvg/iCycN4FaImAgPbJgGL8BPK3mf/UuPHWjMkcyt0m1R70RMp8lglGNHszlIQpPZ8xGVM0rqU
QGgr6qUz6jVNWASNgT83dK8MQ7pCxqDvTDNskyVQd6XPwsFNR5067hLP+Mc0AUZfX0Ur1DW4z4HB
CugOeMwCvefuovNvVIcqa9cJydaGhkVi8lNlGi1MN4TJnHQ9ketACo258o0m4zPsyMOZSRX9iLVz
KT4Lt7FYlf5miQotn4E/+MRbgLT61CcgSW9+0xHqw8mI/Rp3ygG+Xqf6gY6FOQr1fepbOsgDVaU/
j2gL5/IrUKkenQNBinEKxDs7DNbcQAZPhoPoCj/WSoRL5t5Hul+Xf8krSwS9skCaZM/QvG+o2Ned
7e27RsAUZlj6fk6xQx/JWUpGImf1m4lYQg0n3Hqa8K7fU+GQgdD/4jHmZrwDIjl8tHzAaWKDdVHi
IL1zKP6tYr7Wxs1m/ndwy/HhGr6qy4zwpv5HQtZg2kv03iNWjesjMYj4nRo40dx2dNsJdyAJUUhP
z62bj+aCPBYbGknbVu0idDG4NtvfxF0UkPPodImQuIfAt9U3H+1rszW3VwcCcyaK7N5RU3HQVeHj
P+T62bh8D4DRowZethpa/gFogX9u0xq7wDSDjl/4ewj4sTmptifyqwarwxlL8E2gT3howJX5Bwm3
4GMdrSKw0rIT2AcfFSwHKK6IIEjPXEemY+o9pjzKh+Ln9ZfjRpAHKDctwiYY8l1ne1gU70y3Ob23
iix9CkQGXEM5bZidFYnCNk9Izt8HVSz6Nf7Bhu2OxbwiQrBRc32gsXlYcdIUF01gjPr63Wi9Xp1P
hg7JbK+MjEFKYUqS5lF7iJzy1suEBnH4aH6zgUjIP3RwhQoYbGgjFKNKAX8MS98jNTfeMs30AmKj
/TaZXs/cCqNAh69vvpw5PYMTUsRvChuUAaWWGv5E0qj6hx2tIUdciwxDdHTjYBrI6f40KZSe5NPc
rErmnrAh2LmErvOlTl18UVwCd7ERNy57ObNkWR/dqqe6VPgeTybyULRSc0klU40BQ7dXZXYETsp0
IDWywC1qb/9Ci374xrFwrsYJNZyISVb4LICLP41X4gjZCCFf2Qh1KVUo0cJmHjblF1polstPrgsi
jRulzr9tBCwMy0nAKx8loEXdMQvst4tgVK6DcQbkgfVZVLHUbGOo6t3OoLcZtJQLhCdzfR4/6xet
4IGXI/0McGtmTsAc6EWwFSpuMXJdRmI8veXBnQywtwSAEuTIL3XRMB7vTNAocCTlINgVCEyKCrBA
m+JXTuifWINV7k5L3HqCbxJ2Kq8yc3OH7y+TQpSLs9020J8GkxxrUzCEVDB3Qn5XNMUDH0AamvBc
6Bnz9GqE/9+eyb2EQBYyInWSvEVJ2MGFbHXNeeSPyKz8Nl/MsYS/xY933vwpboa6YuqQYHwo2gNr
j9tHjF9G63BQ6H+vh378D64colHi3LlA5FgBGpbbhiJ5vcVo4CLJO218tcwUmAYHX0mS2PVW9Rbs
jiCL9FlXOKPsHKeGz2kyvhjdDfMzMaFwChFXITvZrlYv1YnFPagIXjnhM+vkLVDmgSqI9iiWegVK
k1Ln4/GkGzGMXiKnv+sSG1KmnVMEpYoBTujQnVbkFi3JCS5026N5Nf4h0gB3k1342t3jaGW1o5qf
kk+8FxSJshWIMqRlP56dHGLOlShNUkz5x30JEQ1apMk9Fe+ScKQxHkqga2CbUDipPyRxJtU/Yrr4
21+Lf1ouKGY/6bolajNHZfIVs4JiC99yD7/GD7s/t2nR02yxuGDrUCEhigjw8DcpyOiQX6/nn+Bo
IicXOMfskPWJNPXDGpNCq7WHA0z60xuOp5B63xT2mr3Edbvys+9K82J4DC7DyD+gL6dk+vK2OIyv
w9l8r1nNsoT94eeOzRQyid+0FC+CgYPhd+dC69/i4l3YoJHUpd6/vhonRQMqC2HmprIAFZq5CEfQ
jzn9ZA/IfS36JuGhqsE4YCDdZsrgIEEytaNi5iFnOWAPit3Qv8XTXLbdfpjdDLwQYmGYipG3P4I2
15MdMFSp50cD8Q18y/FsJxYb2yZYvOpBQzbM084dGBkU92t/TGlJTcROCcBMD/Rr+BHz6Ic/X2WY
hhHKNwvF0ucKtRl916Lx6WBk/l5XyM+ryKG4Jpf1MUu890xp8LLBOT+d1hbQn3G280zVJQ8oPXSe
n5sE/CaUIf1iKMC6yANGDx7lh/yvVXAZUcK+0inr5W7AY0HdPEfYVYzKARRuOqeXJa8BJyx61Trx
lHnrn9ZZfWF17QOw5TV0vmCk0ilDAJ3HspbDrPoFEFIfQc9f5gmgWwxonXk0R7ZPUaazXQJj70nH
NF4PJxqHQoauYa4ZOSjklyoh9UAq5EDFqrj0YM/yvI33MzwX9SaD3tW8nfiFJlTG8c71RUMmtvkT
yYY9REQ9JOukZ0tK1z8XtMJiil5XR0/l4+up30zYoxJFxXh2cTaAJQutLXy4V/0ZYWir+vdcMZis
VBULpIxnQ/pJ+G+aHkvAL0n/vlALN7yGo2/JIt+6o3Hm34JnhBKouYuP1rfu1AQHTMaAjfVUoDFp
2/ommEc/Rvp51b7ngZZe8aWpd5k3j7vkY85sK8B3zf+lFZA+Gw9zDoaPMf3hg7qISfuFts8LAsLV
ZAoDU8nmMbuZtMO4kBb/8ohRGhCfXac5xbr6/zLeWcqE5OP7DXxop1e+75F1p7BunKGl35fmOKqJ
EechJ3DCdBXjRVWD5kqewV7TNQBe3ALfPnu8cgQ9b5tyJI1tVP9py3TEBI/m7/nCXvTS2i3JR/KD
x7XoEz161VwXYI2Ry8Qb/FB5pU199IopxgL2dOhPBHHnSYiIzUZ+Euhe8HoGQUpqo4EnzJ2Z/DOx
EmXcMSj91nZzNuymj3C7SfU/vqVyvEpmgM518gtUVM76tzhhvOE66mK5mDu3aZ4K1k3yI5HambZW
EDurzLZMD+GyHCfNWgXqU4InAeU/EHuHqA7bMSYVou+Ne7EepJAuyJMJIUqiIkXwDCxec7M5Q+E1
9IBkX7UFPYJrGk90vWSOQwcJWY1I3cpgFggARgD//0C5CYuew0C9Lj7EagYCZcrl8gohFCYnKEPK
KeWRLp+dOoq+IWa8OtQZPvYfICWYCu+WoXmdSgR0KCOO5/ZT3pwFQfzUX4gcfLZsYj9GCk5RnIEZ
s/xcHTnLFB4aZWkzQdq9+uTJ2Nr0kNExsEg5Aih/RUaHGJA5O7evazyNCK+1/pLff5oldekrCTuH
sDqwINQoV/AF+dmjEDsxL69ZkRCyJzET9KMwlaHXNHoYzIIZTGrL7FuwgYrCrn94BJHs+J8tA/AI
ywP5fBwxmmZ++wFfNnqSlBZj3EdMWO+KNSThCoscSdKjRmejZwrS7Lrib3cG2QMSW67ei/BmVk4d
iJeg1Hm3S9HC5sANuXWBNMDCMHV2ouCaPvbk+y8XS6IzMDB7yzNsK18B2vd2nR1r1qRp84MoWIp0
2wbdNUl+O9sH4vdMs8Jc/KK1PEjJJkqfwNOfGhCo9AwJ7OrmHnybUNUhKPieS5qYAsk5GOm0YgJE
3IQqpzsWAoKzO+ZGVUInGgBo61ky6/pr9SevtjHkJ5Mtwh5hO7qvhekPH17KbNgjGTkjE5QxT4fk
7o6MzcsNiCjT0OztFAV4Vq4p5m4rUHv/INt7qmAKYgPF+9yRvygoFwvZEZaQ/GET2IZpoN7YrHBy
GxOV57zh2GdbPGG2Te6TVyqy9lP99hdAtSrTub0ycqnYVRSY6HNN6UVB3PVvYHq54KUP5MQqcA+W
XjWASG+Qh8JQmgXmkSI8/+Brp6UOLFtcaKXc1Om23gKoo7p+NK2b5MPY+nLdJLQ+kMbt7kcZAbPy
WDw53fjOqxs/t39pntZi5XGeaEPIVZPALmSrMogD83c2e7mbq9KAeWRPgqAYzG6cn+4ShZOb5Hym
z6fO5nUMob9jqFf0IqCczkVvn7qUm1HH7oPiECQ6EVd5K2r+TIU+ftaw7RySiuOZmmCknq6Grt0C
mOkSYmCGQQ1/ebzmWRQ6kb++0kMknntjtAcwXktxAcsRUru5YX3oDtfRQIqlGq8Gwcdv0JutX7E4
iivxVXN3CC1MwEDRws5xfl6dYP7BIICdt0rP1XSVYZve8tM83IBvedQU4y84eVmukgtplspZusQe
tt4UPAfP01k5y1/m0FwtSogO/vvHBXmVUqol10j3uA9KUiBKTYtvAqmvbUUsmj0YALhgcw/DMAXR
xJXxBHfQGYXLLossZTXtbas5WzKpcL0jkb0rW5TqiWuTDOayyVZ6Yxlc4gNawfCV4metf7kNX+Lh
K58U2+aVDPvrnnrie+RRBnYiHbnLmMr9Hiy+40Tsn1rLvkvP8k88/VSTPOgGDh41JkPpb7dopTUS
4wuRa6EHV0nnB10RNOPoPbfiQkcehYQON8G9D/pNW115OgQ3zigpHD4rAoWw3QsfL35DV9gtscJO
EPk3Ly0bieoNniZIRV1hD8XemO+5cs4k0jlw1aCXJZCrgKQUG6LUlPehF+uZRKDeccm2UNmz+eLb
SPqH1k8zUWh7ml++ef1MRPYL9kx6ookerZvQA9Mz7CUsnru1FPIMFRTlibgvVMhtmo7lCdwYa+FE
hSFoYi6yOz3Y+16ATlsHyHgo9U/fRXoA2drMVYb0mxdfr0cBZh17GCVo8yeBz9Z8PuTOYUdkJaWR
DcKSlV8S3SD9IMo0iAI+hgCCA4644QMzjBSEM+pt8ftjdYdv0Ce614585v0SzG6qugwypkG6X4z9
dU11Krjs4aOlOmncUxGDbvaok40EmakPRWs2zJpY/rzput+RZ+ShJsyfBmTQq5DR5NHD0S+fbIMW
r0KsphvPvnDjW0boojNMIZz1UHWaYdbVZt0rcwJMQgof25N+bXov99GE1lrHU+lA42V8pJVUWRdf
Hll5k1l01/MtI+0kDTRCbqNUZsxR/ScPG0HhN8hfKmrtJwhqYIVzNiDDhTUoo394vbIucxy8Iw/n
lepcx60TRGuxuNl46lz3UEZOQAxJKdkwxF/bdwTTRSBDj4ktXEjc1OLLghga9QTybZwR6iLBkUDv
+BthUGT4MqbKS8b9OENWjy+9p+2gFITnFUK8vpxtts95BgeF/IYK5XX+33TFSC8tx8rOykzKMB1p
nrLS83oaGVLCEWAXx3B1CWgYPtuFR5pR/DZSOKzZFz1fKzeyj50B3R4vNobctCUaHAdGxTReos8P
JL5GaGmJd7neZuCN7VJY9M+cakSM1KOTTSZEwqAYDoscHTlwJz53pdcRERITfzQ6nES441N92Jhh
8JRtHIBrgqyd/3fy92lVeK07Q9lFvylQFrd49lnUoNGIwT455tWnuDo2Zm9GD+rq3hDMLrayF35r
qm98rUclL8XbUYU6d90rNEk16Rpoo3qbgak22QV+hM0rbQjFmLQBtzrCTxSpCRDi6SA4TArjkPGI
KT8G0f7SN7Ax1XD2UA/SEt226MnKkGLy99qhUL9Imh2+IdjSj+1YHEClbkHllbZO41izBUlu013m
pQj6G2rWkiVWzQD6Pmn5i0cM+4tuPI0pxM+70Usaxw6wuBfVDnSWujfmp1UV1x6mS4xamTvGk8Rc
pESgEu7yjWumMKpOTYv0h7fSUJ5PDQQfbCPJMP9ppd0aAWdfcok0+pznznD3NEkP70tPClMvwyfA
vt3Rfk9egq3m56rSUaT3vBDxex3BVvjdATlT0qqzb3HIHP5gBwh2IRp8Zc3N5nGtp2afpi1uEc/A
S5Mj2Sci2oED/ENGV/dgOshzBPixbWdq+2KMkyQWQKk+oXU1BDSZh5i9mIYfJpXcTQZv+chcHeCD
WJbvCwIfsld2d9/wURzrG0/kmEgtNEQ/Hj/+WEC3kELKKEMDIx/KJ9SuFEY+zwFXkwz0Jd1tIEYB
SAq5mI5MKFQ57fdeKT+N/zTivKhp1PCVVDUarkxDPzEvxW50gmLM1WryccihsBP8Qu7kZLdoLXUJ
G4+nM2Cd0ufNOoKuCtWjVjEfLI2YXwCqw/5VP5c81rQj3gkem8Ypx+wDSd/DwS7SttKW36oNgL3E
jHmmAAvWxoJOGmtJhNXX71kSk6xCyxZ2PVQrLOKI0A8BnEu4ryQVak9qibsTFxGTQUWAiJXn2kH8
M3GUWIa0rWlc1OItz49xN8QN/t45Sb638dgOKc9PYJy/y9Gfi1Hio8jdXvySzz1JwSJieo5L1dxt
G0ZNctSi7F7baR1zf6Ksw6aI7lWY4Ms51gVznNNB6lOUTeRC7DsPIGRmRSS4GfX6Uh8Tvq4T5R+j
y5DcdMtSAjO8d4pbNDIYebKWIVcR32hTdZEm4PPQz0fFNE/JaoYnsHD1a1txktd+rOhZnZMm8zxH
0T56eV3MRSWr5k4ewkjXFQ/kGTjAEpuA/2B7I+lnz1cC/+GlPZA8G0q2v1PdgKWs1tMTbvKddsWd
19qaQYp54KVY8Z96BKxPX+qibxnK+L/Vw2AYSM7I95fb3pFLMFtToDOnEMwEEP/dMf1txiYu8fsu
CyruMiUvqW3yHgRV65Aqottsd8XtKMtbqJWdwMtkFl1iO7YTM0uXuCdFGfTiy5bib7BvjyPnmge8
VjpZZgKBYHm8ve0moiT+HHkJaUl743GsIb3keVjMlvZ+NmXIbrBKsWjhY1Wl858ISiIl9Yl0XrvV
GoYw7e3RhFE8C0QXi825/YsmBvzFLGyektokglB/nI9wm2xetnAq/82ds5iAzCROjLbolgRL1OKY
XlSNWhMS3PEYZjzRTSaKHZwy5nBaZC+Dkvpa+OSdlRqtWGtuYSJpA4WOG3uqxcT+eNjKdGtMSUOS
ZNCRAJ3LXeMyBQ38H+pv3EEyr/uc0k6Sfwm4YR/SmmzDjaaRQoq9dowH5kYpAenwBXo7ohkOAhXl
61AbXJgU7jnno8KIsQIawMmmC1QLz5riNiRjue+SlPKW7i+/Nn5fFQTOU/xABj1Lff+yQRI+gvXw
ZZpIG8OoowHmTnmQoDlQclZ16fAfMCZ6arGYP9xXPJe5YINUi9tqTBnXnodE5i0Bjsd8MsOlBIgs
2F2c97SzBMySjoba7twM5DcScePZ/GuR0TLG5qd3zcRp/uXG5qrm2caMhASf7VkTf+gnqMZDKBph
wc60HilhJdOQOBGcPzO0kKiil1CIS/TZCMxSCXsFnLaZH/2DDPVvHj1teLt2APsD0Xe0/OjIsg0r
0MlenZq1axzQQZjrWRSN3LqDaztYRziqaierX9+OotLPjRzuuQlIGEU1nf6SyqceI9W34SwIWcDO
0jCfFW9VFezpgdzfgx+LXobe2pHcg99vZGGG4KlRW40N78/boO4/bqJZjb3qf9Xjh2K8t/5aBC0p
j8RRTvR5Rjn9dOekFEPmn7kY+9E04wxzBgngJC2l2kmV1g1oE3hsxVebGi1Ac0/CWAhQx2M8+PkY
8ucxwlRmCDZgmYnIxvUjdv4WikK/zEpi4FXilbIjDu+KPD+Wp1H0AvSd0vCFBducExfMPKjQNEIX
FyObxwOdlEY7Or5wPIUi/PEjIChTfDqtMj1unFlAfbnyGJ7abMXf7MqlBE+9vheOWyam4mS9SbTb
UCEj4euikPzj/rtqphvK6PMocymUcJu5+gvjhIXtS7vcwwUfXRZYx1/IYVKzgEYMeQU6jokUXc/j
Jjke4nTOmgdikA5BKKAzylkb+ntbunMX0F4LBWZ8TT1hAPKyB0dhDiXvEVGYiW2LgqDpYpnMjShA
9Toax0634NcoUTVwXmlAKUVnmNTJptXPvsuz4Pdga5J/7JSafOrRX+mjKrGOHjE19hFDmySlTy4V
H15Nv1xsj+kxvXvFe/6mxsrBvU4ZLey5cuJJpcN/SmLsmSHrWqUQb/XdT/y5SqgdaH36CqT7ZXjy
DfC4cDnq0DLIzARpbV31et/T43+OIqp0MECrl1A9+056NoP7o4ba30gxtuQnf2VLNNt17cF7s+6P
i1LfWzNus4OT++IZgF1SE4UY/RrRQ+tpwb4oBMRL9LntS8of2b3BhCw1oWoJJX6KabMbWrlNPHzt
WW5QSU1BxourF56ye8b+HxYtv6CzEHXzZeecV6DvohDB68GJP0NOR0Y1YKsQv3NxfAMEbrOigYgm
8xc0eYP4ILhh5oiCyDjjiNM4nw5JNl/JpjkVFJCmmwlWvEai3yaj8/JLSEid3O+d4uIp28WaNi6B
A/i1Mj2QeK8znyaGvdrfLV5c8aXaLICaOTF3OH5kvMqjxeRk8WerumfGjSKs33o/EifoXsD5j2Uj
bqkAvTQAwBgg5cPv7aTaDIZ5ZEEnE2SgrJowsrO0w44nApEogqj3xBMzqXdSHspHndXrLUJJkHQO
QP5J4LRjNKgxGjXj0S/F0JtrGqHTsbZlWrkrNTEArInQ32wnnjfQ9+Wq3GpROcW2XMnW4Pt9b8vy
/AIn0H1vmVT4xs90UsP7en6jrQXu2LaAy0PJnmaA+6J8EeroPZFj8M5lpwY9MZJ/r5KBjYJJPUXk
TYNw8yRFbiB5/yeMFad7TLvKeQV+AXG9x56ek9yox32DPIHtxRc/VEbWDZGKmHaY9177PhimXLaR
eOTw+Gq9eL4Zs9VPI28ncQAsmr7F5+Aqc7+oonOs6J1Ay9rYTof1Sw39q6bOGcucAolG2aQkUsrl
yy0k1POj+08LEkLtJklWJVfdsS/SZbLFL6gioTe5lwljykMyRICCd7Xz8aIfB261iYGQknqOdj2K
OrToetHmPaB8A5YDCxN1fevN/sDRPJ3ASyTAMKa0ZGavrRAT8ydVj2w54ZZNrTUll6yr3WzLkxh5
IDEnBDuRPRQ/C7Er5oAJAc3zYKNU24/ofLkhRD19SgOA5rHBy29wGHn6TUuHoELH0iOGsh6+ugd9
EUzp049xvGjVx0s/hmJ3zb0PJQBIbh4rfX2flZ4RMdQsMw3Q8Qk0n/NygU6aQxqseyp017u7yBOr
4APH57aOe13LBTmnuwNCFidcrKD/L1UJXWQhUSqzRvydAsCtt4htNOdQlqj17C2ygpwbKXqMIMjx
l1Ud54VgvZXg2RfGpMhDv/egHh61k2Q30jafGwrEyZT8e6GHnGNBv8g23wa64DWlmiZ8PjqXgWNg
e8R/n2rKLY6uuvBYLBZxXSnwhZmOG0YxK98+vIHms2TVIShOg+Bwb3kRrX2q3+0nzsFB7Yd9867c
Qa/odtzVb7YprUVLQE0TOzU7GGekjNqAhsysNIR2Nylg/rAijppvHEsz8LmVpGBPdazHmksYEOeg
JblrO2K+H+jUXWbhtrFwDMJM0NGmS3FPPEWhE5CtLz6nRw1fkDkdi8cJ5L46rx3R8FkMRXulWXep
MN0x3JBmGXajWxoZu65GeZSTpZzjS5IN8uDiqihKeHpxwckcBGN0ZFf+WXYmfN4LuDeg08x5SEq+
z6tRoZSmiI3oBP6M0WbAECS/m6YXPwSvMWAkf4epO6q2ANn1FjK+/oVPyi13yiTKI+xtvkSUfsSL
JrenOPsKlQlMYjRvMXhbdLGreuM7BnItfwsds519DFAWy0Yg3etk4Bk5A5XTBgUWp9VbYOOfgnDJ
gi38lwzJRdUSeAxeO/OYWNiW79Q2rpQL7y2j4p6aTjiqqnqOjVpv3L/HVlU7PJyZ5lGVluk7vwMq
xkt5c8Cfi9hVBjq1a2Q4Yz/lKuUafKTrSoAmPI9F9dPtcH81iJQX/d/6J6IUhznST2YhStA03uGH
O1K6ue6JKxyke5xllOpl64IgJTYE/hi6QlsAq1fs7XgjOoQPHFz+L6aQ7vAekTDTahKFZi4xRq+3
La9B13NhU3GYu9mPVZUeqKZ1Tl4fH2dvzT6zv8jK43O/VCuMWll4IDaC6NFiTAhSflMUcoyiD67v
TSOS1VPZM/b8aq/xIcTE5XBmi2aqiku9RkypXv7KOpVuQyiH9X0zLoOG4Frz/cZ7fK9nqOq6WHjt
6j89cqWI85XLKcUvjEw0EMU8EiMkZw1FDuy7x0kBZSmlJ2eWC+hCUupdNuSJaXYouVmRKUdZryi3
xAOJfFGzJ16QefGsRM3W3rN3HxGuFrkpI6MUqpI5vDzKn2Ue/ylfjyYxKq8R41itbBgIuHRCPAUL
XnxKoT4V7XUvGjilQRUKJ0EY7n7dzQ4YP3z3vDnJnw0JSZM8eQvWwtyNxrwsJWwcuoydZfJgA9Fb
Jndb/tuasOfRy2DMwq7Do9WtAUgrIPpkoZeMbTd/ZpYGBZ0bzrIQhwXiMAsxOnsL8I4f93G5ei0F
NKLhSrL8soTA41RuDl1xxu38C01tTGJwMPIU8/lB3orb2o17Zc3qntbHzqt7uw/wQnn2iQYcF6Ng
HjECB+RTUfwXsSlUausTFkcgn4egLAAeRu+CE8Mk+zgYEUJQqWejqe17sf9baYW6SmxWfzcHye8V
DbjGNzkQJuu7+B7hUQScRsDP8QZOzmtXxurNygvhKkZFQWieiIZFcR8/ihBBZkRS/Dhj3iT60Qdn
p4kizc81VhvpfNJpwM63kt2i0M9rgxOffTcVzgB9/F0XAZxHX4WXad+HATSxJhG3iY+biOtct2z6
xxZw5c+vQs2QZL7nL1X8RiQaNVz7LBvirQe5QCffpSSrUlOr8gF9VCNQPw1zOdIBZNfyVmsJgm9w
j9x0PpItxORU60Sxsr40HbJPxN+mAhnsghoObA8cDmbeIN5cfIVVzMLnFX4fnSFxj4vMWZiP7h6C
loHXc5tq+tp5AydFflCkG3WZPOppJ7ds7YVSAqcqMKLmYNI7xOSpiFVQHPHTKgh/fAewMpJwfwXU
cOxR27VKqrsb0zBkTKUOAtLdYBsyW98vtpdRuOqyKcrCQCprvpRtQOn6BC3b+hmS1cAWKVbfI0rF
L5Z0+Lm2Rnjecuuw1yXClm7IU5D6sGQ5OykM+Y8bKnXtvuYdrFLYHuHdBJ7XXmheMFv2Jn/JCbe5
I4BwXGpsO70qCe1NdUzrrqXrGrHx0pMtYtZbUStT51nAKVDXgheQO8eXOjjLj4flXOjZ/eP7G8nt
9XNGj8i5OIZIcgnHxmjpfUnaM24BtNn7L3hfKVcRwTQCd/b16zBlYwa65vv94NMEeZkDzI91js5e
4Zkl3dkLgkfl6ebzPytR/fW84/Zzo6MWdhdwqBeq4jv5U30r+7/65spjOXnsqfIQFenJy8eqf+mj
gSu257JbDcNcqlHdg25nmegJRD+a1/gH3eVE9qadRyG8iMmqBsa/uCXTPwQY7HrUEXRGwE2DvyKh
QRmg/d+7GbmyXOFpErl+NvwfQdQUyngvacEXE3IWFhfPsmn87U1sEteNLKvujBKqSwDAGVmor+dZ
VOnHqRHFXs7rnBzbPb2IEt4nt+oncEoBMKK8WGkDdTMIjPJ97057qfAu1VtzbN0F6b3eXVb0dAgQ
OkupQpZTCF2j8loFOediu/884+q3nbcH39UVOQX3m64EhSEFqco7D5/i2lmWGH+KTltri3zE30GP
lBb6NQFlWf7kijAKNWbDt6yxXTEcejc0V1lG6F45h2obdAfkh72awkVReeH+Zq1ZfSRmJN6llCz0
phcmVkG4yEPHIU6S7su8BDpgF1o14oUPqz8wUhbF8jqfmPcVURlbvYAgU6575NT7C5pXlooiHOaa
gubIO/eRALC0b9AheOHC+uCdu4pwJuaUb0CZMeB+RCl6viU1XYPZDwMJ3CMR3X7e1wUB7tAdqDW5
J6dWjpZGXPOj712SJVpQzxGY99hhi5nvQ8yYSa2/PQW8oLdulroDTU2irewVtuspOw/h1rgrsL9/
pVvtcoyB43OQQ4yWFHUPIHaRT5bHp6o982P0nkutVWqP14jPl7mzVdgnqghJ6q2JVkM1z6P6z5YH
HNyGjfC4AUg2HXTwI3jVnIsmOj73tASNE01QnH1IsE7pJUMIMtrbfLrHMA7/5ENtWT0qIZx0WxTo
drbNmhXxEqsVFpVIBGyN9fLINmSVFu6PZ6w41HplNUVtX2pHds0SuTJceU3h/t/fd7m/uBqAb1lC
gGn447n56NwAwjB1POB127EXncwAS9U/uTr6PlOFaAHwdgm5T4e1b8XV69krudSADpw1L0uz96F4
tvp2zOlgJbFZcmYOCqAKc0/dDUfZVxoev7IjTBlO+cfs6t/mn2rGDZqq2aeXJ6Dnx8Bfai5Ya0DT
qVSMOhwsiYti7OwuHjzr4HR+gIlFR/9KnSZu7vwW7/5S2HuUMI6CnxNa9waMqOYl+wBDnr1Gm+BY
4VUBXzi7k9N0Be2wgy7Pzn4+ACoh9ThpsmQCM0GgVhXPPMMGzt0EWEvknfb0VcCtqlAcy7Elkntt
lPA8OT1+BrIId9h5tgvugr3JZw44WL0X7MyDUcUfdFj2t0Fl4ih/0Qog/0qy2rQcBL27sNnMjpt3
Iz2hMr4L8P9mEUWfyr7r9GEy0ju4TIe7Ncsgwa7uL6RpI45YdHLbjK+lGdApJBZpLb8mdlNNZ/32
VwKEV+5fHnAIqkxj36MiTLIwxQhBOgvsjW9VpSzkDoUZKAkrKKVSxjs7mt7lJarSHVEB7oVkBnDq
PSwS9P5NIHWD0i8r+zyjoQ9HYR59sZ3gRoEl6YqNrGjQg/TN11dP9IYoE8GiV9VVMMQ3zXDSEjWJ
2brkJ70AVhcQ9lDD1XPDCQV5QnWiB3ttf9lWMLNscj1ANfDMvgtFg40wy/siquAooidN+AyKhggV
G06QufKQYFJJpkn5cd0YB3iFqRujlQVWe/A+P4k7olk0jn2v9DDwvsSO3D2vPhV/WCwTEQm36/2K
hhIFSPsqGlhQca7Qq2dp+AYMEIE1ybNQbGWzuWlmwjf2yFrZNIsCSlEJ57YiWKtOXgURaaflsopO
kEuuWYRb80TvFNAUD6752Gk3tqz7q7MSw4fzobhpxJQ2tHp30GnYso2CWlkZR/gHWjiN7hD6D/+h
wssRxy6J0h+vMrBQ/4gsVWncrqEbwULddMrlvj0pBQEvo2mMGh55yHaRUMl2ChIJSrRi1g6zBOgZ
tkPlIqcjqVPqcqQk1O104tiw+StoKsBCT4QfcS5DbnXfsLEPpDFqEeISdUOktkOVOlXd385rae6Y
aV4U5jU/NbmFlzYiIuPUSsC4PuPf2LdC4wM5DNrHtZxcKg21bTfwcNAnbe73EdkdF7ZvXK6YXxJJ
6/u4JKdmd2cmza6pf68URk1VVAzR3Dc7I7BYx1e/R1Upeh6vw5SvjVEw+rN6xBn0n24cIcZTCijl
CH5D0FYhAwHvsc8yeTzcOr5/NiE2zKdHrlOt2wVGtXuOd2Sjj5GHTFsWqvRu/Yf6URErqYbcal9x
rdZsxqCZ81vnXCSOzqFS8uxPJBP7gNMg+l4Cgc+LpMRYe6Pr8LAxxIe0Eh+cOCN+CrxdbjMHVtDZ
uzJp8A/t0l/4iwQp4NTMx9B5s/HP/0iaGb3rmK2CSSJg2VIHc8e1b14yKB0NxF3IaLhyF5gCtR4z
i80691dhZWuOl8jZUrKVqHAPWTYFB03iXHt1pqkAOINZ5HyA0O6C4hVHsVhXnTcF+3kYRiJxq+gP
XjQUKZvaU3hIscTLM9MQxivSUC4pCaOey7lJpUOWlwOyJNzv+Y3n0joh271CSxIS69d+cMLIKRDQ
ed9m6dHz8S3qFLcOs4LRsvGuofOqfC3YPp2mC4zSxX/e2fazVkN3Tm36B+7qve+h6xMkNFnLn1o3
nDgW6Qeqpv3+tROrt0U09cqEdsJv74fMyGC38jL8SS6dUzv0T/1x21l1b+L8Lb0MTJ+73e2u1lnG
kU9kFA/T3axuRP54UifZNXAJU5RrZxElgm0PtN4xKTOl0kHPIs+9l/5XjceOFklBDZDwwbmKLlcl
tT+Yopv/stNSErXAOSYXcFT9s4yw9g8aTRohqY25Tzo0uRkFwfVp+xOqK+9oT7rctmw9n4ChF5Jh
4N6uSI0Kpy6/Q/FaMLeE9i3fVToOcnzj/qGcsXmRgXjrB5bDCFAuJOl+dL9AQTHwrsA2JZ1uWeOM
JmXUPrdYTZMeQDqhSevIFd9ZobHYQ6UDLlIdkRNz4I88h0fgLDnvGX3FEBKZmyoO3svvsex+3ogT
D/g2lYsxH+Lt2CVnK9/UpINSmMAxpU2SH54h+sqxS6d7u+BJ+Fef51r7xe7qtq/WKm8ZOa7+bIKt
m78kraR4fTYtd8PaV1ue8uGqovTENpSOniLCK5MVqEqy6P30dr/E/nfRQAykVkBWNwLIRsiBns5u
hrYkPw2p8KX4o62TP/keUxE0Y2EgYJbmXcv79y+mpa+qBrZyv6491Ue3rOwCCoKHvqq++m4HJHUV
cnMRO2xKVFN5KwNUYRFCR10ohirRq+KiP/sxCwHCcrbAgNoWKwGEkFvzFmzSIM1sOn3Ghc5kVnmT
bcQoqVuZ7ZKzTpnhB5FsukJklG8g0wEwXBY7mJqnKtuU3YGR9rwZJLyUGXWchjeCQ0/PkT1LazTk
Vu3GBpNZQxeSAQ7AyGQPATf7asgoEB1PdLzm27InnD+h4Xg5xLnX5ULXxsf4XWiJaEiJOpRb+paE
1wByPw/h7osldXBwVDPmG+bAmu3Vke0DNmqdc2KT6zg9keQjevSH+7bNejdO3KS2fg5YNJNgiNTY
sjhJ4rsk7QRAwJV+FxmcWS4jQI1uIRIrOSDcJCvabaASywlFOUwdv52NJuEDX/ngxpZruBIp3B/s
UVqMrlEGhGlBSGaPN+So1zc90SK+MtK50K+DU64s0Pk2Lspw447USkkVnjHn1atmmK/rMX09XjNL
GZf6LZEmisi1kjpeFaqrPJvd+vOselISxHoMKUCb/p4LGgXTHFyiPOZshai7iha4GnXim5JmD5ke
RRVCxNhO0Pg48FzUfrYjZ7PEuYHSPKte6TLqcMRgYDRyF+r1MIhjKphuKi1p9rb1/b19tu6YBcXr
dZF7rK58BrmN2eP3upJwnSn5MAVn5AmXZ5e+mQdweoGC5rr3XC66DKqVbcX0ZJe/7MCzNxb8MAIr
E5xt4qBrB5tocfee7OZIMrWbrj1+WFdkFbwVdmZhJ/yj4FwNlDnQNfScsIltcv4b33qNDsJ1gUhp
39xwUOIAZ1wGBgX5K9hsMaxJrpWhElEcyNpYl6c8ytsyzYxuYPeiTCzqovK4GvrQGYTD/tsQXEy/
CgDcyf09w10QCR9ZMyyqAtAz8giWr8TpgQT11vVCV52UJM6Tasus3t4b6XL/RssFP49NEHrUiZjg
vmTzZTe+bUfSEM2gIJqex53EfQP2lBLHAORvVg5FqUHsptwa9Nt2PhkHEpQS2k3iQ3RTckz7N9Wh
qDkiG5A+JSVHc4unerEGgKWqjUsjPWK9SXqvV1Xy+JlC2myLFZvGWSyjpQ/TKlA4OjLw0m+EZZlP
Ro0qOjTsmlsH//lJBlc7XsfoHkq2BtNjX9xTf/j/jMsLxjGzxEW11xSaqkbRUzEz0RR2URhsXdcx
IozOdRtIX5cgbxiHW1ODNjyZ2QhJfjFJE5eq/pp4UUA3py/CNRGuzJ9QsY1l5gm0L/dzMNDNOk1b
HplWg0QU5o2tP4tlBRvFBDW9Ldxf9ycTHgrD5dC4mpHUyL1VA4EkbeEfubzHh364sCugDbBOo7ov
cfP2DPW8FqVi33CA4TIp2uGfbOyK0IFttEZgi6hdTTeD8669UH+9PwtLLlb9t+WszHCepzCKFAWv
DkZ4dIByWyaLcEmhiaPr37RgN7yjCy/zVVG0nDXFZSSzpq37WTIivbfDVpxaKk3o/eE/D+VcDDkV
ADv0X1COQVYQuImyxDXA8HzljLedRPpgk6zJfjlC8DEF04xl946iETyKpNMdwCKaUtWeB3J7wKOg
HWM10Fj5AX1nMgHuvLXh94KZS7SWKIfPdyPLToGOffnTGYmk8hUAcAa1QmY+esQn5HolxftNT8ci
XnoNNggDCYLWRsCQoxR7Q55Qxkw8G9HWdCXu5P0YBTqOGVr1kz7C3ZzMt3n5u6Hqbx4s51xr5IZP
dkVqc2+9ZQM0kdzBQt18ynS/wJg2Xjtca+Jw2wGi0FhZG/mB/T4gG+KLixrxOJt8wCmP0Az5+YNk
Er0GyUkQ38j+Ij54NBEQSrNN/wFXl4qUHATXwHML+2vn5LTUrZ3edNTCz+27STubs0GtnEugYwHY
YdpRIbNvP7YP9ddvImFweJhplTwiaADJ3ULRxtiA5Wp6W12MTlqSX9SLZWI9840782onvXDmm80Q
y0CCP9mHZ1LRqTx1dRhcOXw5dVQPnWOf/4qS4HjbdJD08w/oH7eXqjGNle3VDLeQRD6ZeUerfJqC
jjer5YTpU5DxGvMy+YCK9fzhBDE9jtoHLIUipaf1nK05DX8IhEme6P71BPIwcAx+BMWN4OgT5OBR
Spv0YYrJGFeVpbH9LEioUcwsLVtqGGGlcQePpbGtUazG6zjnCxiCYA0cGTDLkvdfysZf2KCqi8bi
Jz4g5LOGXfBz+ITrBpoQVWgFrxxxqIFOFxyJbmvdoDcTAJEfAUAiHeF/pFUWoSpiqp/G85htUaDe
Bv8IuBpxVKnDy8Kv9ohbhvfrAnv8r8c4JTOlT5VU1E+jdR6rVjekREDB+cn6w1Wb05O4pL4eveZV
RtFk8tfXhe+iL/+PoqEldz3PDZKhvNfHHmFmB89sPCoq+F2TAwIc6oM/CHLdg4pZKiTd/zPFH7Nb
ikB2QlagWgjHm5Rc3wPW4nzdkL8Mr6SifvRUjVl0kc68rytSNGxHVrSZLUZrQIp7R95iw+m6bcPR
+UHCzBx/14IH6ADabTs8RaD5tifnPVKg777VjPPTJBXe31sg9kDqRhCK2jTTxOSA6GMvgr+1r/y0
4jmzw1FlJMBTSwCQxHIqjp7qhqneYUgNaoVMwm3gNKydD+T1TcD26aSEk6eyLF04PoW11Hxr4i61
dyYJZwjkdox+i6RfV/CnS3YnugVMem2/punGk7f8qcLD9aDHXtRY9y6wUUcueUaGVlo+yj5c5o31
ww2uvlUq+iz4PSBai0ZZDmHlOPpp5/+zV/8OK/Qt66MtcKB9FT4ukafACGm0Gn2rbD0ADsmgV4rP
VkADofwfHYDvB4LhfToEXEFxDoYb/C7mMjgI7NYUKXOL2mQsdh7EYYVTaZNz/1hNTZSP/ytqZLuR
thbysRRHXWBpq9F+mqszk6Vupe+xAULof1241t/EKUf+j9wK3/4qyHrTeTLkRWzKNUALGCUy0r5X
S/ljhXqPqFcK6ss+OTlEQA1nmrP69NSpkuVDuvfQGpdOUBpIYZ0nIshQ71htYpm4HlUCqKCh7ZzH
kp77y0iiiiPUXJUbHAXXBJAvbzHaXdF3AY1A0DVm24LvXjQvfidWpP243tXYq3WKlVNhIqlh4+p0
Na8QgaB+lN0CCuWoOGVbWQfZxOrvzkWkpJPqt7X8tR4XzpHiAbMLDQWiEojOOi1Cw3sCkHsaSakz
rfrCD8PSM14HpmqrZEw+8MFMAvhehruvlevzsRuKhNi0XtyB6tDf7rzb9ju7iQacGzjL3qMfEqTj
sATGXE/HSywPJlhss2D5bY2ORqgDfuMi+zx0QtFvlPTtPuaKc3kFcqMdzX6F0cSZhV1IK6RF5x9W
UWg8wJohbeTYfvkZ/Gnrb5OMn0cUzw2lVy93rAZIJYo7n0NYEAcgaggdhbadr3IvWc3VwHQyYfFS
JspWQ46EqP56Benu27QfeQJgawThmPsptE5yd77uzHB7UsYj9AXxPlLBtUV64P5Q9iO7rhf10SfR
NcpXrR5hjIgFgbZTLioBwQjlXZMo80WcWFBYlrqTaaO1b9GUk9i8iJXYwQMbzcDbNz+3zEntlatC
kAC9qcxtwytxhOYxa97JMI8g207fbAucmt7t2TnbLliqGlyyg3Z3bNgExvaPqLYHlkVzW7abG1uL
r/bMFxX257m2kJEfas2BMHuFGjq2AT95kvDi1ZFMNqfUIVpq2gTzGui0NwcsHRSUuHghh/K0oC11
QyFtabJLYzKh8XLBVxo+QRv1pB2Vf2Ni4SBx3ZPdDG4cHNDOpHNcdUEMLdycocJv511ZtW1EMtAf
cDd6Pgbwf4crRwBwKWNzdQfKkPAWd8i22MeXie9Dvw6sTnTlPgfY70Y+yQv5Tt6StQ9nINgsTgbT
75JDaRFpVyuVWaxt8Ppck2xTXu64f3TW/okUwRuGlbJkrUJg6fterhIfuahfv3SWpv3uG0TQVfRr
/+iucl/zQv2ZDNTUYD183+xfhZAaxNMTFBfWJRJbbUHN5WMx1J5/X7R1sf6/VnAjuOSYjzpAG50k
ztrrv+QMxEie5GppWmsTI8lPDXZXL5FQ+i5ana3oSLnlLlZ6qOmzeXJMkZOXnQWBm/7i5Aos552f
X5dRGBOhlDOeSAgsNB6JNypTdRDAak2Hcf9VslDA/oTCC+a4dghuX6JYRq/WCWVv18qaIf/L+HGP
3zI8buik4aszU55lyFzOvHxCWivVdFj3lYIDNwOa1DFyz7yGG6bGkLKamAHZDBHUa7GvH5+8j4MA
56dx75QQInT+vEa0uVKnRiOVsCr2xSY+vs9/E/sH9oZGTqDviiMHFwnwwSitdcFZifrGzEvNW1P1
R7dtgUmXJqgDZhQS1wkq/0TQwH9BzSzji0szBlqpmyzaNpu+LQNoz+XlvEI7GFQSHRjsb4dki9/g
YSkSqPcHyrj0Y0qpmDLbQxJZCyrPqEiqnX/2vSW5tMYpHvudQPm1pcxVVTZo4qoWF9S/U69ynhlO
rTGnQZGZZ0j/+7miZtGjdkoB7xRQDoKntd3s8Dd2sduTi+fvB0rLGt8LZAsT9F1YV8r6bryzcZ24
jOZRSUb0KEeq1Tum1OpX8YMagJF28EOp8a+oP/e2LLRbCyrBi+fu8FWH9KirvoBgs7N5D8u8lHSI
2eiqA50nXBFLv/HiSL4KORIKGhysfwsmsR5RqqhNALb04soaW377HpoBYE22rRwtXtdWuNqgJDEI
3tXJJJpFAXLtKr3mvYuDFldlYXFqCeXSuETVcYFA+2IFGxfKSsjR4LlS5JfuaGoN2ijxrK7W1X3t
xGzD8tDqnPm/9F8Azs3oEd497bKLYyJRVUWHN06lFCmkY5Kztszb0jjh9HwTc7FpHbcDcuuAeCZn
/VWJCMM9QLW4kblRxHs49EwNyg9MV2ladPi+sLuDPBBrYDuldxJQQeWyYbxDvCNvGBGiZuc8Pl3q
rTHXAv8Q3mI/igpRjGNIrSMT51+iZuAdVxluTjZxqeY/ksYL3DNnZEHLZ0+6MMuCiIuIBldQ+38y
mNKABbGMU2El/O34nAYJxZ0BOruqGvabyfllqPyJqoyQGRBEDVmHfkxdaXdkgcCoyN1STQNR6H5f
wfCyFofXC9dsrHuf3K5EJqfYdbzLU2k3673rl1BL3Or3PXUaspE9sykSt1dyVLt4/Wd30Ui09WZw
SkQ5ngOuFGs/Ueq3q+CUvjck1IUVnSYqISK6SfPV2rdQ7l5mjTiz863x53HW0lrR/8xsxrjhORUR
i6hnKIFIzA2yGl/lh5GphOC+JfaynqmIp+Gsk3eF5RrMgS+GtSYGj8Hv8+74XI6nykHt8hWLmmfR
FbZOCc5irvr/L2pahvCtQVl/lRWxwa9c1hV2fYHJkcO9oRhnBQs6lX30qLeICTjRGUG3FXYyq+uH
PmGAV7XZ+i+eYlqBftvwNqADQOlFQ5HYwzCVyTRjbMiZnkwOYN7oLKgI9cvrNKwCTArfRgCwmOKc
LZNEMKfnabPPfA6Mlosl/Pj/0gOjmz6HEAPBA2WrwYK8OcIxN+UknEnZgxrQRQWkUI020WUz2+uw
r0FX07fQNTQjCSDzzKKkSecjfQSWyXxSN3IR2x1KrxcVTnNITUeHiITj390WNQI550PbjjGXn+Dn
PhxmaKXen6/+1HUjuAU2h11wbGWKHXYtNC9nJGykRx7mtkvxzJIU7fXtIvNNA2PkC5IL/LlbXeCr
iJFi+7GebQC5/JM5oFDBNBCWdeFG+lGUiYIBE3hmTnuK8LSfL+8vi8ulKiuCIeNVO83NEL08MREf
djVy2D1Higr0AeJSbAr8BxP0NzF5wQcNwPVx0XRtOhbvpzfRzxYQsBiDcKlEjBzWq34cUY3sCL26
mXXbvxTAuuTElCbdaA9A/RIrHOlWiyf65YyFYaXd17Mkjk4bysFfPkxnGL9ZU6UvBiFwoK2eblal
pquXSUfdogpf38wwG+09ixjIsTO0oowNLrWzCCFLHkKq7gJooA1NjZRCpoLQYv4KHxjimANpTF+I
6pSkK6k0WohBSJzME7Iyq90yr9usVM4SdX4I3nS5gd4ThuKHR/8RlOnyS3KOmcuBHrl35QJP4LbK
MXwqAcV5WqLKzWPPiQr3SvVyzathF2z4heOHLj6l4Qi9tTK0KITP5kFazrNpNXDMpUprU/xy4Pwg
woN+7fCnQWlFf+s8AkBF0KD3bvDXjif6d11RfnaCuuTPJldpIVdtEOX8lVApiWPgZS9S4e9Usbs6
wQM3WTRk7q2GtQNc9a3SBvVn1jbk3BXkfS/f4aRoHghrtibX9TW/uyMt/s/N9LhwY2FYJXpGYUfe
VrEA46jXHBpSlnuwLR4GSPu8G8O8FbSZ5h9dAAgBV4e0CF8fJo8mBHAxhmYCx+/VDYhrWSHRR9Uk
99N8U+Wm1bqp1sA14JBjmDzGiXY3XnvnPlYlw/JjlLxnxzB98rWqbU9xLUm2XK5vJ5Zsv8pbac71
LpWwYe+W5AbO7bd9t+WSOa0myCs5jR7IXiR5Pce6PNi44P6AdRadtmQU891J0wCY9s7Cc+xnj/nJ
sOjcG2W3oMnSyupcyFsVWeDjeqFcRARzXA8seN4jlwaAGUzfH5nsSbOBSS3E3JhnqWU18G5Ij+ki
sTM+yGawObns2rzU+XoImrtaC5HkEAE5kntdMJ0Mwx1SX+JPNBodJaNhaFF0ou+EEiGjkRv/71Pc
7KGGlurgJd1+JC5rmx9FQtkFApYS538EhHh2TDFlUZtoQ0v97eUkgJCEM7v2kpf/S2MItNSwvzkX
aAzvkhsRv9tIDqRA+cQus7P6P7RqXxxK0b1wT2HXs5IIPaTCIdZQTIKo5VY75RgUw6ub4prk8pC9
aHj3ZdwnyikRNAMQSX0TLupr4cyXuxuuZpXqMTmxbw/kkalXKyqxFwKjC/RIRiaKGSZSccvmBmDj
1Cl6Pji7++54t7lURVD7LlGIp+bPRG8uEb5k6tEv1BmMazYiI2R/oS0myVeU39SPacuV9dfxIVR/
nY6Y77tZSFSbnbevNJkiQFWfsFBdZ7R6gk5TRDfr1MWUJ0FV8EMED7OZHeQBxL2uXE2NbuctNihd
4JbTqXN2AQw9J0RvhIDzBW6ofMQ1ploZPiGfTJ4Z/nK7+oese99IENfSbkulQjnCIrThs7Mxf6We
YJURuhn6VVPnGWMcfezBUD9HMjqu7eamdAjG09lT4AyW+feYEFQSIhopaJKN3iUJ1OPDRQtYP7m1
J7enx+0lkpTAuZifk/S6V0iwUr0U+pPslXDtdoBJNSCT190ep+JZ9XXVAyRVnMqPJr1DD7AQtQEI
JTHdamOI5xD9hpj1jbEUa69d4YAOHFTW/80rgvYxHd8r8dvCNU7q8uByDyoXPBbxFDcugSns5YbQ
EdtZRnkTwbMzIyeHkuJAY5I7nwFViq/46Uyt17WMm6ZUvudBf7dipcUnkUPdH/3EyaE2l2bmvUOm
EzSB0E+DhN4nn/Nr9Wp4TsCDQNDUTn8cqbf1C5UbYGajMZeLu56e7qvXJw2GDpSUPKGzj0h8O6J/
ox14rn+/4+2H4mQXGbZXXtgZ0q6KQcS3eKdXQJdwFAdukuwnux4PYPpJKJd3ZHaIhHtr8nAdZqY+
lMcv0AFms59M8TLD39XgcE8DmUb8d00BK4c3kqbLQnufAeuIJDvCYadHm7tT8eqthdgaNnG8X2vP
gwXhxjk8ihJT66pQ2/oEY5Eo7vZbvodPbpmwpNzNv7EEu5fovGFfQXTHkVztWhxEGONd9K/Q+lJW
wU6L4d6ukaSKFsoEL/3jye/OAbRE3p9KGyExnN7bUkKH/vE/GLCHxfq5ezxoWQPFN3CIiu59X17a
HfZWjWi3jfRfcj9cSXfX0nrw2sZ04kroddWfqsT+oTAaE4HegFqll62ci5MASkLOSOhSmNamfV5J
kK2IF8ra/IXO/Y1gl9p0aW71A+lQH8wF5ImjJbaoCU4I607ctJDDlbMw0uVbLhgQUkqWjsZFWqzf
yIPMKU4e6K4/aiejVtnZG1M80MWFKc54UMLJbGugiTkPd5LeEqb1MpcuXobbWWZxen1HRi85LRyx
Q4ULlLD1vdxycznQvsLVfmxwqXQlqGmPdPUZ9Ee90r2Zx7cIDRT8Kys3cUGexIzFKSGnnHOFUZVO
zGdfhBa9N8odQgZj6L9TpzW/A7ZZTsDKcnpPc02t9HsJIA3+0grDnqUPWUjGVZG02EM6SOda4yFq
hlkytNtXaGzthb8w8nD1tJyAv57KPw8A7+hQU19Je+VBu9RMwwPYKvd3EAzkRsE/YS80aK6TUyyJ
wQnEGThBb/0bzSo9U4C9VK4Th6ZkCSLq8cODZKZeB8caIaj4j6OSSwVwnSWiWqgfqQFJB1vIWaLH
/CVNY4Y5rAf93z2DAis3W6bfO6VGZzckD91K4ElUKl14VDWRPDFOV3MpAT5ticTOetjK6Hc0uyls
Zu/oxpaOsI4VIgpPPki2mSBIRBoeAAHAmCeZ0ArFOy8NzaSTnKvBJzMOy68I2HaFGVSGGljHf/L5
UQTSz2CYK10YHuHaTpSfbnmUzATUBo9fU42km08+Ewm0GRQnyOZnRU4AzqP/lreyvI8H02Ue1HrM
f3KWkdy371rfe9N8NIrsOj2KanSA1Sd8hMQBoAEGygb8WO9KtyeXlkJjfTEqhWdFUwXLPNVb5uQe
Dqr38NWOm7ebnW8XLwIUyrmtrcdeomOvJORDy+pGwO349Bio6cfkzmDqKmSxuRDMHa9fNumaEYXp
e0qqyeyIcJ1Z9tjJ11irSsyx/DQopWWSgHBtEQCJ7eVyz/R8FpCKUP0hkKmjav30YFE5gTValwaW
Pb7glPlPdMSCRRONGd3GaqK+QzoNMWsn97j8/fxSJaTd/Xi0qzXCi7HKP3kQJAgxieWJPBniywxN
IPcYBFCPmPq0Fq9dHHbHaQG+3AUd1mjsEowkXPQoty87VZYevWbOd/rcqyF8LDxViXJxMoI/nFEC
C81We1yHyXULRpoMExWp3rdP1MEkq+0wLIYZvPB66B/ctM3Ur60msWwwBVViHPEfIGmKcxRokjz6
1t3IM3jtJeW7rs238kdHIuojEjBSTm6Xh/F8HNg36yCIRjn4joPxP2bF+YKU12etiS9qF+Y67U0M
3D0aNikuXm5zjiMLFxAmrg/PhOAYinJCT8+MH1fiKRGkzpThkE99hDqJ3RR6p+Pf2V2qhjr1u+xT
u7C5I8Op3skIvJNNyVQMvn1+IdgnjvTx8q1yeLnARHvZ/fUrbgyPhu5cDcnVO0UYtHixBbnbNCug
3P2Zs6N3m+vnBLGwHakEkxRKK+8LEtPOQWFc9i9xR78ud+1GWNlpLdq96rSTSZexsX0zFqgd17+P
AxX+d5cREwmzORgnTS3J8sPN7zGpkd3RsCsvjzfmzORtbOq4dUDQ2OcJWFkjxI6djYTKh1acdDKb
+46pC86h0zrVY0Nxl1uC5KsLqp1wuu54tP5g57cmzosXQfXq6037oWWIy+yGYPLOK8fUN7L4eXz+
BfqDP3aoKw8GRLEuY/S7ehwsw45lrVrHSMKkUdOUWKfQ2TDx8M1xSZ+hDjY+huSnrDgihMpdvli0
kvwn39BtHseSP6WRg49ELOJY4kqnln0V71cpXdQp7tFkpn6HTmYidKvTNF7vxwL21IzZ7CIb3has
5kdISdNuoXbojyNROwdzLVlOMXyWSlcVldRIOaOSz8fSg8VKSBTCvz5lx0BUDGXl3BT1iFN7yAqh
r5uY7uT+wbpqrPFc4Ct9RyvWkHI8M9PoIZXD4tnR60ActoVuCW5zToyCPAPgPBYrRgLFDQ1jQqMI
ZoCKODbuECGd6VTR/27laYaAfyBQahjgYyxAQ1hC5NQMtaq5U+6swt2cMeeE6eLrFP3Ae5KaBvGG
vujozXc+zh91rrS7OnIhY8+5k7HfKpStLz0tJWnfU7fehdSvwkMudUCvFVYy3dwViifkg0+MAiL+
Ww1lRfeidQGHAHdtR+Xa4eGw90DDWn+A8Q2j95Fh1i2lMNA3BHpeZjUjQbn5gUEHHlOgLbwSl8yp
ytP4y1eqzQDPzksb1ocvmS5ZpSPKlKd1NTSwmuaCpIERZY2AWBpdKPoTibIpRhw3AOSpWw1xm3sD
iFaeaxHEGKYOYkW7ANEQNyw9T6uEJYdBZoi/uBghIQxWA+zi32aal+tKCr+ADGE50y872585nlWG
Ag9qfhLsSYWZkMBParawN9SZwOG70TVOwbjREtP1kqSMcQy78fl4+5+KhfMkSoBzzF0itkNO7JEU
BlpSQEzzYvWuFu47eFb8ITeSRkeZLXVuF56DbfZHkaYxbWXyBMJ0ex4UdYxsW4aGjt15oCMnGXhF
06NvTNwer+xUQfZs+5ORj6wV2BXqJjS7sRUd3Z9MaJd2f8jr5f+IaL3ZdkoitzwxnrtIYSEt3/uw
LekN05+/iuj/qTvqEpXDNkXCH7mlWvB9AhG77RLOAmvZ7d/OW4MPsxvAjchJQz7zY2eTxJEpDIe8
vj82eAzG9PVPwAwZ1XmnqVgxqMe3xhjnUzpDYRiHajjvAngtI3PScqV8m6CvnCgU8tZq2LFKFK2n
2loD9qFfbBZ2Vi40ItHLv5zLxj7Hjz9BcsFQHPmxMK7na69rL6k8Emhje77sSyXqj536kVrcB4p8
xw+lQS2YTG4dDlRRqJomqk5V5/XDeoHfxAYTOtOnMMHoIql1CUMvSdCYMXmV8PtNtn/j2IMMqDwW
alU4mlCg8UkN++N7dgcuvdQrmA+BT2LQwE/gunJoCefhSkrc8Fj3PCc7ZxZZlgUWPJoeA/OXu4d3
zrdUdFjI64BfjkTqGg8/38he0srH6UxRFbY25MpPVsk9zcDWZs5124FMa5gnKUq5lWKU2YQFDOBa
zdkWo1mpzP1fhEQ6SHaamJHhgSzreQ5rB9pBw6FeU3NliJ934JPlHfVGq15AIvv7OpU+AbNxYvZg
vaUgGe2DvnZpo5ZeC6HR7MtqXCSDvOGFytCE2hq+KVzgxDgZuVHSBDZ1SFKNkPkSTY5o/xyjblk4
M9go0NyUlx7he3GSkiWTuzh637aD/ZmEooNelq1ChBhBtmlKW1fF9NxKiiI9oRPpF5XkBffSKztY
s8w6NvPCinHyiwqH4ViXwZ2gvMlwLjAQQ0NZowm77OAMMFiBY8oiHyM33SXUGj6IUmBKHm0FW9P4
RPhACr0UHc9qW91ZmWAEB8Sw5AN1EZuYCzEgwqFhD9pr9DuwFi2tKNAA6dD4D/JETk3lGRLui832
3wZXrwYffWSevDOskcTkDugIpYmcjrfsNSDW9DuCTiYVJ51ElKgVTh7Pinkzy9/n1VCHf6kkksse
HDI28JZSkHKXzPb4WclkKLLne3H1M2sBaW8EQ06+02EKUiymS/bXvGftbyNEuTWi/OBlfPMuUvok
LYvKQpI5jjGe71ykTZYfe+QmIhzinTtA79zRjK7fptsRJPznVBWH2Dqy6EDkSAR5QVCcJrkYOYKd
z/Ol+4UjimXsjm6gkv4mOc5M0biCGAmbNXjXWyhoMbeqB9qwWm0eLXKdCN//X67dkDLblIjjXHT5
iZtzElXITqAKNCYEXJH/2r+Bbd+0vW/Jlsdcb2z64VXNsNM755Xggro21tH2PrMkqA4qveiTS0jp
5+Qwxn364PxjtHG2M9Hxcrm9tkKiIFMny1Vzbtxk71IAmt60Wh7ZdscWQNMvkSVfHSUDkkwMuzQd
wRr5SvA3C4ZWlBcxiyXQjESQmGSm7g7UDGJoW5ulRmGS21j09goPmJnWO/Xn05ZQlSi982hdoK+a
GrlDOpoOriK35Or8bd2VRcXfB7leuB821dKWrVhEwORWxs+zBbORWqN980i2kmD1d374M9pbK+XJ
7rwlAA4wAZpvKgLH8XX/K2L9m0l3gC+6AWoexzFpNt5IjVlwC+PXSo6uaSTOlTtjILn0i6yFNezD
0q+GkDvKoBGgOy+eEOCI4HtBddo8rKsPuyoBXHADafFo/PCVgqrdg6T8j/YUC3Kbq82cyXojSIZg
dtttf304Q3STpJvoP8hAQid8eU/eq7AUK0aCp59rJnQTijyftz4bP8o9ELLctGhXADRztqHa+gSZ
4GajBnwy/a1y1TkyL1sKeK6gYHWmc3OzkA/SW7SeWMx0cuxnsYrFYRRcs879Jzy5WAhUT5SrB5ww
jUiLcuVgPc7pY/LQ32Dw28mOT9e3UqN1ozKtbGUM2Q5uowrM35naMpb1KiarTCvAnw0xpwBp6idI
wMw/9GHVuelcRwg6Myz2tKXFLHokL9hyLIQqzMtXWt5K5qN3tgJQAh2HdhXWwntW3RnNMZtDEZAZ
gaj1nE3YB02P2F3U6Pjpux1QMEbhP9V494qZjLO2ywLYmCvbdJKP3cuJhUrO8oKKi642fu0MBgra
zDXqrgSTOSKLbXsmtzhNN+uiY12oU/Meg2ErLNHWuwDETk5giDwtKUvu7UwKVqonHs699TqecnmL
it/GG26NA9FhC5x3zfA+Hzmy9dIzRI2ooZwFmYUq3SnX3wU+mn/OJJ+dZ4jsRFx+L0oWorlvMYKC
8KYJ8Kb77zA/US0S8DpwTLYX1PQZbL1TfXHcXfVj8VohTNiJtuh0dvJyxllvwGtnc7jI7jik6j3E
LWxByJUkfCyP1ZzVj6td8kO5JPW0A4H3hKhEGjlI+Uu+KiL3H47ymAdKOXf0+lHYz61EV8ckwXXG
22EHNq0c5JrdIYOURayuq+9FFxYoSVNWqP7jxV4/g+ce2wotoCb8oUT84H4X6Q8f2tMaKA1mbRKa
zdxhK/d90dAlB7rXX8cr2gADaOAjVXWuVgGASwBZPCRLPnOgqHdEkUCIetcwys6NLDcl+DfdlHBf
crFPV3Kt6TbaPkqcVgFS5fi7qAVvR4RvcIaJbXtubh2apvICQMxqQDFZ+mr49THKYDAgV+0YiDv2
Gsn4+byXelZ8LD2Kqw6OUdMmQNC5ljRk0hrjsZYgoU1aUWd8o53iwvzhEIoe1P7KeXrn15mZcJit
kelKL/CIsTBxCUCdJXfSSGNaUrkvvOroZzvxL5SAcg7pf4JrhBi0e011Kjz7PbFUn04NN5RZxtKd
d563mAPwQfFgsFq/2gArLEMr8umEs6xGo/vpiEeW9w2X5ZSvpOwPfDmKeeb58HnOZCMBCnESvxhX
yetdHoX7N6WbnjFeutU+A17x6uI59rkioeMxFNI1ch+ew8RNt6xOZQ6P6XQCG14Zmz98Fb9j0L2x
t+3Ppq+772SXWunEjDG0Lrad1ZDEceaEd87ZqIyH5wG/FnaXuVGK9lcf9rsagd8X4jYga/pkSe5n
BHcaML9jOVXPCr2hEaPetC9JPV9Hxmjd0N9jzWObyoQ8KzwLdD25EhaMbsD1/F0n5r201UqEQEzc
GUzagaLu2JHMMRtGFni5vuIMbFiWwxmfCqI+27G7jWWNu8fvrC4TeI09B05GDWOFtYlFWbPnhl9z
OqN1TP/5O98rEzuGGIkINmIAYTc20hKuTuaUp6KxKWKjb0DK0bSmQ1Qn1u9k3RQObjz+IgPOL2XN
ZqgK0KTnFBzlyiyTgAB+cTIXFHDTcMZVtW46B6BklCvNFxhiv5/S3wwrhV0/QJt2yQ2Xf2DnWmeN
gkMyCjn1CeJArmrUjYckLKHlz2tES5ucT1gt+Gp6wiKra6/kkuWb5lS5R/C1ar5YKhUfmhthtush
LcvgXKxbf2MrAE8afIAQiQZszfnkLc8d8QlkHxHhMViZaTi0kQK/w18iHYRWj3rZyYFQIjEdpYla
syLuo0yl3WpuIriGk6pThF1iib+iWAnrXfI7TwyOvcM2AII5QMzgLl0WlLZgOIf2av2WuLU+Dn00
OMSkjbaTUJdFQxDuLu1bk4Thvuht8vhYVyimUtSmc4R3mlkI2c0J3CfZ2Qe/7zxmY/JjOa1Jktf/
rOrIdumfG5k8Nt8fD5Qf2m63GxZszYi051xTxoDnL+ZpH8zpJaitw4ztapG44KPCGS1yq/hP/xPN
/1yS+Fd+rqRT3iaTpz0em+jOAzMwCj0gopoMPDFx+umEbJivLXp826A+G98bJmbmOl7EDj1IpuC2
FGeiMCIZMPz+6ykjE6pClrNlpG/HDlnb0YK2cjiT5ROJc0ZVKHllFEM0QvnD5LGgMft6yxzCd3ca
ik/21n8wMLemSywIliqFMIb1eIsYav4cf+dAI8AYikOrW94j3TQh29P9L5bA6BDhlYAJ6K2DfMWn
6Kac+nK3u02jS/WIXLO+H5rHixVSJD6o+6D+6fuLUZZtShKSiniIODjKwPiOz5F1rRYQBqwAyHzw
C1KHfI01tepoZgt4qA7Ghun9uWyaAGy4G/mlaLubm8dXWlfnPPm42GvZUUfwiBqvCJyHoFiFvRVB
co8VR0CDdGzC0S/xcQr5izS5YOJ7f9CmN0sV8ZY0JmX6SaPXMvnrbkCA3/xOpdMLqfqvv3vwzVEK
45B4mg3iMso4HvVZwcFRao2ShmP0jGOxnFaj+Rge2XMBE2FzO0q91mmEwcOn1MT9T3B82nAI4isQ
V+hZGmJYXUX6Vej/SpgZLjL5ApHRZW+uBSpLF2gltnhYjuGPM1j7fbdu1Xl73xTqUK0LmJWpUUi5
0qUudAhc46WLD9LKYs3jh6Qz/PCzYnX6TS7uyWgN6l1pfqcIdRGd4TWOsrpzjmAQgPwjb9xDraU0
zJktAqLiyINsyhS2avF8s3ukdGYCg7eWfyhNBOj+Ku12tUvqhrCBfOE5TbrFnFjNdikZ+Gugieds
uI1JYe1b/k9U4rlM3pu7aWlioqZs7sDwzZLIIJRhUw/qVWML/dUemwCSOtkwGzWCeVM1z1trMAb6
nsIX5IVbRUpp/g65Z7XpXG/sH/DNK4AD/xiocdw+MSZG/tVUDkVGmbtJrYj6nu91mMFZKEZtExYy
JCe7ygXvUznXPjhcTnktZMRuG+Z5FJyIaH5BFq7aJ6IgeQQIU7+yARUUAoU70xQYIqlDAMvkkbDg
vAM+AvyTy5xKHvytNDqjtAOXWdQSgIi6aP9JGOnvjZpXJ4W+man5hCDr1kATxn6/J8+I0GpKSNJg
zo1bb+x/qewIDMkvJOvQojEVHECUAGN8vqzpq2X+B1h57Ln6KFxXSkwqDxPO8GRaRRspUg7ZfisU
DQMDHs4/e5qHIMn3ZtIwSQ8aK0jCS8ZynPyTCol3ULaKStiaI77etR8N+NSpmv5P19BZ+ziyiPnO
NxGaLOV0lQQeJdvmsgF6e9f6EXdmtDUBjUkfaeBaN4Jyow0O9KAeyBj2B53gZpaXmdNOkjU5cYmQ
dtB77weV+3IykuGGZ3ClErS0FQjhLRfu4tUkftb596/jUowHQXecEPbr7DzEv88ASmEmc6Dy7lei
snSHIiQNlwugQ9jMMKhj5jSfprhjS+B4vZZ8pF6QgX/SUdrJySvH8e+jzRbx21M9//ESpkiQ5LWF
czTFgVeeqHXB3208lOXeN33XhR1QuTIYysrLgVPmSqMkXlD+5XcuzBT8eOZAHAsuKows1rX5hk0h
hONjO6YOg+zviUA4K/GauP9AEX0dPygcONAp8MLFzOTREq03bnpB7bWKUxUMF5p2YEd1xIpJ8fgU
5oHx4LegQOvAJy2y7dyT9PjQygcRl1IhWH1xwEjKFpT8bRxmIpNj/nCl3R4wlWXPH0FZ51S86+ft
4TH7mxtr0/CZPtemKx7WNv9IB+hDscsJK754zT+NCryaJDFjsynvoSXF3L+fDYExT5M/vnMEEobu
LZtb/WA2SSm4PzLv4bOPStzspQ0SepukJGNGCgzfhON14kM+ywAhcef43SJer3qnLW6GjWQ6f9MH
ZsFLZrASQbM9uKpHcA19r/UvZ0W1erQfBX6jYe2CQ//be0BuLQvYSHxug20RsROFCLk1UseITXbI
OfM1kaFKkBmm4ulbfiBavjP7g97PsjJEKNVv5fFblpe9OYyZa1tIqxI/yDG7YQOZWdITSnPZ++8t
Jg0d86MbF5f5mxoaIne8o+CZ73E84/Bbmxbj3q4IQkGb9be0/Yql5tcgp4VDYbepkl4wRc+kgqPV
qRequGbN/25xuZpaekOOqvmJGqKl7/x0gM7EuocLvdiR37OQ69Xd/kLirmfaSDGfNFmIeY+ja43p
tsL5z3JQ5UKYVUJKFICZPUotdbG0DOwm8lepWoOanTtHaqrrKZVyByxXVWkNel2OmPywQ69LA1IK
LCB0aTACPV0L7S+l/hHZTca+TQSrUapEV0bZfNU4LxePJZQC4ldTjcxpQVE4OcY3vrS6DsalkV8z
fmQAlkWS892H7SO0S/Lsd5Ynwn7n1xDnjpe2HwpLPoQAOb80Rrs+dUmxxHRD1kDJ6d89yttnx1uo
sXlLUAZwkkZtndeuZFOTFIeibJe5GQevw1h1LxoshK4jNsZzfJbHykbASlkU5IxFA9wVaVBlm+VN
6uI0LodDpaesw2ZYVirYhqPPFXv4zxajG/I7Y96rQk7jlNr5FogPWiOu0XKh9yoM9l0572NY7OIl
w31jBIBdFZZ0qZMD10NVQY/ZKyWNOgIt+ZvqukBdyqZaulwu28CBqjgd8ln1/MZ2mokTkezcJKg2
JnNSK5kydD3EXjn+7iy8G/4Agrr7oQ+I/rRzPuRzGT5etiCAhjlHw/RS5+8QPiFckerHSmicXqAx
izhwedQJ9yo7uiySjm9Y5w69fcgqSQEddBmBUs3zv5XAHktAPyRWrdDFOsnkThYOCEldAxBI9o55
rta9fKT5PP2Z6z6nI/cnRceHEsB0iZ8eyroowZRkwbic0uFTgMiaOIFJBE1t5TNdK5ra34af0fQX
HEZgLa3zA4CzTzjlp0/pGnOtQips1wVv5rJRaG8jL1KO7rosF7nTMWIKpyorS13yQTOCfZy76VJI
OsNF8ZiEfr0wVZb1GxRyACWb0AmBDoHGgFdAfPWvHIee+mkHd4tvBMn4aMemdkVdk3xwX0Ci2QIq
+uJgunDWIrc9MpFmDzGJ5Y3BS0Q6yZnvCCTzYefeGlcFmxkNE/hZIuRFxWnJmPPrHMlhlI2SGgO2
BpVRjozSUPWPnzxjeLQil1rixmPh2c5vit1UL9EdO8gzEXgffp5189CdcD+BVLIrB8QVwPIsWQ2w
6z2jEye9G22J34s5kyLWPXnfXRuAcZQQrEz05MvHQGQxUsWIasyhERtMl7ymAwLAd4vMJ2X0D04T
oMSyjWeY+1+SDMV0bupkGREWL89Yuu7/ICqbSkcbKuQxrQcggnHRcP9ZN4AObAr6Q1qtWTPRc9Jc
dOImLsLmwSvgyxhyQTNKpYlLIF2LP3XWOBvTpSIP12JWvwzhmU+rUb3VZYItMMqdDq2MBUz9zYHz
5FsLNqKz0atTFNp2gpU/wxBCSL6MbHsdJvqOgfqxxiFi1oHIKH0IX3PSA0KqT4eBhih6fYmiUadb
xHAIx7mRNWd6lR4ZZKxkDfnk4zWXCP+YpOXYQEYIuUHv3Hw40w2ER5sYyHweK4hLLFGE+phv8pe2
jcaLrGZ9NcTyZC/XoRnG50PYgTJ+iqLDkVZI5NGC/jtESxL8/y74BJRovN/EfPgr06tEHYDnttM9
PFIpWpTsRqf99EWnXfXZROlKOLu7rvQse1Lj4VLxpgF/0q+FWOn6BwltWXcVXm6U4Ytr/QIWU77l
eY8FxCVx1jW6RTqskfOqxCkYeRrbwDEPsqiJuwOrbH5F8yrLjXyMZYfk5rSn8EVPUdse8jQBRyYh
chV/6PCR1ceQmApQ8U3Yz0kRR9pGprvwew5RqJxDvit2Y46RwjNAlcuHXk6soF5A+8zhG1OIa4bd
lmTuPtPtZe6ACx2hgR2OmMW4NJHFJZa+xlJiVg5U6L2M2/oEi/+490elY5rkgThphhcloCDxtsqU
meog1gt2RigbueR51hit1K1olbC3MQeYftMw5SyOqqiLvJFy7qhJZNNF6HF/W3DjvVREDiZtadQf
O3toJM5OQ9pv6Bsk1DvWEUL/kGIxD59tHNsrXUdInGMz19SrNzH6JJx6E9rqaId3o7C0WvaP6VVn
DErM/84DdcYwNuBymDzCEM94SzRvg5axoJ7iyAvwdxA/pBYiAv+VX+Nz/h4lyQyVL4D/ZkwtgZua
n4NTeRUiX91+8KK1FAkdfazv5gginigrOceN04qwG6JAwyvuxhJS4A9d/7jDNGxoy3dzFQeBmA59
vrBJdifNQ7dBElDxwJfrjo2+chjhvO68raaoEJWa6yPKR1o2lTvIFmD4d9uhFuSv1NZ7fRO6sfEa
yXcY1T3f8KCwiIxt15KH1kPK44UzFfzbCNzcWie6iNikQS2nDFotn3Xj5/xMHwNQU6X+wxt6OX29
FjhxNM7FnLSVQaefmgdODT1PlsEb4Ofo9IREk81jmk2tIsQiOgUsc7gQr3gA3PKvbaHK/OtkI1u0
3W2Dmd7kXb/JfqPxGcfjBrvFB9mg6WYhWwQxX0/FomuK1Ym1pXUuownsTpdT/VI12iczMiml+flI
w2RJz4rYqkY2pefwXIBYdIsAkaNLauYL5MMr64hMeUbfy5a6ytIlGM0obt3J4mnWTu9mPXM4mmxt
gfTueGLI8kbICC/PkserrBccXnVwQQec7YzDgzbM7UCQp25ro2b2PuSVbgkqlCeKFr02yWo1mba1
MrrqQ9bZBm0LubdJryy8z/CK17X1XjjKrMpVtaH7A5zHlVh4ODlQvz0t+uyhcqJbVzRLp71+YNgr
i7Ar680xQ45fKlANuDsH6BwDEN6RPrinH2swj4No+ElKv2TmvYTubEZgBNWvdejw5ihlJeIlWkCX
6ZohbqHwjoP665qSfUoHiHiRKMha6b9SCtfIajnFPokM1+dw73dhCajD0S4tdAZiPeuIlb1N7eSJ
M8haNvAvOL8mEFC0/WB9uhBh12ct41f6PRZYLtFLWSKyhDpd9ss41MQ6BpZtJeJJrL/TJcVTVRV9
A9Mmg0bCgp5ucUA3YNgNBTSSO6h+CqSmnzW4QUcUs+L2xcmFCEp4FouJvpGUJa5EMbMkgWCCgkpb
5ddF17iL2DXkUpEn1H/IjVIL2J8St5aD/WDVsuMTtSeecY1c9GMmdJjcFVxDHD00/7UN7t8Irabo
osy/b9B5cZ4a5PuMaGbHP0bvQeLNiDy40G/MT+qyGzYMybD+XM/3lWhQqIwzNJCaO7eWm9ZEXrFk
TXuh72AodVzp8XxXZKn+NL1QsUYWs5xLG/VdtBk7uNCEE6l7VXqjvrGsEHhFPbqS1LbduVVBY520
Cjn/mryz+6zdjQqEZOp3x+iVwZZWHb7Xs6WvL5ixg5XpE8on9KieommeQmBNbqBq+bbVmYltbJ+u
nXx+eqsiqW45Wv2eQcwXn4XfZ1IZ6Bp2gKiFIg3D3YR17qLR/rByTqm0+2kMMaRfb5n9GoW1I1TA
z5ReWgytzYFtqltmpMMlrWgz9tU2lNbICBAFTiNTc9e9/Ot5kBDpRtV+OV9XxvugMvujjiYDdyyD
Cz07CH+9WYp03OLglJPvJeR9UYSq04mjyItz+evbcTeGe+kyh8SjvlI4B83fRauABlHwY4MSeVcP
P+KGGKePHWQdLzG+mFL5KkSbMYux/wfB0DvFkMzK2HzdUjeGUvtyf/6jtpgbdJnKrqB/UiNt1gPQ
1muC+NTkBPJkTjARsWq/BUkarpMLPXb3bghtIv/u1yiGMcATczBqO73yIXj+I87i+aBI6rnd6993
puySBvW9VE5s/q74DQJzkD0NQhejkjmJoRg1f/ycvm/4Ilch2P5W/nChtMzxK216vaXGQoxi2OWO
5xNsU1gjqBTImLzFSaV7s6S/tD9y2LgEvcoayAxhAkk1tzV3C+Zp90ELEfmVcI/+zmXnr+3FDDr6
fWMQs5JuRCKQvb+zDCalKYI3/r3UZonlfPk/oayOk5xkNYL/0EwaiYdGjgTJZdKHCck0Af8u7qNP
W0A1vMEwWXcnfCh0O3RMsJWuSntbCvWSUgnG2DHe1GfjwfZ6JV+L+6TlKJqW75QjoMj4MZEcOJnk
vTzwLVlS/6Hsw9zzJJNUQNShfnWaCyBizOi75EM/wW+wN2B+tp/uqMU9YoJYGGdOou1jVdPIcQB7
9NkbpvfNeBzBnIykXdolBy/IwadOaOr4MTLtjpEn8CiMZf+NQ0A07oxY74wq/lOt9W5GfqmAV+W4
/emdy0+Cbv+C73TMPQbk0UlGPPyHhf7NnLB3T+ONKCU2Am2Yz4D0ZNmi7HTRkuaVEEAZQGzSXY0B
tsavCTx7miwF61HWyrL/D6fnpprL5bo0l+eJtmB9Lqvq7ErCqNZxHW8ZZnp56sBWj3LzGjb8on3Q
sfVmkEjZYxsd+fMvnoiByGLTgnM1KMFXvm2/8SwcjENC3eoNcpcygmkdj+AWa3DGvS85auCvqCmw
QxtQ112E5VUZyWe1NG9tUQgqVnXkzf7p9nlrmjxyRPJxcepcoQtWh9dN3jOozz93nLl3A86hI8Df
KADZ9V6pz2kPQNBKBzdpW4+O8uegWmIz5d9rxSs/E1aRlgv3oqJfEce4Ah0IYwHXsuWuV3MaoFPm
0nSi5YWT/VupcJQ/wbbTR1Jhy19JBL7gkKeOsIQy1SaCNcz2PitVtqpwXwut63V6qKIlLO62boWt
/N70F0KOtV0JE4dWEczkzpPDVcCs7A/+wPRZhCjtB0Q4JCFXiwbusZZYa29jX7R9Kbf8OGjVti/c
izt4RSkVgvCfRRUbF6XxSopVJZmotk6ZwHIFYLH6wI4/4EV9lAxyDYbC4VJieGPCq177Kbkb73sx
B90Nx6fR9e2D/vAD+CgQXwJ7pqUQhrVT/78eZjknNh+LAX9dFDYp2OojayyBm9k2pmIBdETrvlKS
2m+U+kS4DQUOvYrAWwcOwuO0mB6cuk1kGqYPfx5IWqojtuujAJfx/T5Zwvb1VPlF4zQKxPhot1vS
e7VI/3WVBL+J530jpMI22MD91TKoCriWAw9pUOQ+jvPainiQDt4HfvOfkGikFjLHLuPGrHejEqGR
aGKVXH5/BgVF+nY/aFDOnJhI4m9a3/Cc1idjviYTSTr3DITHiaGNxUO5BGT73cf25f8Oay+IaNxY
FM920JQSz+4HBiMftkpyPiK1I3cspDgtH85AClM2UTkZsC0Yprs2caQv+667edaLZZ0gaqCuilKP
Ig9tWV9mpg3BuUe2O9I/s4iCk3LzxT+RtSHmBsHetKcDvmmDG7kG5j+oyNlhZ1eYxV1LX7dxR9z4
cc5Db9L7U9WoVL91xtVF3y+BAkmsTXcdRGgaIvloRBAszl4fsBURClxwg22dl/+HhS+B5WAC4yDw
RPykVlUoC+21AiA7Uup72KiobUc6zNJMTDHergty+cnNRJUNhQcKCJEyCDz9hYliikfxa90VtJCB
3IoSQg/pl9XgweF4HftRrNB0mTG+WsTddkT/yM6lAWLwuyKlvZEUL+H8A7pAFOjWHmvsxVKVVPJW
F+XkDIy7DUcoB3Oyf6DHrUXOHMNLUEPNKZrGNQWQVf2xyJlw3BFmqNwM/otDdwnZy5Eo6osdmHL1
agiWDvSN+mNcsW2RS+14Mikpe0zmjN9lVc7Qgo0Q1FPDigVjgOHsL8STxDs4NtdPRfiCbiOZmXJb
19FAGI3iXNzRvxUHU/V01gjhjciB5lJRv/Lyx43J4pzBneInA3eDxf4I7N5ULY/k/rdiFSLpqQRF
wSeLd/rcmBj9iAN0IZjO2jWcrJbiLFHeJ4FZLRqlnpESJ9lhRDzMGM/QO3THslRr03Wz2cSp16GO
MdOqW+KT0r/cYLZTnxfvQEnqHM6Q9ULBvSsJ2rJPRTqksTLGQi53oDWQNFHoim5BwrbGwi82aQEu
A/0rT6yj17CdM+PnhPL2qFWVOeCwdIvMmr5sCw44u4rtEGwQsXPS6P+bF6PSeLxw+kBsCX8/st3s
bEbR0nv7+QfzGCe1wQvp4790tMUHhrPV2xkKJAk4H2D3qCY/CzxNSDSCvwb40MURsToQS5yoTBW/
ksZ2TbOgs8HUvtN9GwBsOt4gdVDbfmv3dQqAVF7fg0TUjb0YHXrnvGUD6DXmtEgeizdA1F/6yQ9w
KhZ7QntC43nTw5H8sl5QQMkV15JwhUQ0cxaMtWG14E8enEZ6gX3XcYZoyWQoUvvqsnomAr8tobOZ
bpU3Xu/mgBPxdl33D/kieso1kEdxrL6vo/Hn5q290oqnsvcDtBN6NoRnTEbXcLnOTAfIOhn8aAiU
nUmUD5xpqC1kvUgQytqCyPtKPqv4GT1HGfwuijdzh6ksNY2bCGtJnhJH0OC3Z9FaEpcRAPDJn2k4
01CJQV2esNo7NOqOP+aOM1NUO2BSKQiWQYLRY6W37gcMFRXxfeCG9z+WeBUoSxnSmWNIb4fHtzDn
K421Fc8+RJOmJS+inD6Y0C4kRfnMJ9RKLOGoRH+4RYz7DKdHu5x1wxAVfchEF1Q+RmDc21jmQq4w
nQm26OzWqDENa/LnP0nQtCSJ3SLPRuH9ntx4w9tHZiKpYWqxwv2Wm01GEEr1ZbEf174+m41rpZuh
Xk/gqhtT8kwsbhN70ToqMFOOiIE3eeLsk+lnakLbWNttFH1e1+UMyJtDbSRg721wkJiv1EpOqapF
0XnUjsNIMqBK8IAyA9tuts1Py3Ig8o2glWIb1JDUeCOCOC3c8WdnsYBH03cEUqZVK0o1LhxH0xOt
WOLXM8FyFwNQg5VmivTakZIyDNXwLUN0Ie82YNRF3jXSmvamrzpc42zO9RXbR9AcRxaZrB3v4jhq
G06+ImM89Rbh0QXc7ctAE04y40DYLC1sv6lmmOGE6W1PJtGio+T5x+IRjXdXlfx2ALUy/wnUaAP0
I/e+09MCSYr47bk8t0yTWRMVHEfIW4sQtKBNhogjIlpJC9vbGDdWhSyW4lUxC6NvMsCg2YnZbJaU
C7hDT+J/G3UaK25GOgzT5MWVI3NuGHJXInNPwGwJuRIH7KSl9nFVXSbPcBi6FVTHqk+RcD/IUq7l
Ut30YxphGasQuqvb7pwP43KkB7A1MO3a2U6x+0JhCUvxddHjPD9uos8l7iVFGkuR39l+iWdgXO/p
zfQ5zK+VFR0AOLKkRbFemqs3FRq7+R9hP8338bq3NU2jTXVB7qgjfsIlCip87eDC0AwYtEMdheCP
Sf7JqEdm3RCNQmNoviIfLeA6YKnaPuNbr4RdEzmHtBtBfEh+ONUgJQexUqysfnrO/N+gB37Ts5c9
7Mt9KkED6MveN75J5BSkRC+RN9jaunkF4e+DI6T3RkMf0QiYMfjcI/tvT9lygsp+RB3zfFyJwM08
bULzOfS95XZSioI22G1h7xfM36UKLRJApMMGvGQriPtFYbHiauWrP4choe9XadHFtUsVrw98FBsa
nrXtsiUIZIkuiq63V54pgfjaT7dOzFQ3Tka4VhCcF/KFyotqfhMGdR+aC+F86+7VKaZ6vxheW0v3
DpsNbAhbTB8y9njhZmO2Pfee0bA9VI/tXawuwN/IGfvzXGEruSYR4RmG7RALtc0wJi+ZtSHdjydl
JpOMjH4ipO7eb5iQBZSD5H89mQA1J59dRC3tPC/z4LVt2PPFVE1AM9HB3HNJ9oasJxionwYC2p/p
ur2+/0GJTarXrfJ7zAxu6U5TmYXW8bR9AyUuhNXsz33u5Vc4/OC0tyYy6jXDGkpe3qgOVImO6tma
rinXhgsZ98se+nj58BB8ERPjOKHQUlw/2JERQWTTbuxVMlezN1sS/x7mTio2ry840kBJ3GwNZKbV
72Ywjyh1sjti6bR/L98lSen8/bMwrp6btJ1vC8D6saD8VaKlIzkITU52XU+7PWQT/nMOPobk+tD1
DW4fjwYIzEbVVLv3i/D3jWTvrODUoFVwOoABPBvrg6VszKKDvt6VX0CxhZNQ8CbylHulNuKy4sU8
MBck5GD4i/wzfh3a/7GFmRfs/pc/g5mNfvRMAfyAnN5Wpcfrs3+6edCkb9c3RXRsyn2hcGDG0zgU
vzbNK3qR5GB91JawbKUoWN7yO+39oWbqJkvc9zdSfHTsYCSkCH189GeyJJe7Wv0zp3YEzQeWyAHx
0lqJihHkrQBaGjelStRMHNMAZTCfGI6ZUmHfT7hxBC0EdcwCf2rjBZJebMuFVu7ahIoCivWQr+0E
AWqXwV51iokSXne94R12CFMddfvb9Kn8GsAjNXhwEYUOF8g4tF3NczJL9CUBdGBAfgzqQ8oVktRF
Mvj6zba2Mkau83t2staNr1iuwuLPNjCSq2vbeoZrro1dkSiLZOgyyRegLIW3DPFH6UgfoA1QaDVO
xMzBP2SKe9Lph+h+U22m8iUMVZ/7Up56xeDrMM9tCdliTiO++sgkntnYVvU7iTq7+UzCZ+jxiEWq
O0fb85ZrbM5mfZg6JExnvjv9LzLMSPa7R+ZIzSqZq4fCSmgxR91LANtVMbbMJctI5hnZgqsA/ecK
I1dCRqERWgR+9nfb934soF4ADakxcYnpYrZqC0hA8VEvTVGf4LpByMOWGp4Ulttwk0oaG88Us/N0
fUd/Ckj34WgH4c6mteXyoaWMu+dLhNRcchN4R6nEgnFW8IX4cMyo7QYON+fa2MpBkyR/7KJP06+P
3PXBao35dRIuWYqCOSR6qeQvmASBBS1bBSjhcbMh/+gJTcDrymmqVlqVV6Ab7X2PF8RbEeRYx8qQ
KHQY57aRsLszxozXfhbb5GH2f3NJ2rlygcg1YyXO6Vi25BFDaZo0M5m6NxsmfPtTurl+tLU1pVHN
MwYtr1UPJ+5corvLZP+yKVvXBmkM4svzaYSc90oXsjUuOwftogDy+bCr49v64Q5rJ7Ld0TUtxwcf
9uNxc10m0Kdc6uMPospdKwTbJTUJYPk5EpQLh9XUDsDkCaCmtgUQoxN81Qnvp0FryyLnqtiEjogx
tfQuqEPIewRe3AJ29dIyYIvuDotmZtjjBIZ6ySqEOZVZZQyEUK1dictbU9ZlKj4xsXUONqteXz4a
yUIZiPiMXqI33lm8wi4+EbHRCXCeP0L8EIVISeZnYND9unYf0Se4u0afANFyHTZSK9oLTTdj9oJE
pKEobBErAjP44d2qTj7QgMO/e0Dg8buy2iSRFRZyKd4iMtAh1j/QKeQWKdLm7rinNNGlfvLH4KUV
zSqBDD/26sFQoAuINEkRGhH7QrhUI/6ptFOVBUxTYModjoB26pGJZjvUj1rNSksXe+1Z79VWbC1j
QiQU8h7cs88LJbjTf0CrFpd4+cUMnJ+6L2/VQ0aUhjK6SppmlMETEN6+gk7YEnU5qb2xxwZm2j+y
Ys08FUtXvqXrqPRw1Mn6m6FOT3E0QwID0HnzWynNWQswaCWMsd8cAQLjlTxXOZ1skeKGMZkf9Q01
FBuptPs50RmLP3SfMxfLCheFPv9peEyGIUKFygwxjPBBBnurFWIQXlhZHn0FiMiIg7c5gyV7IB2e
GxIcXeoho95DFBEYoG7MIh8lY5p7ZRHyHgQ8VcGzGOCPck5ISm0AmP/n5/dcJ+guyxF8gp2F1Dhj
KDJ086ldmSzWSFfePG1GJ8PeYuabp/yL4nw10sz5E2/1Z6Kda5mPli9IbkhuoE7OXR/T5YFRfwFX
4K1Mp03u6SuoIWICYIJNmGYK+u03fsJF8mJI+CCy0dXhhKqMaWi+0TTKyblzRF3n0dA0haT9T0E8
l7HvGGNTiw6BccIb1482J3WvlEbmTqexAyEQafZSXKSLzQoiXWdYPmtunruwxjQ3CdrE63M729rt
dhV9Mw5OwG1OTmZ34F026ev2lN6haqteafwSvmf8n17RvGr2Zk3E0CHN/ksLDsqUgNfTxMcrXQHF
YOlSN6s0VKaW4wZFiRyJOYVxlXa4Z6AFChZfECAw2VWjEJrEkD97e0fZipg/vP1US5irTzmGdSE9
1rtsiMIXlKK+lwC+wzVDAHQxNQpXDrGsqHv4UBoSXcJEaULhakdKQuYJ4fKKm0PHIwMecmlWueWv
upDBMQd7gv2BwDIrYcvHWqVSCh1dkXUiLlxxhS8o7kGOiYP6mD7Xt34m6heb+4zEIq6o5hQtMS0z
lYuklyZUlVCpksP8Ave4dSfMTPN9kyTN9til1x84Cy/mNeqCnaJpZNkc7JRzcfW4RisBIE4im6S9
7kQSrGRIrd21Zkpq915SpomNtJ4tdMZHmp9XC7ipkMPlC+zrWYpqK3UivSaxcZatOv6fAvTjgmAN
a1kPbN2DKmAOkzfRrAThiOSc+uu/j/+NmwzCk4bUlWScJ7W68zD1blcxNWUmvYTxZevaed8HwBqY
fhYPQCfuhOPX8MNOoqmzcyxyraWXuONJC+16VR9K/K16x4XUyV95pqMz+PVbyNvXghsWXn4vclNs
DWmcyPTV5gktcx224L+TYPuOnEQkljOSD14EkcWtL5NclaurOU8GvknhU7DfehM24ckYbFy8s8VJ
zTBHzccGqJufU3iNum8RwCrhTQH0OyxszFhDBnsDP18ypqTbZzDty/mkDDizKAi0x7DesrgG0T9/
/vn3G/yCOWcTKk9YW3fHIg7SDQSUW+kWMGu1qDRKVYAYD5ZskZ5u/7LQyy/hkB9GRxOVIy+FeNQK
5NpjjQwrcSG5cVy/xgVke3VZWKBYQCpOLz76aTr7lXAliXXO5pSFojyFGSEY+o+zcEVXL3Cr48aJ
oUvucH8FPWZiZzsvGyujpTqFvdhtYVtsa++uF8yeW+MAKY5T/JMimuE2I58JdYZJiCN/c2Xbvhwv
ijBkw6zukfmenqO9U/WrhCoggrecYtQa/YY65hxR5HH0lZbOB8O6ihCCuBNwJOM8w7U82vSP4eTA
g6aJCRMuuqAZHN3Zning7u7/c3iOoaHf+ToVkq189rf1jolKExeHdN8o+a1B0dsrKBvJbTqLGw0W
/b6JYhQd3CxRn+tzu73ez7JYSfi8hrsmLSM2MBVTy9OJvJeR6I3lia3bCLVqM5feHZHX/+0gr1hs
v74yh6+OjXzDeF9cwpMwAhmqF8LQWxp4bF8PkiNsOPlsAGciWPE4tskUa1ZKtnJ4DS/I5Md7g04E
tbctTURpce6G0qP9yS2y6BghnJKwHARenBmMxq4fViIN3PaOckLzxU6Mw5iBlIpI3iNUuKVMxjhq
Ov93ccrLwf3m56Z2IFKN2+qPxZJDfQOefWk3hXH1+L4El7uuHyzUpbW5yYbrlwHJHpULo901/AeP
ox9uOYV6wNRxD7XGy2CYWD/7mgP70/u8towxgoPrvcAAm7ML4IbDF8P7KA/FLEONkVhjoyWfWDEx
g1UT8d7EtfnENqZkLAGf6Ipq33JEjS8h+i+6gHs2er+nTkg4E/bZn0psERIZdewjWH9c5OcbHiWv
aEmaxa81qXrsFwUuXY9gU/C0lqy8ORuhUeus155dH6TiLRNoB9+pwoTMlWmBYkjxoxsGjISgnNiO
9FZ3V1iBkCf5ba47A3XT/UZrBT9ugbIgO9p3Jeuqwy7Q4rm43sxaLsU6By78cOce5IkoaxDa/NlR
qnjtEeh3agw9PtPqoj1HTNzegvHyG39K/TlZWvoc3Ifzct1BVfp3wXrn3BjnEpZwRxzF6e+SuFkI
IkhejTPYk48JbrBAVfuNYaEZ4blKsawVYwpI90W70D29pCVZSFkRQp/ETsu1FJalKu8h6qj6ecj0
Tf9+W1dBadhl+DGE9HXgEToddeWN8teAu1TVZ6WLsRUJ9ld5h+v/bBdwd6u6hR1XgC2HtayaL19J
EtVQnqnEvYFyipE3q7QHmQhNkCOAQBsYYvaE9Up89JR/PsdWidJkjK5ZGKgQ//anUlGGRq58tspW
ygVSiLSdCTZZ0cobpw7AF/YHoZDR0uj7/i5lKM1VOgCzy8eWU1HlxpQkpsvFdOy0LZu5cpPrLur6
lWLhICOVhf5XFS5MEaPn77itYPSqWlULV0/1XETfLdArNSm6H3qd8CcB9BHZNcW6pLqIYL1Bk2Eu
n1PFi4uvU9GQ1+MveTLDtpLmPX36sD9do8yWLMJku7cfYwUYNntdcF6BROkzQLpKAIXJF7NKGVoo
cAWiDXdo5Popz5HHjQhMuvMfIh4vBjbWP5q5ud/T3a/4MiXRetAgtRjK6CXIOwcePqHmp6UlJ7+f
omcTDqo1vmadDj+/SYJVbyRQ5GKKcET66q0Qo0VVz6nk/zu8bglwK62cHefa1dCl3zm2MF/zd3fA
ExsJCZCaZyqJTeJPSp+Es8iwC2LJ2Rnzhhsp0Il6XYISHkG5cmcRT+16kr6VF1YrRZJe8UqyvbMY
u8wvAKA4c8Igsk4wEMFUn15KXg4H4SJaDk30kTXPtyLSy6w0b0zNwIKfr0rnMdbd2aKCsTCG6KVr
Ea7ftOE5Rb7YhU31uQbTP0CHZXOIPga9ha+TrppltfqXLW2cdyATxvvTvTdhPn/cLU3zBq/h3vT7
P6397ra+zyG1KKMDEVjykE0G25990vlwWWPbIJjlDQEKuVhjRgNioWZTAlmQYa3MCYq7RjCvUIqq
Wu3EHcoZYAnItfcXv/oReVnR77eVrVX+gkab1O8CmWXVavfG6evvm0vvYLGUfA2CJIkoAVorJjQR
b2nHIpnFaNfkj1AqYcgKPfzK4okKne3nO8Ljs4IV+jvPyuG64zJ0fODF0G8m3etngvT6UohbAjDW
O4d8OTHS18XzfKEMR2vRCNxtOxF4q7LS8XJsbBFIt0y9setpFgqLlu0N8Z+Tk4hT9+StLDrNq/U4
PkN8HX4O/U6jh4DzyP1GkcNGh1JxArZEELYEp5Czu8kbRwyK4Nomnd7ye4eOnhL6r0F/QfjPUnup
sTna8lkUPKpHf3XMjUiTJMQ1UrMJPtDUfDtGGVEYhVd2o85RJ1gHLvznyf0xq6YcMzsw26vSidvM
uKnCz4o7BiMXwtbHnOSgkmgmK3lvDb2HHhJneb7hFqkKDgVTlDVKmiX9XEqL83biuY9QM786iNN4
GfoJ6Ua2SPXMYKlIVCiW6K3txnKkozRQhX+EVNzRjt/ds6sGsoKASS1x91LEAcdUC8emhOuc9xP2
pegEQp7ig0X3FGQyQXHrR/ynYiPcvZHUgyizzt+OHxYHeqN5xCEt7vC0CAt4UGWHhL9zQlwo+xiU
Wf6f0k+YFV+LbrO/JzU/nxd0lkZA9e5+X1qk1M11z6QA2Bkxdofo2JcfB6xi60AFjbehTDQPv5F9
jA7oYNgzR/gVCy3Ak8KeQtC6Gs67AoS/6JY3rScC6i9KnzV/4A9zDG7VTdWSkJmqafcJA7Zu1FJL
DagdIgfioOI55hJra8DiE1JLky0ssaFkNzR1CW4K+Bn4WTpsrY+mexAekU+P02dkqX1ARQvgEkz+
XqUvvTSqdyGhr9UYDu9E6b5qawAVkvwbrx7GU360D1145b8FxojZkVivrbEt4pkwDe5beCKexLfy
SPVAcGmG0iSdcXdHem69vtlj78hf4BwHNhr5a/Jlg5kMnoeRjP01mwSHhwn7DRU48sC39Qe1Bzs5
pgvCv/THCA6qJ0kfTz53lrFRAYqi7eYEdi8x82uUoJp+vBL1dPZa+Vh9KBvU7y1iipww5dAi2ELe
+qTOftvpmQXSA0QgpwtDzwxFnPx8Kdx6wPP+8/FtjrpFqk98XhujTfH6t+ZAdxf56xKXu6/X5Zai
ikbh/LGYJ2LaIFw5ZojmmTJWSJYvj1gHSd5yN6nsiYDnTYTs1u3DRsIqs8zCuvK5X0y8cpiDqgmL
ksXPRYwLLsbmoZLPCvhaq5qxhIAP4T/PV5ZbLgi9E2aQRQdLlVhtlO40NikLlIExQWtqjn+2TgIh
1AlXWVu0QtnjmVAvA0W9sT+LQRiQpv42GPjZtIZcxgkrwjkVM2VztGfyF+qot4DV5QEVqyNjSsCn
b4XjWdB6AVuePt8pHVSZa+g9M3Dlhh2WNb+CI/rXgQzWBk0LtaHNSap7KAg1x9DWUAJIPNfEjEtr
bO6AiqiPAC4znXspsCel3tvpNvmjqGc8QUeAZ/2hO+kW9eQ1tK7UA1kHtIIafO+PbN3pR/8gRpH+
J85KG3zZFy3OnOxU/boGUBS55cPvcF6AmNAXTQjrCrR75dQr+vFaEYvMEwS+Xj0nW8w9HJsXfIrO
eRvdpeL8OD9XJwvb6r03niZu6g44fpPI6tJFjPn6mk59V+DoI7k4hL+moPM6ucE29dQ9pZoRqvN8
SSzOA6yBiNw45XeYYqhq4kQv+dYg/UWwZO0eydAwkDLDkchlQSkPLf5qtfhdX/XM+PTswtV2O+QS
QAl6LuDWbGpDqSdu5MyYdEXn4nGD+GWOw0UqAqjWWCnIVY8zJHPBoIpLTjcXj5wYiWpAbjnKkRRz
brdiV47rhgEeWPZCdQGQOwm2zYZuFyPcqV0SgSamE8+Z6KHILfzWuEDZyxsqA2JBbiFg3+ub5SnW
+BOFGZ4SuLj5A5Xx9aGaBBEmbsyBDx/awh4sy3bxRL0X/aEvlgDKo71EPgVj8ybx2QrHeqwT1tzV
W8CV+Tn60Y5x1Cp9TotkxDIE6+Ykdr1g+vFHQI7I67TP4vbY9FvGtAR9US5koKkqdiyADqjA6F4e
vw26DWMuqM8cGJ8QH5koaSNdmKueTri1+Zcs3vkOSN5UMn/onzOkN6TTPVovtd82JU4/uy0Z5x+q
cbD/C3ivE/UVMJuVmd7DS4lGVIKa8A7ZsgjK3lYWUpjiAaIA3RESHZ6h1w/5WlDujN+VRuleg2J0
O1KYq73f3OdHxasRNaZNimRjDL33gDS/7kBxzE87UWAEIQwPIn4L8yhEBpLPxefCoeJ0JvM32mt2
W7an+8MIGFlEi1JhuK8g/E9/aOKC0nMVnQo+JMZPQs5NvPPVmHBNKTTMuHVKGcBFrIY8XROhGFkP
toSzYZ4N0HMbGJMiYVjLydn2u0UmJRYINR4fvN6G/EWVwGMMxvg9SCfGRPbLCklSlv0IW+eyAPCJ
Uo/ZW6lYUSD+3syG+e+xZ1U989mIxaUqtJUTifmzbTSFUap+Yg4G9/ewLm1F3kB2StnBDEePUsNA
T+U2EqNeb16WdDHJ2aVRDydxJfj7vZ6MRnpCBsnkS0KyujimCV1r+6e6fSqolv8P/p7Zg39LTZFA
5A5fZF6EH/cw/0oB7cPkiA7dFSxCYxTn7rLd703dKpuNi1LBjpgVp/l5j+jrO+kWveknlF2hI1Zq
bVmy6ky6sssPaJJ3Fe2/ZtlkutAjVTxlkx1dQ8Kdnrcpge+xHBNC0MjelQ1IvPiK7TopjuXS13jM
g3cPu0uO3nuSxAfUCBnmpSpNVSM6sD5+vGxtw8UbJ71z8PzaU4fCkIRse+zbI3D2HqwBusr/FghS
eduya1tKODPSh6NtkDN57j5TWqKP9JqEJySPxUict4rxvZwsck83L06oIJf8aX598E8UZbY0A5TP
J5UK1w0Yt9JSaZ5FBjuvOxqKFZQDBgNehxlWTLyE0V6j/rlAVvAljYtb8jXYaXk2u9p/khY68fs8
rN2gNidUukw1fHIgjo66MZKtyvp2loNvE3NzjQTT5BPRV8eyRKCIBQ7nqndEcRjt8g88PvmYkEAG
aWS0tu7TMEutckt18oaTdY9f+7I0ae9RtzGjsY6QcufTfjkStVGaVnydGDpJFcc/X5F8jYSRzEP4
3uEJm7xiiAZ+OGyTqyFVgJD1S8zZuygYPDt87Jna9lCtXKQ3IgqaE9a0qg8vJXfLDaZWauIuXGvS
mEhtjhB3qF16QkTWUBdTnaMidMKCP+4qLPstJJsmf2x1KSaIR10kEAhMSp8r+5jxs9PUHKvDvCcc
EntKLcei+EUg3VV/1k5ZNbCtkRVG8ULAziEC46uE0ELGFArarrWeLd/WfAjxmmKAkGpWJ9nsKYGA
Zyr7DdAP8EDu+Undk5VavJ72YPUHjrvQ7jSBqtpO7/wm5uHpLQJrZhEMidDTyhDDMtLvKkZ6V7qw
5yjEfZDoToIMHXNS76S6zsWXBLcg1Cd3WNHoQA8+SJ7qA7ArrOTDxQbNvjpqSNVB17B6tOpdjxyA
eYD3iadaYA+yzpaFDw3zM0zYXxke+O2+TMkyECs4uBfany3W9S5vp/I8oWHj08siL1oLLa8HX1gK
3yGayyCJwCsF5x8d2Aob4Nn9bTFuZR2e4I+/acW6bJy6fArfBzViBTJh6S6EbxDpUwkkuXnrqtls
vArBkvu4tNeiXOGhg2wq0JDJuUin5lcFdtmG1r+49dZBT/LJAN9LR4R++EQUwPC7fFExlvOmtJST
PieywMaJb9zA4CIedWhgGnFB/01N1u5yn7VvK0R4DwGAudoVuT4jMwUhkK61aWyYBDGvOOYczjJ5
dCRB4I2Sasp7xhT+cm1ETQeO6NOqL2w1WpidNpqHlkF8Is4FNzkSSBVHw+NKPzigBUxG/XeSARci
Bps99g6rI049sLNr+XOnjFqrbvDYL1ZGatP8gS3c1rlyMiHmf6+Txv6+BX10FIWNIAkZ6OpzK/Uc
RIzVpclgDJfr9ArDw7L6QmTGq7Gbuyx8+6SK8qhrJoGjsdOh+MJwMpWqv5p5CK3r9fpj0eR9p4NQ
fmLH00BSfGvMDK9SG5L0bgRmiQICIKGPPVwfrvi/0qw7UitfxfmESVZr+WhRGfDsUFTubJefre5R
kvokuV8lw3TRICJKLSik9ip5O3DGjaN4syIAP/t7H2L3eVzhFnrUPCLo2c78R2ZpBs/MqYiKP1fw
5s3m7Xj4yg9szoS1pKRK2jY/iyS/ebsE5tH9wd5LyEb4SFlV8N/eLv+Rn1Ab/WRF3LITaM7QEc35
sMo55FK8Bh3nFIqdQkdA7L9rBysN/HOQh0UQ29Teg77u6zp4d8VKdQwJ6VlZ4/bC9TRD4ZCDKSfv
b61PJA8pN9aniEfsc0DgWjgtjwkmua9mUbKWPO/1coe6U1KL5hOcB4rMvYWvBkiWZe38duBlaChQ
IsBwOgU0ihZf+zhIKBvu3eEQIWN/3ZDkhk/jqmG0ZcaayEE2H1DviiHPjB6X160QvleLh5e/uZOS
u64oF5pmDyLEOM5ulaOuRnaVNCOiQVa70sQ20IysYSzNCgS3SAg6o9oZRRCA80RWfPbICWfYW3St
XV4hLWHQ8g0vxTeJ0LdLJ40o4Io3uPM+EuHaNgnNgvNuRfz0PhgYhQCNtbYKt5xap2B5eWQknpu2
9XZbrf6/IBhdfYBlAVrYltRKQ4m4SGPLVBjjHQTat2B+9NwRZSDJ9lNKtjV7q3Dol6A6Joy9UXv3
zc5n6rWGBpMcM/0Kk3Mp24PxYBlUhaxaaMkVDJC1Vs7kK0+LWNiImTgEfqlGjl7bqnAxrPYEFIbY
7fVWHT0NeNKJL+4QvmKcR61sBLl1L3TEfrv+9hUSFuWTmgcb7YHvUaCTgFRJrOdhgUEQA1IgCgbr
trH+n4oPbGTD0vbwozb4R/LFv3+l+EiNuCw6kttXdPZVIlGQ5pm6iqxY7ksC5S1estgTX6Y8qQnp
26oGnNhY05LiEH7liEgUlPtDSmt188ANRo3/OQkTzMv2lNBPT4NPi2zi+ZoGiWgCk5OC4T/e441S
3x1Ycz8J5NWSRZC8mLD4zS3n2diHJ9hdN1GODsmPuvOjE9JHJ6OuX/++TE88fAKnp/dIc2Fv/S9S
BWloabZVhkNYK/sJLyLgjxjxzDOoyQjJHubtseBmUxNBx9bzkFeae2iuZ4Mw2wq5P2UBmPu3+V7h
vocnhbB1nFhKQTyOSHPB6Sgbs8Zy2LZhJoN/G+w/da39Kxaas8QLoQ/fE9hWIkdmhpg40AZJzz5q
Arza97FWm+e42vcewFo/pv2YSJF8YghyQgwCuQL282eON6bZ3lFqQw9rEY8hm04+zwneQZU1PSJg
i8aAEBbGvCtsEYE6s/xZed0rqdVUA5my9jqtK0ZHEo2G1jfKZ0oqW/Vw4gkw4oJASYWYADw1esYb
FZ5+YIT/uGdxzsDNxu1kRecKgLUIkqj4Rl93F8pRo06mliDj4wlWLWCsfgSR/LP+2VG21jAzvd9w
bgm7z4u83+0KXB0bZiU8MtRX9hPGpuAWkvmPck90nslCwT0VWnrc3NX7UlyaBsS5kzGXVZe8SF8g
D7L21tmaZUTpUrLP142jDwi3+8bcwH7PObG09z2bt5Vk6X0HhS5wSzJNqxntqERktYY5S3Dns9o2
prhW4is/Ge2zUTQIeQ7r1Bj9y1XxIAInyfm6mvZdSR+4fQR+4AP5Sd6mzrIG6CI4T2HJYZS55CqG
1mvWjvFPA1XhRDFY3G/+/ciddEWIYodpqlbhmIkB0A4XY1XKqDk4zB+QHWjTwU38TMS/CbxIc5ie
g0Jlyh1tWy2hfWxjEfENLVEOkKl5czwLVmdhGNd0/nv4gjSL/PGGLwh7vrwOUVH2a56FBKsigRBs
N1+pkECtQyGNU6tbWlLZXmNjlMrhVlyaM6IsI9zPUOqQyWqFvYlJjxW3oBZ6hqv8VgmTXbnxkV28
PxiFuXwtcg/N4i/FxcoDUSTeaPNxa9R3NsOoq+/AGT4q8gYcIYLM1a6n77CS/fmViPX3hX5mm2yz
G1EHGJqFSY2fYSuNMDdKDt1/cRL4SlUV34zEP6ficBNI0+uuH/69fsQUlEiiZTTSiMi46MpVf9Wn
9UOFG1vfUl0hx67bZVuiVImcSSBjgWkENDj8pVd0nQbLNGtFJDZZHSVjsTtHh6NaF28j42RA6Q/q
JYEO6qoL47+9vtVzaxs/QVwM+oefTqU6qBW5bCky28AjUWxazIVPbMHJFHuvriyFnRH0SR+xE0k5
V5CV+mfZfltE8xCHDvzvrvzs2+zA4UG1XXfu/8gDGfkroE2b7E9FQTX7S6fMmFEIwKzHigbD0+8z
jn4h0Q74FywhGLpY2V8kwNcDXvIcM+CmS7pd4YQyMLKb3+FuLKo6hjYrolcKd0dr2MpWWiJEmrk1
F08GBLiBxRu/2aymq2myQaP+iXGrs7HOo8bhaTIiFY7OeyCN7MMXMoTqPT/H+XT+SQjnAIp8tbHp
LFI8BkZ6qXC+Af61m07wAOTyWR4k7GevW3FZb5TKIWx/sYWNzl8kOzFDinpW+jVkIwnZPq6fJQBr
5JUEqycvx4i8m0HiQqmz6B+m6xcn9XLL3M1PGTBOA6pPknQY+twjuFsV46gSZdSmDVdzT8y7iUmq
SAOecjLPr2yzBooUAEvQaFAe/x/wmBK9vetoA5mzyFmZyeP0tL1csL2eKsFNuuMohnyn5nr7PliE
c9MFO07pU5IWlZyxcHdSlCuQRST3FSbfaComvzggdF0Ku+nj1pNGLapBTVjGyAWnMcIkXhsviVYU
TY8Nt1fevEB02OorWCtAFgP28nZQ0Pxz+NABd3NqiI7y0Daz9+lr570oI29A3pAJgzdd6vId3dXt
fhO/HPLemFi0MItWrnihh7u4PH+PtXnhWw4BIj6zFMkVroYx0zS4e/bPuHvBk36BWT9pp+uW/+Br
95m+jDMDllUOi8Te6VHtdSqcnvM4W46G7X3Zrr0g3b4JP5JJk13zcmkZGtpHdwN375IMjyCBh3+w
hLx1uRsCFjN+aqa5ImTdKXyzq8pdSR6PtHOrLO2uTfyA/NYYHmwCAM2aMT4MXKBLATk8tvFyF3q4
5jY/O/G906CPIQ0ap1KNsElkMUtJl7jVJcvP7IvWacTMnixtDqWbSPQ6y4TywX+/fc1ntWnm2K3M
fOPHS/qBmAyfkggRsIU1SiuQFAu6lawKQaWiaHrytK+x1JVJKDW8DvIiIKopqdjCZPialncguDB5
3KthhZibZ2NghXPWLaVB1nxGYheIRfzvviU78MUeuGzk1Il2GT4P3yXepO9AtOkFwKSRd26RpuZb
MeXgHZuzfnOoKz79QmVsFRuHiWywNntRvOG4Lj9UU4YliEtKUFJID6Up/CyBdgLnsVdabH0MQTQ3
c7YiOMI+Uskmd3BTlMkFJNjSCOIIkLJn85NiA4cTeSb1sdidwVzJ5c4BJqKnfTS+477lyJdTF1UC
9eCYLX67TGyTdBGKK8gE3h4MoiKxLGpOZ8YjiJ6EuQzomfyTK3WcdZJygQRRfA+xn1fF7orRMuSO
4fHCSemMZJX1Fd5hyb7r9OxBj+jfNpoCAqYAoYUWoMR0W4NF1Ns61P8MrY1MhzTjqQvN6Kd/qR+i
AY6um7tAd62a7JJTl9yNIWVMYfrXh4rys5+OBU4Zt5nfjw+7RYYspf+NHvMd0WlBEuu1ELAgz70Y
SxB8lQGCdrUxmeUe+T5ewCsFwzb2fqJoSEAfliOo+7LpZ2YaWrXh9fFUgsiTZ409LNClvWK/qvSy
t0Tzm+T+ueyffAW7Px03z5uF5Fn0pvWvkcv/mhL9+zMw6yGC2XEP4lE8cyH5sA6CdQL4Fq8QUakN
DOejneqIsZqFfL2OULSu95IQOaDFhnwNiRXxq+vmZXVF3TLphn8MnxnH16AdXBhhddxeWSNvZJSE
ZfLzSls1yHn43ejV/GMffBzpvHBqtBRqgTjxgW9BfKmrBJXLGUQwtAxjl8BF35SMuFm1CZF3iLYC
LYt+Y8lIIGEQY+d0r1qcQd/u9fTHz/bnFdA3+g6J+m6Q1dQKd8aojFOyJQeTECDQ0aO/A2c9OUCJ
5AckpnpCFmsqJEWwQeHON80JwfOHaF8yZ8k8V7bc2qXjAgnEOlxiQ/lvPUzDpOdxfUIeoYEQAfKK
Q+LUmYdBMn59UruNUQLTts0hkdRAq6PXHk5CSXoB7pJbyrxGfz+3+8x69UKFJB1DIOIlpGSzNl+A
sFQwoeodx+6q5XJ5CBTZBJpLaklWiNTnHY5h3ioc0FnjAJszIR+XNaSzoe1sJqUHB75+feZQLeHu
D7SZ+s2GtVEG+zGrs8t6GfVKIelDkM11UDjGxe6XDQnYvgwLGbar5u1BAmP68iCe8iamnS5zbaiN
nGBn4jMKyzCdYNaTcnnPCGzm2+0xnXgoFMHoRPdpmy+GYOweeqyD+04hC8oMSP8sROgy3OzJxEMA
itI7dNtIX1NeLhdWv7HQ2iPXwQaedEVKlzN/yoJQz7/N3LDjB3Ew5zJ4I8cjPejeUcABjjg2CjQU
HtNbFFHbrEvwqwjjil103+m1Te3r/vKV1H1MrR7RXsl3saCMk8maoBSC4LvLTVmWLUvWHz1VxkkJ
EWM4LSse333XzfjsEogpK4amWWyM0/PRVUkSHYdboFFdmLe5jmCo3batMJe2yU6Y3SGR5EZ/0qGL
sUhVchLdIvVFflZnmYqMHHKj8bAr9W3LQ/XPy4CplBOV1qNBPa39bH34X0X3LHSTgz2CJZqPnbAy
rgljDidzJZjRoadMbEmWXN6a/Rc2hQyaJ9HJpO0veD1Ih8zyGqsF19LJ1BdHouFuO6pt7HgS2MMI
8QT/ekY9QWg28QKMsGSP7HIschd5+bMdyyfQoKYUuhniEOjXY+r2eq5uUeceReNrpdui7Pw8yNuD
W9LqyEwLwcqbEOnXqjUR21AJ0fID3C03SPdQN6qSy2TAjopgqV5QdFOC7sqJyo0kRQjh21RIVEjR
0od7NOuSmM5RGssrp3GrG0Nbh5Uzk/eHJKBmxQcy7aaeCVpI/W2E0Y9AQhbuOQ+joKb8twPO99ns
qpusg+PS0sEX+GTqMkEfT4RnAtlI2hXWnM6MsM76rs8qVSEQVXLyjs7UxTXanWn1RZgWYGyQqV4s
wJx7jP27iNOD3glaLJ21N0I+uHUBpac6C9OqO0DUHQtor1SLjqs2M7GedmyFCfhf6bS1EVrOKDQq
DMScMGctJ3K3laYGjf4Q+xryhyeZZhGjxJqU7vJCOkr+IJN1uSvai4TQ66YtJzMUZQ8XO7CCqnZq
3oskx0srMuMYT4j2HF8n0g7XiLZFe42XjM/KgcYgnDJueKsVSWp1watvD/N+Ipc1Q1yxJYlvt78i
fitUS04EODZ0nGqFRveBUpLmSXvrFl7tOqjCvBLo8PeRj940xv15rxcztVir/O8FvpJKEcmoQadN
tKQqenuEAhydwT34qtNwsVSbbTnzQcxWVB9NWl8fDstwTs25QD+CiYbam2Miy40pBVKpa54hssUs
6ZR8pYEoq4d8mBkX2pHRWjpmh57KHmNWCr8NubCjCiqJ41sGAGK4Qk1N1K8JIMKStPOjbl8y8TR5
1Uh28HMJ/np4NulT00LszRR/kEEmkUSKIjNfuFtKbx9SruuAZ94BQ5WkOkaxROdMN3JlKe290qOe
p2S1wqB4sZ8k+17s8uBUOvx9JyPu81si7Qv+T+gXGHD2DVantHB2I+LQugXUUxkaZwF5m16P7jZI
DgQxl0kHHMNj5p4GMHpwPzjQENxIZGakcqJhowPM9LKsbEKPMGtt64pdi749ejL/eaDkHXXJXBms
4RWnPoEb4wIa+CfUtarAzdSFgDZWeyfUS+GWH5hyuvqtSI/NfBKS4vAY6lfgD7eTqXuZsCeqlL/v
zLRI29thsF2+BqxIDOmFnvUPwoRRdlcuSx5BJzdGeovtvLoUNkcQxdxpLmmt758wR6IAXGp+I3BW
CQLLqfOXSsmNzL4OSfodGNSZH1KdGVO5dvODy6AVAH4Sg1EjFN/h4xGMIbnPABpJqv3eZCSH+M+I
cSDRxydSqh91VA276D7StMAFfVxTY4aYyosGb8VUhhf2Vgzd+XF+O8z/w/CN/zubnRR+HQvxp9zm
FMfj2q8PbMLpOA4LsJU4hNzzq1dwNssIGumOO0wVwRGPy7IPx+8JhZ+ipeJ8aHBftJ87egwQPyr0
820hTR50ulhtTwKPBEZOCU+Q7LNQw8D9LlUlGOPZLYtNuy0nkLuu06dMntLHjCNfme6eT1NRnBWW
9r1bI/7Klwwculp6QXPmlSGrR0pG+PYoW40loi37FApvVf+7Mnf6ux6BGU9ooOlPKCzGahHGGF1y
8/N7r40jpjA0BeoC8xE9tdc1Kc9iMMksqQjQ0pqnK2aK31fuGdMUzmVjGXMwpwy8Uw9yazPj0R+p
7NWYPKEqKpemhvXu5h7Rq19velpy1OPQzF5Qke9PZfEsl7h2Srz0laVW+lN7/KdIUkHkfUpcWR42
sgk24G2XzrGZluE55Q9/uyPk21T4RcnOXF1F2l7eQhio8XPu48ai2GvCvNcIo64ElHLh4x5eiS5I
FHgsvH5X7Ck8vTuyTDHjjj2oYsmZ3uRj6byCqoit0FRKEHrmck5v/55J6Z2TupgmSfsmjQobnePc
Y6vEcmhgyvVB3OEnrgIPJp5EPcNGYl5GQB7olrrRJ3BkIDHnsfNk2io0zYrxzvEPfDFi+rtis/ke
3kBAwqTS6o/HqszqtmC9fYPhLu4kkz4mxjgp5cubg7+Rdx7uk2jIMV2NNQhTyftBNmMZA6EgkjHA
/grHYzrz0AC9FRRrsna8jrFMomc/7+LZep9DgZSsr/IKc2aXxGaFYtm0t4TY/ArtzaNj/CWJGXRN
V6mmj/Gn7lSRj3YpYMUX3Wn+WaWtAqeSz98fN+tBsxmDKc5FvKlWggq7gzI60LiKtY7VupfrmqWi
ieLz371Z/Py5zmWrwEcF+RS9ZSkduTrn+QqKKbrDdwlfC/DijHbAbKjvmPATNwJKHsCV0QyXN7X8
XFVfno/40V2zxa0usQtj2Jh9vmVIMvq7RXQi8MoH2+EB96Mqhdap5YnYN4mpL2x37v1Z/JaISgRg
kXI2/zIUv2mGU5AVQiMP4y5oUSmLC8ebicB8Qg6mS8V4MV1vGZLD2ULexm8zUw6sxpe87p+JZId2
2TU6XP7w7K//aBlf+Ul/NoN59MHzjmusmVpQyA2zORYibev5eRVvp8IFwXHIzuy2sMaQ7B/WvEdT
whieGx7vmrnYPro3J0PSY9O0PZcJBj54xBEjr90xKJ6oDupe36g2mYnv6p/9RZHtBkUqFcxI7dMA
DbHIMNPdcQqN5Sa93EzeDzHbQSm+e8tAB2wF1kX2kufckqtLHBSIOXDL6pd3d5fnXDufiFU7sMDq
KWTdcyHIWMUAFWO+iF3JRTqvpP/TcGgO8uELHgS4Dr2gyupn3ilw9CBs8Y0saSCHq0SasCszTA5h
jTJyCjptzbnWLrMtGUxLlgXiXZ//H5MxHIHQQQp6bsR/p/e9ymfpaB36kMZx2etxxdXTwyBpYLjX
0SXcx7e1ItVXSJAz2BwD1VgaReZkeOQUXcTfaVF7ItUQ4ORIdKCjJWGxJG5SFh6iqXQktWYIJLOS
2worOsiJWw9lUtEox+kLLbnRSI4RhAETC7RsHMa/3Iujc1uFWV0NLiDalhxAVx9D6dlj2NkXoexF
K8xHD7khchLUCKO+MhNcTShBnRfP4ondAsGvpIc/WnWMli6dWR6NJ4QA4NFwfvIUliJRDvOEHYbA
LUSLpTXTHS2a5lAis0zk6k1bN0tWRGTkYb2I9igu1fY3iM8oWnXIsdg5umZ8wDCJyndGwcXVOIJs
WLLsTAIOKb9ZL+GEBBOfC8iwHIW7G0/ev6HZBMrFN850cx7ZFfLGza3PaCj/TJUF+GsFzy2mbtSw
QM6l0HmT/c4Ve8N9dXFPLqzA77q7nrgw1uqY2BYH0bkdj5N2ttP+rMOPhCI3v/x3ujingCVyioww
XpPbk/HF25grMqoyPHoUp4NsqR6s0wNEczAAEHpwLt4Ewg/l+J7frhX9ynJ8oz5irwdqMm+1mmG+
TsEHfiryDRaC2dG1IwboqRSr/YLtGsF8yqrLuAlkQmHB23ap+hE0HEKwPb6H7l57e8J/D74zCZTT
7xaLj4yIHGb9eLXRtnWu1VVAOIG2cia8Pgz41vtC5fCxs/bjuo6s+ibjtuwIUDZGQBAVzyUlZcM3
qtoXsTF3Tr2YaWLljt0oZCXYrZdDHpcpnoQXfRyzmv1BThKEGFUNrbh24+Gb3k+XjjtEgg4E2PKm
mxoyvhoaavCIOIWuCARK/egWZlQvvUCwQRg91LOEv2NXJdir59DtakmxMywOqVa68JcuPyKgh0YJ
cu7j9CMYUq98hA4R5u+TmXxdKhrHMx8nYftGRQUiv4G3HjYD+2bLS3IbcQpFI8slRpUq1FMmv6wf
C2ZhzlKAVBO0iVSszpEy2Sc8kNc1Uivq9VEKrqbdenRq6f3ItqUG/sCBjHLdXG7um4cIBZa62wzC
0paqHcSWIJrOkQcccFR8tKTGF+73S5T2t1kb64djsrPxY9fYpR48i7lcpnD8ZkZzXBr8gdQT5P7Q
6qCFP9ms3CEmHGPpH14NimxCH4KgXXVMaAh3N0pSl4CNVqERhjEPnMZJGZf2XSf1xuP3GCa47hvD
T5h/RTR/CxkiN3gf29xVopom4QW3r5o08WlbOdEHiG9fNMsh+YIgYR/03vHe+Hi6fWD8FIpsW4Iv
lpmgFWjdUXoh0Fb6MTnSalw5YqhEnAYoziBZjQCHWIrhfLapzkvXebsabJKqouCH0iRsrwxJ6XNy
3RjMPqYChXTyvsh6skVekIEpQH9IFjcWVr7LXdHr0tldFC+bNFyLx0VOsDri/ZY3XDT3mwoogXZY
LpMrViykOKf4C2W3HADdAe864oLKdk8Xyphf7v/0/oSapj42Ns6zThLCeu/y/A9y+NoPT2A18yQP
ZWASQscyoPIakRHW3c8A+t7hL07JN9Kvg8pAqSHPqS2SSB1AviZ0OAlQhmeal6eKYBeyIQ3DVNvV
9TdPyH0HL957w+FBEKvSsvRFTEuIVBfEn4lpbQ4mUnPJ9fjhsSFPUj9EiTRJf+JemR9FcG0hgKsT
YbXVrpN+qDYcRukCzreRsj1BIHIxH44txZrTtCfFI/y8f+Nhi9RwpDlHEAa5gXKMrA2nb4OiHUad
q72bb4oKxDkyPQEJVF4vBPbQP4hoR7LSTrJGKbyNMQzjK/zjzuytFtD5z6jBbhC+oyksA/q9MeVh
6KMd3Y/lamXd8pv0ldCTqvgVn2OMlGGemrHl95hl+pqrYONHLbmKJcZh2DWsNIlCeqZ92aXhtt34
24K3UU5CufX4Xov2rW9dPE0U1oy5u8Gymm6mKDO3vWuu1D+dhuAcifSeHc4w7TvJVpMShuZk5bAt
PqINMAd5XKYjvvjeBSev0/6JmVIkHUc4TZUGCt4MMOB5+5TjzVfubCwsPkca7UYYaJ5a+G5N/0ee
DqqsL3RGjhvodjWvU8M4xEvxqaBqiyEJnAO6Qa30DmLBWokeOvmDiRJVBnnnq86ukw0gjibRuaXg
P0RL66tNxur9sLqu6UlYOPAkjiQE1gweBh/v53G8CfleaWJVRzoAQKsEl0mDOSjkJdBGRAN/XaqJ
tv1xu/k/xdm4ppFyotpqTvB+JWQ6rhkYj1n/3qLKT4QTL99K1YfJPCxMypmx0kusKv82czlPKnQZ
6B1BQIEjD15KHXmts9Cd1RAwU7Zfonwwnwu7VEzLkeSzvSxxsPGg6SKNWaNP8mrXvsFz5YwLCTRL
Y1+Lr5Jaqx9CEDemllYizpa4fWZgKNGC5bx30fjY5uSyQvXDwUd9lKOSx9XF3Saqge9VgpuIyOZs
lEG9T5iDQVAP2wyUhq7Du/HFRjazY4URXXKd2FwyA7t0DfsTYbv8ViwXqZK8NWutF1BTF1yPPase
LwR7pEc3Qk4WawGxM3M1GgV2nwEev5DpeEC315QaEbvU53Lj6LmZDcUhFzopqJRaAJJLnaPbDX9l
uKYwkM6iAO0a6cnhJB18ZWp6wjKC+ihGA1RO7GQWtOojG/64zmUcB+pgtCgf+vWbgElcfYe9BAVN
f+im7poqTiVCyS8Gkff/n9MkCO0g1mSBgYIcS4JAaLmxRxerybxHOKE5ZFm60wXO5Nre2xlO5Z8+
FKwFin5i88GOB+HBNTIoczOpe+O2RSem2kLbD7BBoMP9dau5bDK2wvCCwPLeL6OcrbRmUSyEm1pi
LDcXnlwQ8rUs2UGNQViIWUSOOVh12dHelsV6ydNNPAQqNLLXzftGRYILF7I0Yq/zSjaLDoRvZyS2
rnvqcrHqutS5PaTSi144ynq/NKc0E/Rrk0t+VH9F1JGKhQjyXM/kgild5H8joBwXARtlpPKjdCQT
wU45yxda6EOM/E2voJepxSF5b6K3twqbsnXBU7AnR5haXG2CBiQDVZZ5ZwlWINC0YrXA6Wm8I4CJ
IAx+sj8Oh2QXKCmvcZ0gLIpuBIqbvFvCgQO1bdLLQmKdazPDlVQcY3okXp0kk173NifGsYaMu9dS
zUNzlTjnze9594CGZ+V4LXZV9jpYwz02IWZUbcILQJ/qS+aD/SJOR9o/YmIOaUWGINaY0i7TjoF6
g746JKPAq7k7WEuHa02paj753hRKuYw2sslWMvhx0L9xSmZSFLV9v3bbzLfxpCgFp122bclSsmoC
0JTmcSigI+wTXCmEUIczhloCHLLbYsteXpySjeB9RtZqEqGkibTnlvJcrO9qRddisnhudCftxTgH
ofMXWOR/yoRod48pJfZfRsZDIqv7yQhf4qAQfU3POj3+J6RIouGmcLf5F4zRb2e0HWbxKw8cMTAO
WxlXJ/Ykzzhjcu0MdCi1SRMJOhBvZcTjSTy53NLLpFgLedZs0/Ang4wy7dM9uxIyy382resgoXWn
Uqf2VzO5D2WZDNgAYpxilhOmKotUaunx0DPwU8u3Ce+UnxaRzkjS/dtqPoIJrdUOgsm9DuviI5vP
TPihlrenqLF0uaemjxQtevH5oQp9sIWFkVyObE6kgk2G6GsVfffrNot0GyWEd6mKd8+EECQ9snYp
B2j7kCHQXN4tGS0Q2F7RrxdY1mD6CpCByYNBxzKznghl5h71Mlpqw3ktpi4tAFjdUMR0VG+Ck3HS
yvRMYcECOatzrRZGuFC4EDFgzRJ9vIOfb7+wWyJTmFt/7p4/d5I8M95SwKmglY3VqxmSxJqmPZll
WsxIe1JKLCx1nHGghZXLsEY4vl1IXz+wEByjbS5KYcHUVJw8wCaqVzhAgcvAqd9M2PL+/sM80K66
zgT2moEU9TS1Ml4t5/ZZ5tHVqg04KUJ3vU/e6JKBVV1soX2J3pqL4uWW8rfxalEKIn3HkyTA1Ez+
UbnsPNTGDqS5B5C6UnPLRkenTG09Xs6sc1mOkswFutswpY6k3GXG8aGwCF9lAXXHbX5/VAUilUDE
PWZBSXMzdVsKFcd6ONFl5sJkrPeinJNSJgopnN3eb1zZHpqkXaCxNvlgQulomql08iieg7+HHlcL
RJWTYiUrX6fpUYjL+6uv/e9T6+tiN8Wyn6OVkGa4rOZbf+SjfencqhqGgKarCQbt+EFf4BODMZS3
FJPZ/SV0ep/tnHfIxTwhG5VjCnNN3TNATnpXcsf4JCQNNJR/Vxvovno/xxaQhi2M8Goza347zbsB
hHo4R/VUdmXJ9Lo4wR46pwaTO4Ay802l9elnXjdHIL4B0aAEbh8NrPI2KfE2L3e+C4x0Yu1XFNpJ
5CEQJ+AfD2fk0mieBZncSiQH9y7kovRTBGL0KAlJXshgeJWV2AEdG/SJBaIajBTf/Xo67aIRngia
o0UF19ZZ3QuRddag9NhkPNDef+kE8U/N14f1wTtL9bTiicNh5HlBm8RTRF1zKOZNKyoVxcG03dBJ
iVLaf+FdpHygKJG82obKtmjoHWRCoYJhLeA+lKqNUwX/8cZGKKaszGbzMmBTlYITmXcVE4EJK5Bc
TGRscZWGzyRHEqPcOsc8X0eLBz3M+fbiWsKJhEZijtke2IsjMqUtwUpyK8Cm7GlnKmTXnIM7WX6T
i8I5xnB6Gccs55baZ6lw3Q0/3p5uonF0mrmOw11dKLOPwZIkc+uP+39a9lbkDEPL/hJ3OUlv8Ufa
iCpWGcB5XW/Y0byjM8b819x8n8rBkpcmYIxQTUi9PncVFmW8r8UbAnKTB1BR/xFXYCrNDh3QEer5
fLfw5Gq+9Wyo2DGxBraI5v0g1DYkoTUDENRRIzjrUyMtn4rWkeS9RvF36NzuhV4crj0kwkHHITSP
UoGpVnJgIjSqlt8q5399a/JIPLmopXJoJ5SHYN+SrULDvOqvspJcjN0uODXhW+nfqS9a5kMEFG6K
YExDrcYaxT2IVf6a0TgAEtGItiwxfsIXBvV26jhUxT4eThxTTBccsv0I8NiqKKOX4t4WptV9OEpM
9vS/yE9Lju3p9iQR+lu9t43uRjd4/dxarTX83L8dQVd6OpIRgVlHC9OlkbFAC4VaAURwt6sa4+Ls
KGSZTzXyp2MZlehSYAlhKNgJAKo/zZyaHCuLLdlAa3IUCYz88c7Ck+dWIystD5TYFNRZLmSuCCr8
2Go+uPDk9I5w1bqSbq4ppdiTy968z6wLJWvxmbwBVCp5R/9NcuYk7PhXS6eWiHza0Ctqx/vq1IDk
qvR/3CCowbnZ++IJYaJB5Bp8l5hF2pxtV+SXX/7xx9/T9GgWyJBvKBk3VK89FYvGSyImV48ZBEWM
Js2istaP3/0npYtilWn6n07ZAkq4rs0A6DxlmIPXVEU7WKZAdDFu60lYjTHwmEHFkYKQUDQFxbTd
CkTAn5l5F5QUftx4QvjISmtQsgCpcMH2ntxkLikK+RYqrCKaizBfPV9Q7ATH53LlhHqPuDjHDMoC
ZDGdQ2elsB9VDk8UnSZEHon1EuwaxIrAxnE1iWGaLGwA5gCFJXrq8fqWJxCRcU/QVMt8K+V3mArB
1V+87HSvmxPzfsmxLGeE2GuEElfUKTxXXdN3U/p7Rsl4hvn34VW4DZWY+kkhGq54SZk9hlufrUe0
O+tJhgXFvH+v1gkYOzNgbNbSmX5czSmt+dCebPimhBRoFbFv3WUp9VwJfl6Ik2o59G5laNe13hBJ
9bxsFlaVmB7+WiS0pO8bwxJmXIK4Xkv3atdmjXC7CHQtwufg+WIKI63WnjAuCyxdp5IrjwDQfWbV
JFRyHOEvD2pxk9M0w4Gdw66W/7X/uRXh7WfYWKtTVpV/cIgen4amOCCniG6GVqXTKC0raJ4gpTSK
HZzrRnoXVhr74MHi52LEOEBP+TzuV0B10o0jKSzESTRWgxA/puz9BUx5jlqN4f5aGHqN5erUynF4
9dBDsWUBiecOAIDNiQGcKxAPHc4CH7BEmvR0bW5XUxFo+Aqpmllrjd5hP/BoAehcj0P412NKXRve
ay2SBhiKr65z5+dmOnHxiYvfyGnZlUHkPamAsLhhebCZf/mzAO57hV2iGuRAqKEbsrEZVdUHBtNO
w/Fbt6QHigN4nyUruNobVHcj6bTGumbc4BIQX9D3/lWHDtP0MLDXpBqTH1kISQuJo+OXeiQsyNvl
XYEC+wWHxAVClKqL6kkbfTMI3Q/YsNPOFrkOoQ1kHn/WjQfSqgxPYdVNISN718JcLRzA0CZ/Y9fD
NPjCT4VkR32X71liMQ5VBuVSdRaTudjw23Gz5pvC08RjL7tJLaeGO2Ie+keQ+pIlrw0q5GMhaDjz
YzT2o0XgtcuqFhux8KViN/9hXXUJ0rwD6zWclA/rJRuNzqkMDPFJlbWADjfAqG0ZKoWSLB+Tw68q
xTO29F96pru0ooOFUDT5Jleoq9Zu/c/qL6ohCN5C0TZVLsTG2npT73ZDoQApi8ZxjoCnMhnxposi
1VsmXgvGpnMdNb8NJkXEVl7L8cqJkpGlvQWveHY4PEApsbYpuPkxdMt2J7rUdyX4CRIeqvP1JL7S
JJsFCOTYwN+H+7fArNvftjdJzBVYFArJ8imlHuBABD6CvAgYz0f9fvgKkf3HqdSAocmN5F+jVJ21
0CiJCwdiZU1jMqiSaawkpOHwpoMSjsSKkTlLQWmDX/7uhrrGjSO2Wm64HjZPj7IM0z98fII4HtSV
0Hsfq5UhlArnTPQnBMmGLSESss1VK/n8pcxKodHZnr+XfNTGsQVVLYzpsO6pnCfw5tv9V1+sHHl8
H81dDLiVHarUR2KcBdVJz1mZLBY7Kb+Hbr82MKXHBy7F8/IWTV3Bf4i8EvSQgUOq4XYIJTe/J7Of
TgCJu65MUjvV6Frh4nj2LsApbUP5pnUKstl8CkC3RgzGR82/1B65UrpjZVOlD3HLOOG5wew6ZlrD
tOWGvvtuW12KrUpuK5Z8cDk4lAqTynW8dDd2rLCS3Vp1mgokiaTo/nN3uhR4XcLvnAzTNp/c7pUj
3Uj/wqECRltyBnNitaK+GK1A7c4RdeDjwgd6zS1yYeyqlzGutwf+6fUC9zxb5c0K3PZSXdUlxa5h
TUY2Z4gNWVTzZNSGlpfAKMEqXTcsEsiMImMKYgvHhb8roRlCLlFjngxdSACPXNvym9ZHybe0H2II
PkTaT/SkKhPfEqTaP1/MmCfkI6Sn7EgKmArDbtw2Aj1wGa5ukVQp8v6b/c731u1XPMGP82QIRHmF
qr7CdGHmvGMotEBAnij4sH80Aoynec9eXa4HCo+AHT1HRtfXOzAY97NZH65OK2lln2Xf080fBu7B
NzicyZ5lr4YbjFP4vxTGDGi8WlhXq6ahuEq+2JFMfPKJKQnUscy1FCZolv11NkE9cVEpPTFj+N8f
VD4/ZfV6L6ilfFUH3YgbwnkG8cAjM0iNMr25sF1wGopBZDk7JhnMRbE9UwbvtWFa82J/4lOkdlox
eR8/x6B8ki6+lxtzs3QuZf+gfBj1Tqu9s2USuwL2bxNETbRDYTcppCwmwVzBikD2RfMhdjgcIVxV
tRRpmAbSzZLyy182DJfh7kOTyfJrKxenhCaSw1HD9g5Y1GG9wuf6/6S1F2aoBqwhRg7J5Zmbw/qZ
1n3IqjuzC37jRckqXhTnpRGv02xFKT7scpJDqseKkRZQ0yE9H8IJkv6sy8I49t5jUmaviKicsHKU
Ofzpq3S41Jctka8BP7io7mnsa7Bw7nKxJbqoRiViM6VHMzPBUu4xpnxsO4i25nWc7Ql65Vz3ovCE
zepf+U1pJ1JQIhC1nMvsL+DLZpLs/Dau/vKQAQTndrl+3aePF78mVvYdP+k7CCVwIkVnbISQN5h8
Kp8OP48IBNXQ95L5qKi9fIWeyhoE3pfemvGOSaEq3xhrrqoavIZFOXE/xHQTm6VTBvv0nXd9dFH+
Z+PlxTI4cNybI6dPjiJI652dqGq2qo5s398cTeN3eaVFb3y1Oes7HGVyAcklX5LWlej6GFSrM7ds
DCoZerra8Mh1KQgQvoBiMiTEpC5FbaleTJOGT7dVdhA+a99PDeHYMmT6xWUsRNDL2stjrWdKhBlp
zrmDXr+ZLyqsdD4ClP6aNBydxI87YNQb27wtJ7FcVXJsqetTq0571G8PGtYg9P+atKA4Ie493cKz
f30gOG4mTA87IoG1hZorLrty+RtdHKvwPPkb+/LveDGgdmFYFhmqCkoRrufc4ovZlI0CXXU4mX+o
BktebsdCK3ORQz6sRThv5QN7uXx4dbZFiTX4Kuq1BzSSCmHeTVayx2kX0vWG4sD5fE5Ajx+oN7UG
Zx4Do4BkdMESMa682WQR2sP1wc6FB31sDvIekhWvKOay2f6ngGbpaadmrQSyRE33i4PPr0CcbVzY
cf8mhK3uDvV6eHBOD/i5Lt+ud0bgQ3A+WH2ELCZW2syQeUnr2NGpRWjU4WNaQ4697uU0LQemsh/v
QsEQxfXuh0IdnO5D2/8stfYSdy7l2mZMxlYyIPJrmb25tHDqHV4BRy3f1HDx8tozysMAeFbqEV8l
NnjAOSUoHXQK07N0iD9pe16YUvneMm1c31BySzY3fpHMhzXuEINZ9D/B0aVoCt4Ore9GRxsuKR7z
6qnkwWBbUmdVf3thMOw61Fo3fCKCD1Ipp27j9GlQqtRC3XRirHvDPfic3718PJwmw6G9851rExiM
kQI8v4s9ALBcPLiYYbj0HT+s3JbsE5ltn1GkMV2IhTe3/w2vn7mYr49OtUEIuvB4LF2jYEiyCQOt
AjuLROUC1yMMdgce9+34Ge6orS1L78/0xoxHYA4Ay0ZK7TWJ7V7rXLVy0bfLlGjj5kLXLbk1G1vU
aewj4s62ym5YmW3uARsbJnLeATrD5Ss0swM30Q5+RBYROgSMn17f+6Cj+G6hNpQ6a3Nf/Oovc5Iw
8lrKAejSZAfTQm5jld6QE/N3ki//1IHZsXMTe0N3szv4MF/ykuupr38UEdCtK5gg6i31398J32wZ
nYxr3pE7Mv8zNVSJ2HWrB3fCR5+kPL4miUfrlG9Kxrv6+XGM7tQ8/4G89ELE/PKQ7osK06yqzlaW
z6bhxKy16Jc0ZkIr5uypE8LEC1USxIy9VyBgHBEy50GWA3dsw2PZ59nFRpkw10ed7i4V4L+aq++G
VNteoPRZHL4PYTq0LUKFvw6ysDR85z1dH0cTv1WhFR6ISBGIZryvAbLCzqwYRav8T4EOeIrpPREV
hUAsobPaRCQ7LusCzJc0iNtwbZAyHFbgQSgie/l9J8rVQKPRgnrZuH4glpl1HLVHCT+l/vI5uvOe
WEtkjWE13Tqej37wzxAoVaCt2oHArtDWyd745rs/BtGdZcugq8VNrDZko16KpY8BaQy6TgE7Wa8+
oSiFEG3Dfnz/vq0TvmfbALzTxvTVCMGLD6QiqhUhZDGrFuwYGgMnU0yL2ittydtXHnp2NLnPZLl4
O7Mic65LwfAUL8TamRz59goiYk/f4NXBYXoAEvEMuimJ/m+h7MOo5VjSizOxjk4tiyqE8qSI8IzO
H32GSRY7Z/PuhRUCoTDqdCyDZIHcHUKIxcVq0YNzP/bzkDasQruAiGzyS2ctX9Wa/MJiFZ4Mf4T8
Ca9YGViyGUdWO1rQZB3qjqJXPn8QoVFwJv+DDi/aHILJa0r8ZeYoZsI9/dsLEeyvOc81xDP2uoKL
3JbHG/QjibSyjRvGyTw86TOD5axH3DXGlYlshmz8N5CSjZ/wXA9DUaY2j65+E/PQlffhgcUc6W2c
ngU2SNqts6UqVGRh1KCsxwbZ+i9iF0OepHTX/hWbRL+VeldBZ74vmLYXaejwcF4VaTpG0DivvqCi
yMU81pjh4Td81k9mlqpi+jxPIzULguC2ms0DUm0EuaeKk6WyU1fZxXrQdeeOD6Pl+FtV9mdwN7xT
ymeucrrHpXgIaZlkKILrbg+TWGA+GOxJGymabIoDDAll/DGzLOwEFtiblGa2QS84GunvkWsuvKZk
AshiTt0xZIocwrR5m0Y8uu7ro5PM1TCVS5tWIIP4+tYJYpmZ7sCIEcggcigdGzHCQ5SaKREuJmfA
YbS0QuXLtBL5NhO2/KIFvGjeytEJDaTNf8N3nlMbu4Kd3ghCutBY+5TMJs6Y3rbs2o6kKFIM2d1J
uB3BPJgdMQqmebLAd1yleJnfQURMoj0mFPzqZubTbVkoFDFy2voUUT1EAHXV9O/X7llS2exavpXG
KD+G9+nzQkr3cz2FB+aaUoqJa1OFHry79y2pbMURzgdLCVQpEG+l0NyCv70M+vFQpe0xfGNtrEs7
tczh/AiHRp2iZ79UReivEw4pa08svbknTG7ALj/iYlMr8w5jQQTxnrPS5ijXqsMYwwRELxZlAtdx
t0oHOQzPQkzuUt60pcaJZVF0ctvqPPqGva/n4VCX0ui3pYxDmxqghEP0ZrW5Uaf/hIkl02OOgxh3
0p5Pv7wiI2uIOrVwdtagHim3QX0ri84c3pGBdfww92Tw4BVprISBjZxGghBPodPxdwVQCdjejXJ/
Z31MrEzsb1LaQuMTpJHjGltO647IDcOErWhwL3NBftaFJU7XhimJ6c+GAXkn7JTH1eF/AokTvnpC
f52S1kkTjNk1XJ7bUBvu3rvZBsZLer+4Ujxn917MDsZsIeKjB8JrPDvW96AvGM7+hJUoCaIEoaVo
/YMtPggzK5oh4v8KTYuqPJ5amaolLY93fe2JmYqY/5uZXYvQ58JcpbTJGDBlEyqMOT42PM2zyv+8
bil7bgwS5smwLh7dSewQokqH/ERBCXfqllgXQPnf1+XW+9U7wjy7Bfs4y5pYdBFDx4iWb+M1YNLs
WCE5IauiUBxuSFRfA+FQxIoybx9ctJGvYW0R8C3tdmYusobC3dtrUDoqyA/ELRaEgxfgWdb9rcsY
A3SCMWY9T+GQGTIAeSHMpbqkj3goQH6eSB86V4QbFrlc+H9fcw1CK4vDRDQmR5RLJBlcpaMP1euq
/+hubrR0WefMJLgQd0AWGxcl7vl4GMeMMp24HHBFaR8Ah5MF5fTAGk/XMsVc15kAAHeYhLtNp/Ci
kKJf3GrAMe4DcPt64T0ILFdS8+SJslhr69A0pFKBSsCqIL4SZ6W/OwnX/g0ci+2JN89XA9riBgNN
zpnq2rCptIM2FWt3akOF9zwWCTcWwwITgF4jEp0QYPsPh06GXaygIi8suKZUImsxRHYg2ovw5b7S
zDOFSZfXjtnnyCsv6dltyf2QPaDcR/K2OkOD0L5VV09hxfPHy0Un8ZvQn7MempEmr7L12F05N5wr
FpTE+MP+y0OCJ6EL7JAajCCGKmEwT2knQrwxEL/ItHjX377XTcroG/k4iM7JYe/gkeatZcYJX8dM
PH80h0gBGrQ0JRbEJiZioxOn3ojgPo5ztnjZ8dPbWa6hizoYTD5lnnQ3HMrexuupGgL2O8/BmcIR
eupzHm0NhCN82NIveLmwjqflCt2PgP8Wj18DSfebVYA/MjKJEef177RJME/KC+MF7NxZ9zEHbG+3
X8SEppsz7YUI/F7h/HxMdxKh4lf/p5NJ+szNpk8ewwUsywxhY2KLwcJeVF0QDnFF5K4XQtMzOiw4
Dkr2lIOgrbm0jlveUNf79aFjk81WQggluHjvut4oP3s4GgPyA6H46/uHBUntCO0z7jjAZgOv6qaP
3MgCatUlfIGFbwz2JPLt8emA2GsBwllP+EXmlp3i8nvbvTIcGoIbKt0nlaiLzshGUdOY/m+rV6Ho
mIWbNZYg2REeJiiVIcAXxk2ff9pHxHrN/rGGj5/rEpxk6xwL6gCPId57bbmBrMLVVIZXaQpjMDGK
e44jZXeV7mAP70jcTDi5mMPotr/JTDrzBiL4mmwpYPQKETfNIlBYnDP4perEuuGNKl+qXl2QaLie
cJNcUWWTR3rxv+SJIPWdU/nbu3pKl2adBe0h88cs5ZKNyDGKpfEjpfEShGeOj7wAMjn8TjsP3p/4
xctYrcYaakQwoIOp2QBxaF9kRZQMSnWyUOqEe+CwzLFo71n2R/8DfdNRKSHKQPiXylF5J2r6QKFu
RfPo1Ut6YQHU/m9Bubrh3SqrPZQ4MKAQIRemECEHu0GzLNaCWjaC9suSvWk1I5pzK7jMIpq7GAKy
5lFzQzRKsgDjrA0fOiNJoM19DTZ+QJ8HkLe0T1zS68PMNKcOPGlNpkp+S1WZuOlHAvJodHMoH1G2
7YjaSfR4VVozk/8sF4U96gkKrkbJZjWoczRHgX+MSeqSBGbd554ET1AmKy3dr+EUdUcud9JqoXP5
WUIV0MQudDuztluLD4nNe3Hk9Mii+smPxJ1xzSqtahf8AnfrDpoTlUQrT5Q6uX7bFF331ffiHHKL
7TQhucahQY66m8MHJ0got5Yj9pSBKCUyB17sfrA2xCs10pRaTU45Wkwm832KCCHb55CtsMTQmRAu
mBs55GIPzRAj1W+g6hiIyLzU9NuVEjPsrjkN/CpL4vHutEFi+qTiS8WjdM84aGQS5Cgabha3sTdo
KuAwnzbBzwbXE9xDa5y7yhr4SxHta7SpnlmujjzVRf08tH2D0dulRL0um7tA20F59t2BcAPwEQKz
eM5g9x1+4hP8t2OT+L627q0V9ff3gWpPG22bzx1MJ+4EfQ03g7Ib6OUe290fOpedq1LX0Q8K33nt
Sl+7AhZSlHafcYbY2cFvKucELPBjNQPMDGK1Nz/4NGkLP8/d7j7Y6xlsmnXuqEf9JFc5Y73tWq3z
xJ4Yt337p89VvkR5uhqszmi0vzNKmlj28MlRJvOIN1wQo5QY65xpQKjFRLb81AxpLilkQLUB865X
UfXn8CozQmiw04Du1sEw58gVNXay8hStNi9PalS6twxo1WGUXES6voW+Es94BM+y2jrQInBS/kdR
B2LqFdQnJy7EWBja9CyIku3DSx3y7RZc0Rg9wEx7T5ywKdAiVHTF3aUfY0vKNUjM7W0ZwvSClWLd
W3s4QesuPn75fr6OwZ4R4OW94TuQ1NyEpz7XJnb5cwruvWbCEXOw1joRW61LAtY8oJCWAgkTLVzz
iSSiBQoESRD9fMmTpH+sqN2Ne0tZ0JWOmGq3P6th2Ce3sl0Ap0wpTI/zsucolNYFqWuDP19e0Udw
AN5o0R8ZGzpY36zKhZ9q08Hllae2MzzZ5yDzgtXBCeWlOKV/G3BjT2yYshdJLP4pYCYP6zHZh0Mk
cxhLX6FOUtSDYSmRIv95ef6y2J6I//Dgt/MIu2+SxKZerrbnbPOLzZrNLzQtt+EyCB8d2ElmwT8t
eFaHn6M74aZxe8om9PaS0wGMThfHHvWq9TDPQUKQUGtIp0XvJh52cXimT3qoGUU9LHCbS5R1qJl7
pqZxzMhlBDKIvfPtjfP3lZRNvLLn3mdlu5b+CjosQ78/cPM6O2UkUzRnEd7iVMDhQCAKJaFSXt/G
vTuzgVf1mmblkSzFvvaBsbvHAkQIkFhA4Y4PL+FZR4JpUBSwE32kknNk+nRCWUgga6m5/P+3Aac+
hq3m+jTm3AEyhyA5ZSOYSC9WSNGtpDeYHsaYfq3XPwKV3ry5SNh+O1bOBVEOkge0ucbF3i0ePTKZ
rrtOqmS2i4dAtOlf8DxXHwA0BTQB/AnSSDCs0FX2eT80m3j1GC7mJmeVm8wZaR3wNZRgprVOVt2V
a8UgvyGuBrpbI9IpevAyhbET/5TRmBJn+SuF5vdIXhhvjCW5+wXf8sARnaMns9qe6z83Z9YsZ8yX
qO0vZ9XdPbnF1392s0Nwl1yCTSWSqH2wUx2YgsY5EpcP3ka66JNeIQBriusnN4BaqRLLgTxmzLXh
yVZDwP73HWoXLPchXkfC26qKKOw057FtNSQTcF2m8dk8PqNEkaXxKpkHeX1INmU1nifbxYrQuXtK
VWDf1IWHZnq/pE+WOmj8BpW0wfL6T8v7sMBtJsMLfPRcvR+2OpW2h8W9l2Jokd/NlGr7Rygyj7TU
cgWq+aMUIJ3TmsWsjWtcJHE8CzLw1+dV8Qxyl5Nltmu+gt/R/2VLHPDbBVlmaP5a6iKE2Kgdrizw
KVqrmAWso6WXYVLYHfw22WkPmhxQItYoYPALCAkJ9U7drVm0opv60QNO1qizJWKSLQdUURViPX1w
me4HdfKkJQmq4kFIpwBsPtN0Mn9CfM7ykLTqmWIUN66mC4mKFDng1VWDYpD703OvzViN1T24cDD1
xNf/f1ak43kAgTwr2zW826ftJgEyeqonl2PJ+TtZ7uvVDoSBivh9B3eclKu4KajC8ao7rg56CBrx
wEsDQNUwJPXUeBb8HQK2Bo/4Nm2Apgs291CejBrfzwDWfYmZhmIrzPGjfTqEP/zEfYd9joZ5C1Zn
BxNIsDbXtRADf7DBXid6BaVAJ5+3KLiYH6/TctKu14oZ8Vq0vwacVIhh7hO9yHmvNpuzh8JuTXST
40zMxklt0LufgJPDpMleVVBiD65FzE6psw4jbq8LY3Y7ZlOKjeXwzi3swo7Q/i5d9Yup2Vpyahkj
WDbT6kPb8DQ3fmGzMlOM+Hbm08eFBRsRZFYh5hQlskRE/OImsvYPVXXwUw+3+Jd/LCIyDZZKIdQH
2rXL0I+RcxeLbxjE8hQWsYwlT+IZEqQRbKe2uKL41x+z7AaeRFQxPsTzi2Nus8svhr9KI8FTtf8q
cihuBet9shVPMWntyAkOdM0dRZavkIQZDN0EGaIGJ9leEMc7ZVLv/gNK7EjujKnaBMzlGhm/pmWj
KgKQm3KeAV8Vxb4h5GOHbVG1FAkq7OKVLj7WZ6GOP7NW4WYqly4erlFcYc0DE2qF1EQigTOxK1YT
kcEQI/PA7d8s3GBGHW1J6SNkP46dpb6c2NNQn42Vhg/Kwl4f9UZ0/Qf8gmwUQyycxLqT3pW+tyzl
aW6jNwfPleQoGU5Jp/sBA7Q4635JowSl3R0ES3w0NKmti7wxh4AncYwlB8aTOSEQNjjfdG2Vntue
pgo26StqVE/cY1/upnGNpqN8A1l6QrDRDoElMs3V16ThFhAoSL62K6/PCcztTfnueozC+R2Dsh4u
6Z+iIDeGVXKQnIkp4qgW0wPECouHQs7oovZclZZm+J5/BlJolMofd0A12cbJ474dh2qjQs43cTCm
8skurf/L3DMjs62rFTPAlB1aakAnnR/aTRRwunRQxNk0vunOqB5/PKUS3OmZKLsf1b5d2scBbGJc
d4Thfqekrr00FylqeBnfav3ETqagQNV65QUOsIrQfzV+OuAHVbZ+A59FC0wkrvUsR/eJn+798a1x
TPqPd1oi5vfEynYdnV/p5FcDtP717iCV7lS8dJ3ad3Vw681x7y+qVmcvEpKNa9Xp3/N7JwaeX/Ep
JRRtoDCtXSouwCxJ7ba4AZ4I9Wqvw33ivdbNTo/z36sLwvW+Uf2zPTKUK6SPCst5QsNrW8xwmgs3
mzTvw6qhTSrwdUdLEIXQ1MhOE7oZeTgZdpqBoQ3stmFEpUvUiOeMAbLzUvkdPMgjH0UnoR4zaWwO
6f5T6T1W8Plxwah7WLPigo/QvyrKiN9qWsV6P5gi6FTyf2k9xF27/ab0ra7/m48tBb2C62CyxRkf
NQKRNggZjXE913JYjZC4heN3jLdsz4A454VcPhuTKV9YLuGSc9h+QySV3I8UcLkHDsKYy9pZ33TY
ktOPXnQRJpAzzD5PetFzRP8aPR9W5rombsziV2JqlDtskkS0KJxopJN4Gt/i7KNkFyS3eGt70qGP
NzPjtHAw3WgiFeCg3nT/btSZKiSEwMP2KoNsS7TtHRv+OyoeZWPGe8MnsJeh/BEJz2XwsjqWeteq
e/hzWj5EiBKo/onm9ESfuDB/HhA9P6rNwaAyQEnFl8hNp1V7Opl7yXGxOHQAsd3MpprIo1mU7lbX
+nCSEdRcrRyPZG97xvzXnX+XLLQyCgKmFFCga8oSMu3ix+07GzEO7CXUWOfj2vRB9TutR0GA6AxS
B2TKDtKxcIDa8cnyY4bSS95lIUen3iJry1414tNHDtRxg5WgRqEuNBCgdHr+8YSG3bqzt6ylX6wZ
qYkkZeMkBPAC89aBrUYa9CW/UDTllloeF13qo8wenQu2r4uGm3NrACnLz50MMCPUbNyfNx9jTCct
i1qUXqKtig8X1uw86FG0fdDA8KsMFLqDQeVu1dThWjRWh6a9YXjlz3ShRiWEJniSx4JTDq3NXPG9
Ov1+GL4r3rTD5oBBjxcYr1ZbYSBihzxhfJX7Llaz5fKxtCTyvlF+CrBtbYHfgS5OyRGSQw1zdFtP
MgQ6Ty3mQ/mTAhFlw60GVxLZzwZ7TUw3jU5LK2i6GIQpmkcezKx5Zj3/Lc8vXR5h/WLigZ2KvCgT
4ErM7PQwYG0Ri9mnQasImgDmSXrnvQBVS2rJu7iDGueoeQAzApLsvyIhJTTl/106FqC8CAqdk6N7
VRxx+Ksy25NIt18YbDqCCq1ykpW0rTyBFNlzwhQ70fxT+DaVe8oBrBytX1Qh7SNJkeVLhjG38RPb
dIlsxDZUHor+srICN1upstcol5WKTGyL9s+N3iH7yI3wtYE4zuzHYkNFsEeRjpsoU8KBbqux7AiQ
KkC/QT9Ce+NuHbeVYRXOPuWmcZzsXoNItu0aBI8kP1pkwrqb7U67ikRdhGSZ0AVEnUt2DuK3U0rz
L+3sWymqR6ZdPUFmdv0b5KY2f7fjq7fjOUoX6nrExdMoxNTzikjH+/0BxghfPQvDdCSI7NqG6lbL
xTux1PxeNDi3KRC1VpNM1Y9c9d0JqKqSSrNkJmSr7BIV9aIyTK2m4mXISa9RKpWU33GzzxRhstHd
ib2NKvy4RyUBDzEFoqEqHFTjXFvsQDhXXTwFg4s93GeYhCxcyIL95PlotuwOD5ITqOfdgSD7BbY8
xxxMoW0QfeB1TKk3vtXPBXgN3jd+0NqWUJlxGUzV7yxhcHA4gGiN228WVZCHPL+R3InrdEmV+QpM
jAfekUZUK2XFGQvPxzMaX9plneVH9emFPCAX1LMir+eTDFT1YUOwTT2fVsPH9/gI6TOeP57QQgCS
BkggaPSUe1RU0YToqTvYAkOGzXQGnS7NOBu/dioL62OZrL/uXZSP97fYPJfVzOQxFp/KXevbhQyi
CTQhe3Aed5nxcv9m66A1Clh+yf7Z10jALB6f1ZXpl24puDqH5XIVtHI7yzrGPnppH6fvucWpXFI1
WfhuHNV8LYAxcABQAlDy4GUiQ+f0RPdy+83TnEbc46TvYZJiF+OB3lTQMBZNqh6HWCBIvGF5ix4w
CA76IVwUL0JKQallfTUCpwxaKOH5v5CWCM9T9ynP6Lbrzc2bTuckm0i2L9bmWu2KmmXfEYvW3Sx8
BvZ/z9H8sVj6pQK/0/sfk7UOciZWUFu1DTmLuQrHhTiZcX/yzhgHHtXGRo/nHtwkjKEQvBChMhOk
GixPwpxi+DOZHzlmipglLa5U5tfU7RolZ1QsD3hw7jA1b5YlV6o81inA/IArcOGxONCt/22tXBPp
SA05xVvfxBx3tBq7aMZm6OnO04QRVx+zixydaHdWxEo/zH15NfAlr7Qs605zDXdb4FCrw0nhFBwD
Ss0RNr4MLHwikhHwi3Yl5HvEVeoWNu5aKG541tLVoIAgrDfaukYfPdQ85XSLOFLQwKGdjEjUsjLE
jKX2a0r53YgymkQRkpD2m94zibdPPk+0Mpd79rA+d5kjbTUUhlbZEUCsrw6aEm78Q7QGjzTdCJa/
nv7rEWJy4oWrPHe4RPPIlu/MzS7y8ZFKuLhJ1Wh7aG7s5p4Is8aIhjd3HTyhUtkltVsrhPK5U6OE
DdUrSe+191qqf4QVWup6gfpY3GcBfbBsDseZO9/UWRBKbcscDdzAgS0KryPbBjac/HT7mzfyTL5u
8bQkvAWl2La1mc+St+awrRdWT/TC5cruoQGGIiNzCF20hAK4plhiaAzUg50T/l7GGn4wVb5z9pGc
Lq7QDyTKi/pU+pQThaLAbA/Mq1xH/zyreLjzKI8DX+eqjwdzGCb3OXYOAufbZR6+Qwu2WWsMWFxi
j2xoois1W4EIByvHG8/9pftFCOXQaADRRMyLVhM/x5fv+NQVHLLQVO6leyH43NJnA/KdgIg2B0aJ
aOJrq49WmyP6UEDxh1wts2j1/Hc+SteP8hgipd6TzzuAZrnROQBQToW7VfE+SxPaZuh/J0z8MIkX
9O6cl14dKB5TBO3Wl3GvCMut7T7dnS0pPdPQ+9msXDIoZfUA44LSrQHmrveWPoctqIXZoGOjvChZ
BHwczHKCG860m06WL17le/ao4w3Yy7EClOwP7RyJjCXKjrN+vkusOpcwsrErtnjRcGaNy3vo21eY
wbOLElpZsVEJhfah6vZLPcJ8962KK/vcHQej+XoVw6WcZGtnzwQgwAhaXI9V8cAhmk/nM0JzhTdJ
E/3DEFft8a2EAJbYhF7LiR+h2YoMBEUYB+TNw+O0VDQG1Q6GBL7i8sjvwCChtFQN0YK0dkEzWCZJ
9LVOj+RSerKeSSGFjjw1Yv7V57HaeFPDXiYWBBc4l64KtpTjq6L5qfVMPMfxo2cwPqgQAEXqW0jr
CGD21NGCLqVYfK5tCLwibVDUemIBtOJf6nThNeKAilmYxA1gC2jcogomTN5/ULYEpUdW2CQIGpzQ
PTyUDHrp8TeK2ATkhgh59uFV5tbJGHVMTbF3UfWxgYHNZSaPQdoHdNJLNZWombrj5pHIHXx8aXfw
6wMt+3/R3glrjthGE78PhmA/86+TtuvhwSuwWTF8d/bDZJHtJnyJqvAks3h+FpM0aFilFZagdrSO
teojgXqwOVZ2/OAqPf5UbWXwTnvpx/j4FQux4bFtA82nuoVpk255ZpM/sDdIEZ4Rm8LM4SWEA0fY
trxcq3j8w8rUUo06dYaigii4nsI8COnsHtuA/QMHbZBlOW4BfFl5aX2Bnh6FRKBD/BTK6ljWtE8X
ZmDbgcOKrI5h8fSDOgLV9IpX1Kpwni8Ts/0ACnwU8vuvO+EWFbH+hqH36FB9+OLdy408FGwfNVHa
H3DjJ0yPU6LEnQPtE+GaiOPn+FhtrmzrynYjZuEcOVe2O4fhQtRLR80tXsi91ps0PtyU6uLPauwI
IsdOmlRlX2eYjdq1kKSfPl+IrxzzSIvQjIh+vUdXsbyHrgZDJqmSQ6vqxKucEEUjDWIyjdu50nXL
Rq4OOMCJpiDHlcq/cnn6LhrVnMa3iuuIVerEYvnpowGC9hXuv9G5IBmI/W4VrqneYNcnJ9Ibpp+6
jdVns7nUIBhQhrpgC5CUjVL1dxeseFMBEiUFc/Zp4xZGyKGX8+hBMz5ANr5F1G7GnW6/LOHHVOdO
5ZzyTwcVl62X2cpNz63sEoMKBeI3wFtFCenoGNgAjBvUCjoOy8+1z7JGuyQU4ZYVocM8tv7kpO42
TcWC3E9yMuOn3UDGsbtRsK6/ZPFnOLGTmnOQ4+gnRwRnwoGjtUCbD7Mqm5oH3MeJFRFGedR37BXn
WW4E2scFLtJuYCFUTo0TyJ95X81tuJpWhL47UhZs31Z6Lx5RM9gzLMgyyUMnWfkDZN9TgETdE0U/
uc5KRzYj2gQmdz3APqvQ+UCRfm2jWD8FEiNGOz648BHXcZcuZh1lL8qwwTIcdm+5cTCe7XJbKTAF
bG6zYmGFZVafHx4vdfWNlCIekZzh7zBRE2Teq4txlZFnkd3RFN7DeUid5t7WF7P+N1tNw2Wq9CJx
LV6m8udo3rF8XSV+iPUEP/BcTqb8YVCL0xdI/PHrn55nfubxNuPmZonRc6pmGQzlUxOeL6V1R/uq
HN6jb1vjpr1J8IDHFtCqsNAJF8hLDCoHcEGO+YtTUKRTKJdW5mMXBbRcHGm4AJc7zQjDyW666sFw
VFkwsLNPkAWtGXfMTADi2Df80OxxRzH6RS8y/dpD08uf5JyDtDrdFpIFSArz5ZyVXTfXeO0siemE
lDbasNsWfgc/58e8Kp6wi0ggu2jJKFe7xNV/MV9OYaVZao2Bay1L8T8DAUdGwoSPDEjVijvR2u4W
+/k+U6IhFpiudGoRBMncFxhdrT4+5y2uz94dwYinj6RixL12yk4YUgmvfpEkcTRZVjN4HSb8GxeN
QHWMwpcJLTK3bmDXZ5o3/+cTKQbDCxdUlDKTsb9VXb500t5q/4U2YLM9mMmbe16yqJemrnIyrx28
4LKGxRo1xLTUegFVZRQhamhKQcCv9x6g8O5gzk10ZOmDJhkae4fsNOEUiXTbODSK0DwIwSYEbivL
Ji7QLMuzDw2g+7Ryur3DaXlZfmTIzF4WielkFvpBghzcQhaYBzis+vTrWqz8mT6jSD3Je0WX3s/+
at18idgg/Sxunew4e/bRd8gEkUdEzY4KYNkI1iOzDfZQjcgBakKlKyJaQgwbZmU/e+bMZAPsn/FU
0YQRyfCx4k6XKJ0j5isAsu8cka+m4q1E00kT0ap/sUsbEblw2Wb24diXZZm1heU5hQsJGqla5Bv0
3R3ipXV9Jo1UnYlndZD7oLo9iAygHYfnXjNl+YnuiUoAlUanoNY0BUcekvZnYvB4eX0iTFDM3hMZ
ROhdkIG/pzDxOpgkbJX9VpFhVfQPhQ7d+lI9vDt0X774vJZhcB7yL7K1D35ETvg5sh1Mjv0Hvlff
kNEI7cdterZs+/mXOq5R93QULWksXGvYeWD1jAbpo2AaF6Z5Sr+qYQ3PIpxzwMmKIvxNSQQ2OOIL
K6CvW0UACdcfUlqV5RD/tEKDMf2IBu0fzHhM0uRhCXcGJ5o/NJgoRs/mFHe+Xw2JPIZlpvkYJ25P
cjKNLSJx5Df5b2fXP+kdjUvsxHRmbJYVUaEn11xZxmOKDth5EU3ILiwz97cAW5vTEQyzuI4F7Iae
PMytlvp4yk8QaXEzxFEoBOes8/aV/8kUns3qlPQwgvytsRvylzHZiQYZ52gPC3+Wdngc2RJgEuMZ
o/AuzQfCxUPUSu6WPv8JFW+A8Jq6h6v9ujoM+YeTLjpYzyih5RHVa61fSNhNphvpSk4O0qkt/Q0k
vxoPiw0KBM9KToxv3PIc9eXNfCyrceCylykZqAEWwKpk+7DAJUYD9xztEGC5a1UbjUrQYw59kWNL
GD0fHvbixIGTG+OCtNyviG0RQ/E+k1+2GHQ/lpfLUkuzbhCZRCA8r0v/F5fhi6HwwUHRxVyhYlKD
SI2ufouhSpk1EayWlCelALlrYyf8OOnkR5WfAC+xuRV07XGES3+5yW72trL9qiBxh4+WZ1EMEsmO
CCVyCzW9AKyfSRGcYD+ONKG5sNXG69bUG3sTA3J5FrIIC+KbDJRnzb0TR3S1RLXut97EK1T+m5Z1
0mSGy1Gp2v6Yo1abV0AeCaNY5/NUTLV02evxCW510qM/cze88sK5vQozR8fJjkgtIWyD3gRAE4rU
fvleOImAwI1A3bxlZOAAUfkHc++M7BuLHiyxQUubCC87sUZsurXIPN5cSgZpw/PXd4/1QGG9tlSr
UliTgEGjAQcY/9DebNz1yt4GFjBBhV7I+cqxXPpXrYoX503I3rWGtzPLBeKhMO1w10a/jtggXbq0
sm9zT3vj/bzjYWWe0B2raJfAMvnKvNW3reIi0vwK/4llyVzlxvCY05OsVZBaZqOZtvSf5GqL5J8f
2C9KuNqvG/+Hwe9C7/Aqk7D+dU8ZDJy4RiO6v2zdmWe5W1yNQy0Cif0FmPhNfQfAFR9tgr1NdnD7
bLM+7Wo5aQXrCmJYImPhHjo8Lt4o3yUAyB3suU58xccctcAmqtWSHuEAotuNcYgAln1kEWt9Aohc
RSeQoghj0cOnGE7ivZSti0JgMMXMXwlUj675IYJ8YBc1ZIqJfvWGCn6rCiQ8/loky6U5TROnhMcq
PJtCY51S9d+csUuSsal8iNmgzsyVVpXXyDXmH/dQ+SwsAeUcx1tl3zqe3h7ex7DLkWfKeiMfQof7
mjeR/VS2YOy7T5N2GZrB1wAoQcKufBWnWUpHTklTKwzh1/BjzW1RPc17+2kBmjoDCoOc17Uj8xeT
tcjToIEpcagjYr4WyBmFqzjP/p0UyZ12DkoXTO7DZlEsm+OnUuxUPG0xjeY4P//P6Nols09smmeC
mwuwmF7/n8OXvdZC0uNP1QK99s/ReGF3E0nhneZFw2L2Upa8EcPc+If5KlRfffEybz81JyYVvGZ7
VZR/dL8km6JURS87UzACOkmzDiWfbhzWHMEDNmg/KqKvpP59l4bUNyCVmJUxXGbzH85IYdxMcbHo
bqLnaCRrliSg7WEF5ZfIzex8UEPWc9CIKZPFed4k3JFdEEoGVMNWFQuPeQw5E+p5Oam+lbftA2Gq
VrG25bYoAwTrtT4Xp44NAgqym53C/RxSOKpzTNwEAYZIeVU0aXFEDEMvKAGp7uor0kimdbpFC7cr
LHPkPdZuN8qeDZRsjALeEwtgjKWs7q5Tq5tBn9OubJYndGK/pxU+PBxbisH14Bby8uR6DyRPBrf+
n942zHAuNuZE7SjtcwKCbt6aU/QV33y4TiGaL+T7m7rLtt/d/KgL0gHWQY5IxKyetkBNCA3W3m7X
ncbnD4WHY57Xy1KhIFfM5Gwz2AJUuN5aJlXO8Y7vu40dBndd/uUZSBWYPCcP7a0OU1pocCxWjvy/
X25KAwnAXre/9nOvdR5tzzASEiK0PLgM6exbd10DAIJp7vi0lYVTsj8ioKR2zjDV9KX+KihXWZdA
0xivFvYgMXA+fD2ESxZ1IJPdcFfrRR9ItK6QXtsoOPBxziK1Saefq+Kr0Qx7qZjPAVpyzqIDLC9i
8xazWJKnoiE3xFJfSMAzDaHzEj1x+DMOwUX33pCk4vFUKeR7KxCMZMygKi4BjBqOZbS8tzIv/AQD
GaVZDgOrpEw76aDtiCRbltoHwaiX5qBa/yGQFDkVzutzM+uGBHkXEo+TyoOex5NDDe689504k/bt
KZdrIlmB1tbAtRjyIZWpt8lByadBUWDYdhg8fjlw9u4YydtVU5fptAWEun7NMeQIcP/OAyWn+B+b
TXXY/XfpAlZrjVvBanc04pd8DMHtcnl0iSXWcj+ssW0aguLVrLQBDRw2TlKzTCbIuX7D+Z06BYly
XuNA9xr12z6WNb1A6Kn0SxC69rdd0aIzhEYyvJcCaVVzZZJ9r/4k8dQ9ylHTGZDrNkJUJ0MgzaCu
EblD0JCql29qvyO+s/lXQA7Z9kXBiggYr/dWbfQnO1gwAzBgNqVULfa8oljBFyOOc1wD0n/A7FIA
771WTaHhnBgxNrWl+uLB6oKA7rcUwiB3wWk0YzlJua8fS983vjn9me06mMh7JDsk8yTklTmjwB4D
6MPZeXLNbsf+4WxSctyDPTsrrT0ELHkBwwKqG5O6yjeDoye9mcIea2BVt5/Hqg92euZD17V4oV9l
7yDq4x1DdQtGiYo/fKqWa9p0U3VuJZwHeaezc74pVitGzu3vGjKNmfVCXfnzILiwiX3vRxwrnXFs
uioISiJya97tl2lm0kjGn9hk5Td2yGg9fr51y7uw0DkMzHJz1W4gEdYlsJR3IpGbBbWCRBB04OuJ
+W8DGLajSIZ3AomjcVdVFbhKDVpAHiO2p4z739dn2gsGgiD8WUkmBC/b1sXKSLmCFEuJIsDg8rXy
1+TvdvNQJ9+945Ej0ZlTReaUybkenxhETWPKfSrZa5owr60ClffIshKgz6ewVPDiffk3bceUqVyG
VFTgO43SVAXDxIMRf+/2e841thZNCVohW3YZ/cn33mgYFhYCFQeh0cF/1snYWYxtXes2jkzlHf8M
fMSXdFYuMA6eNWvEo0VA4mUHpacQW/BkaGu/HIoyn1b4fkXszee1p8RKJtaHNVvXRCy2W06WHutw
Vv4aOywoRm8bBokHPYmV15OxAfGavsE2YVPr1KRMXTu1GAs9i6O6U/AwNCpMI5Z0LAoQVNauIdak
8AAmhFI/kSzXLL310q6bmUnXE99Ruve6Di9NqNeaqP99eHp6y27HWoGb6RXHB47UrmL7YnNS+p8z
eToRDRZUjKU3wJna2VM5z7bkPCofRAvcZw/kk+Tzx80FWnUarZC31pCnBVrDPa7gwAWaJOn6S4zx
h2Agj9uVPnc0jPRboGDCK6RB/KxUQr5nknd7Rp8JAEY8PRFP1ZpGmXFRHQ3IahKtCNZ4TX2xSZBv
/8KJzBGy5LfXQXTndnfV6+0P+rU+Md4ayPKvcgIoTpeH6+3hlxTmWYfWZvvRM+5qsMrQqyc6iaqM
SuXlsEM2UAORaSzUI+c2ZNMEa49WBpzngSI0yAydgwxHq1QM4hTJBMh1MeFJQi1OpfpG7Ul2rBE0
S+TS7KQfFL3MD0hd9xbkBiNrEIU8wju25+A5qLAvrG913rDqabXqudP9AWmD97+7EZ3cAddZP9Nz
JAyPaqo/9EoHPUa0/eyvv/AHTdLlqTBT1rck1Cowmee+t5ZgH8pD5o0kBGsO0zSGF1ynKGUaaIVH
hrhxYPoel7hPBavEMIzk0fHQGnwXetQG4yQRN8tgORbvTTpyjWFsZGy7nRtR5qk62KjEWdHsgeHj
80D08NN640ScLHY0z0RBSOL5UwG0fZHwDtMwsPzJZOSM4i+MBJaQpMpNKGZyy7WSIRU/BfndeIiz
F6hXshD/fLHeU/V6B/KE7TffuCsFUWvJiWJPyouZDi8lusjjV28u4OyNZYJ0iDh+nqIVw0Gk435b
RiDpkSx52O+3W1HVAdEgvSaNV1MAbTUS5SG4SVD3d7hRzRYmoF8st7maTgN0PcOxqJ0UwiqD/Zp6
GYNXCpH85tYrDL/1EebGF0wCIbQIj8j4rFB9gc7ZuCg/mVuns7oT9pV6SvZt+awpH3hR/hS364gR
tgiXBRbZ+syMECPC06x3dcNXqnlsFIoJzbHNoEsGdc5tflQbAPWrOmOsl+Qn1PKkrKPcVb/tRfBO
txYdEkFkXoc7HE/34vgchR/HYQUiuXSvYTfN+uejQpLKalKJ8v9NCD0q1xl08TPEvrRnSceMotgi
rVsDC467R1pAdu1B8LyaOQIdJ7u5UoLS6YMApk1FXF3I3MVsyRJYXcwKVOYAt52uEIWsqBsAslK5
8vaiBGemvkyR1lPGtb47wNIsphWTV1h6HmeoETZFvc3bsp5vLb/qUIBsaIW3TdinCyRSXDYrRDXM
nnHVMLebyMZlAxdp3t46nRo5sqhg2hK/bdB6475m6QpuS5tDLwboaw3ULAeV2lcebzG2c1l6eJza
CTTYvjG92d+iruiB3tN5A/NZWoE7IDT9WjhgtnErAdSofIEeWsMXz0QP4e74w8HPqSV2aLkMnht9
PIREbAXPrkCMIPnv11OVjGqvIO5GRGR/KErcul87OyWfRLwuuxhYBZ7rsdKfb6YJMj4xS8ogHZya
uMfmBZvnpyWsATVJ1/WE6yT2H5a3AdvesZ79mbBE+FFOllHrc6aQa5rVmw4L69qTzK9SxK5M1jRW
OUuIdkyF0EiWI9VVYvkN2M1NGsPsCn5UGL2W6k3R/T0Hm85Ct5hcA8nbiYj5VV6qcaNE8BiU/D81
/telXixstu6GEmCd7tsYU6BaZ/P0AnCWQmpWswq006t2zQNWkh+0jVKJ70eWBXd19aL+rzQzuNcZ
MAEg5FelydqA2k0DVGUkEfleE6L6zCFN3gJaq7NVAkagt49qzejC25hn1oYgZV3/8Ic1QWY6nwKg
qmKzjPXO46B7ccugy/MLjIsjkuiVm2cEotYcC3p5QrElEZV9nqiSp13brPlrYSG/b9GFbadpKN5v
hY2nL4ICtT2zvpyl7TBcivA1ZDXHdn4B3a6XqWcUPR1Ggz1pqHM6Zyt4JJJCOl8nmC333O6XLIst
WnsRj9a3/cia2bgGsvn/ZSS43TRKnNCV9E+Rq56n+uEIJGgMe1Ikyb8eyu185NX60osvdnlfYuDw
W8a4Qw07HRS0m0ziQzxuM6M3ZlpQmHHCnD7veKHQ2v+UWkRTb0A/1gSbotpBWN2YTqpUUPt/uwH6
vYj3GsCO1H3H2tnGrcqHTV3f5s8TX9BfRFwgH5u+FbNZVbttmZZ6gnOUVlHV03+ddDIB7B557USb
qjTwcBnNv4Mz5tEMNPq3GWKHOmXg6XXVWKjFod1I8wN/KukCskoeSAdyD1drlJTn0m9mkM46QkgH
FlXi+Cdo0HBLxk0wMR1me9TQz+hAgTkq4/7jy1TTR/R8BUiLW89xV7X0ZUi+LiVdDUni8jkfLhFW
UgpSpT+XnV40qxgyt/qLhnrp5x66clileTASC4MVU8UZcYz2f25jmy3MUsE9evYE8TcE4ipM07rG
y6vhU3DreugIPcvABXITfZPSJv1dUIX9cLSUJxXryELwRitGE70/5UgQVEn49b9ROnlj83OecYyC
5oxR35B+nGBd63PX9gu6CRbR0509HdHd8tUnPBXjPRfWosxmEAz4Q+fX/+GTMP3YDAkKXdJSlZPj
8XRExciiRtdTcz1A9Kfn45QFhME+7ihebOlhyqnURsrY8uerIsKIAWgdrnb2LTWHqxHiaAabvG2H
LEzSXxbiGWysoWfOkT5ioeOhmc+/rkSs0nmJhobGwEP5H5ueUFlAqUpwJ3LV6IiRQ1Ei1r11R2kD
TeO0mbw2X7mUKZLTAVD76A735CtIv/lqHt9+3cTQezqMvi7js0bPJ5pBoedkWwrbb6AwJbHfsMsg
WHMaL58+RiplJ8RQRqkRlutN1oXrFrRxGF5sWtygP29qJ2MUrVz3gfRYI00BMT/mOCvA9dtbj0CT
VQBGO03eX0iPHfltIu1ptrCY/Ms4QsitctKZHYRE4cXc/EhwtxnHMqf2Oac8hIJ/7BjaRy1Kb679
2apqNCw6KOg4q812SH8l1aQA8WgghZySRVMa4jg+0rThfwr6tqXs9Q7fvZNC11lyVljOkToN8KxO
azCv7fzC89htZkeGSg7hXveRXnCEg1Xjz3unDCmSG5gcGyBSnwuBuW2lAHmNs7HJTgycVeradj5V
0VrP8N4oT17AmKPX5g7KfOAUaP9E1f3OQkVxf2aJ8vsMxOXXJjrK1IiCtBZiwynTAE9Fkvg89WvL
xN89JG+760MsOs0iUbLO98WFpshKuFQRTsZgTUg68MuKGrDdnYtG8AWXbExkIxeHyVM/YzOQctpU
LzmoE/4HiKqhcsqjdAnJExMnplnv70eCP1Ny4RebvKEenm4fqvPcd5zzK/FlkYPyDuGRO4UE73Hx
72jh54T1eF9/nT7FgEPKbLOlC4CRknZd4EsrT+6+200f6fDNsuBp9TDCPiPYDL81AzZVQLRDHVDJ
e+sm6hgnqM8X9loWpYRepB3/O9djQwejha94tncaRhxenwjFfPfnX/bBuHuJrWRokBDbE3hnl+x7
5yRu6d2YorGEcxKVzD+1+H7PWXe8lP/X1w1RlsFiad7u15qwJ/ifHkFLDInNl9PQP2lKTU6WvsDl
yt98Iw5DYR20wXj+E1xSG8tsC/qochFHGPQxkKkTllDSqVE0msMUUGvJ8SG2AAmflajCAILwofwu
+o/ZYKvrBha67sX603mG/EKMtZ2Jqujtitlz8MT6iLltEX6kvYyPdjEv0tj4U5n8xIhiMWlPFwl/
OP7meoWrR/EhGWpX2DaUHnPm5DonqRtiu2DiJyVRhxEfA1+vEQt1LrCcAZ8VnIF9Rb/H2tnBLG9+
K9IxXlpS/esNVER+F9/I2rN+LTXS1MN5HzfNvqTSIkNfUeMg3w9XzxTtlom2NFmec6W3xyr8V1qV
yNvzihQzhBqgvXPvf1E6JYURB9/rSneZjxkoHYJNYGSiTHBylj8XLCSjkb59D+PcZW7AgozMw0Kx
kIRojT4RyaqqzvpGbGndUNgaSqILCSxsP/JBd5bPLaVdts2Wj2AsxjtY4hkXXBOvQ63XeiHdk3Qv
qOXuF3OrNvYIFVPby0f8I6rg5UGgjR0Fk3L9mH30hFzItY3jZb3LDjSaEAZDB4IiNziDVyLMxhpJ
bLeq8VZdjAefZ3CjyMxpcWm/Y1iaknKG/b6osOl08bD7DcpP+etPY90ugmKWttkzUuEizs/j0Yx7
TIyuP7PTb5lxj7xGQ6t513b+WqwnZDCfNi6754oHlsEZgj16FfzDCoxAOJWe8z56b0qiMrXXUiwu
LfOgeoogY8CM49clp/jdCrqinr5261Xpgt8hoHZCbzymK9cri7j4H95sYsbHe9HhbDN4SPkG/4yb
KkCFHgGnAcnyrebT3IlOFhFp+XsxxpgGmOaiF2r82gCIfI1bKWYrcLiBJsCfCMkqu1Fa16FHu9vx
kEtHFc381nHMjP7Dt1P9RfETCBSFecu6yTlYGAJTUQ5Q+NgfRwa7FnrLBBUcPruBHfPYpZxbm9QS
EENt4V4O40hk7s6iWeeaRtQeOe7MycGQVVVKk9LtLkLfN2Qc6fKDLIGAiP5TOIiuxkv3CZOx+P/M
tijmxeYuDqoBf8lgEENBnyJosr8ppfmjCiemFYvM131VXILcCGg0Qf6ehRuZAjiT7lDXTQDXOS8/
kL+IQoehGxcN9Y8ZIbRZf10PB/RZ6lFs669oql401rZuH+rxAW+BOMBawdlor/B5/8Yd7Y7cZUQi
cKU53ys2EV19snaH7z4mNhR7Fia+F4TJJjwtyobaS36tYUz4KchVL+EEVjA0Zzvg3tVR2Lyk5xBG
YYJvGc+rAe8S3ToGcAlY6c8KMVH+pmIAyvALoPA1Pv23lJiXWu0RP42oqEv4EzpUUFPhvWCPPVag
u63YMv0CHnsWIfYcRzPO3vgXN2Xiwy1L5zyQmQ0NzcD8vWHuNfQgpLTZHEdQGnnSxNU+MhNVeG1+
gyxvi7udXbWZIXAAPuNC/lbnPPHn/Y/vLLfe8DLr6bALpi7z1BfOkfZA1ExSunvPaS2vMO8K/79P
vnoYNVX9tS3vTEgN50W2OksSjQ2qUI3pQEgLVs4rBf1+t/SzPUjxn9T4wEJwOfYTV5HyJaVbU7UG
apk1y1m+2Z+E4mQRERMges8W7KicrjEHvoKfsOxOWCnP1600UfhfYa5OacI8ris5we+SG1+BZGXu
M8e5ts2SJyIimYxHwn8e16mp6PbWWnyf2GZH3Li6L3IHD5c0JB5/nN4xDnhpbJEWYzM68HaCj6rO
rUsSiC1DVgoDLUlZvH2zZKdeuHmKlTQRFtN0LfrYpfgFE7dQhVBKyWp2yQnS9Zs+TwtCX3POK+Pa
9X8/m8R7xhRufCkA9QMNHyc/VOyBA7ujUNzTwtcdeuXjwexXHlmfqh6JKxtGpqik2WUbPBefmULV
myQNEC8y3yG+JSGmFwjS/n7YbADI9HyHo7XJjNqIktz50F6IgS6DbpEIVAy/c8G6AMKRRq8SWFCP
BGiWY6EJ2z63wVmDqYQUYxjPIzdti0Y5464neGYDHdGUOxjxkmGeG3pDKeFknYi8vpJa1qcSicZ7
mUebFnNLjRGi+VIE6HlTTZdeFxjG3nUcXhXZuyFk//+frKeNbZ7qTu0a2VRcH/B++wrx4ifVsnOi
cKyeen3YYCn93SEKb6yIFsvJie5fwDOc02pGrIfy6P4X75IAXvmh615n684LwSmO1gVtt+46XxmL
2SRnsjusNuuyKqqVR0mFtl8Q+bLzXue6+bKQehjCKydtNMUd8diZNbY9EirSATYEfEVQKaB27sG2
f8YrQGBCGDcsw+I1jnX64vKIeWaEpV+1qS8Jhl1rCXcHgUYMb96cypRmN2QStSwYu8Ek9GSqfaXV
bWsx3q0jvXOQtMfGXkZOLbnio5Lqo3GTf1iFAPZKFQDSzKmWAsmeACn6pI80CksK9VvlekVheRt1
IdT+fvNCIUdASd//FXFF5MekwTqBy9asA4I2Jm/v9x7D33D65N4rRfjAMp5LTeBrfYkOmgb7oGmM
E5HlSgLow3PF+s3a8wXeW64gxaSXWLLOVs3gwlDMy7eoo8dZWxRuXqRLWdaWPnUYOoFkaj502q00
pqO6yQzqWph0Gc5bSRBoNh2ouYJrVN9/WRxv0b5mdgMZiOXsYeV9pfAuXd3kOTmwLNM6zQkbxKly
m2unDYGlubqclk/8HohhuS5GnmNJWayOOHsPzgyaOhCJjAy5w7mdeikQ+g7imNsu8GpVBc3z+P9O
o/gWi8taY2JGFAFV31DegrOe8vwMCoDSTrxJFNe+h3y0UmvD1CINK98+JqMqo6FsgaZyQcRNtuN2
ex4T94laIaRu7wo7F0h+9/80YaUEpwh6rRG0vYP63DpYYn5hNgJVNiLoGNkT4QKKcOnIxLutgOjm
R/EzlxVl2HMjKykNxBiMEYeouQlTSFd2UsUiftQNaUgpbypUadwnBd++EOOMXUUc6P/GaSa0hWh6
c52Ehu2IMrtdZqjGTUMB9xg/zMhGtN52YZYZ7VCfh6LobvjvtYcOpCZaUcd54BpbXAACs51xOOI7
V0w4OwvMLlxmqnf6+uyrm46UO8w0W0GLCr27y6sTRh1w4n/hggTdUiSMmhES0t9UxdyWLo/4VATG
tZkOVdYVh6r1Oxg8PxWNhchJqQzM+V1vDEHaMGhac1EudxJoeZ9Foz2IpsbiwOUGfJoKo36DvNfD
eCuE91shRkw7sUg3b6a4VLeKjuCtXvNNPv+CK0NWseXEfNWDF1T/vBPBdZDaQgGjdVM7HfRmslxx
owv80YzW5DS/e5NbosKQcAtzMuKzsvmT73FqKMBIWRcOnkm7bjo35k+KxHP9lBJdxSOtowKoe1fG
Oj+RHZnGmdGstC2OoQ0ut7SCTHJqca0NiQNJrfgf9KZ1VxR1vFoCK2Hvh2SrYfXb/FEv0ylj/ouU
2H5eTueczxvo5/wzpvFSV3JbwAyZesr+F2zxGYqSNoqGN/w/Fz4iJInic8YVodF2TF57rDBzuItp
9GaejTw/saNBrGrs4wsK1n2f/SU6s0QGvZQOuyA4jWepw3tY2mBmro31ZM7MEwICfW5LGkoUnSH7
DRIPflT0KxRa28mr8qDlmE/HooZwLcQ/BqE6JIfBMQ+ebw0LfV/xmeTDG2fDtFZIKMWO0FRk0PPt
V/sGuQ+K7G5h5CSHUcG8uPOesxA2nrY781hep2EYsd02Rqf3EpUGu4E8i3EWK3zhsOLe9/J4nbCs
dE3r6cUNXQmidk4SX7DfSjmPFkDexLOm9GzTPlBrhvFHPx08aFHNfjtc3u5oab6yjg1jNqlSrYnw
t1OAuaIfxG6zjjzufIfUJUr2jyvB4BqSzyRH5bCU76x/q6xfRFmrxLAYskT4oLwxiyJSsVX8CsaF
rZR1xT5dLysBdVj+IQXns8yo2D6XrqULTd/08gh0dRJaNZ5Y8TRDSKXvx6BybsBYJ6IMGC3Q39WT
f8LRR4orICQMgXl42uAC71fsm30tcnJODOP/stGJd88L4ZoY97sdtcBSwTjTXxMw4/DodSraSmMm
KYgq0P5LiHAfjRsrFUVepW2mpc2icOfn1gRytUDM8+hOuQIEYC1cyK/kFKpMc8xWrbQThW6M9S1X
oYsA13s5PZaQ71z6+8wCtvsWwiXnYRCY8gGm00j3nblv4/Em3DWHJomBFG+WcnXxIMP7CNClx46P
+9Vt9UEgYH1Aa7aeCqAEJdLhfQC4QDDPyKje4U1ZSuAGS4VHWXbOmxI9wNyP4TQPdZSuw7wGENI7
C8KRFUNZPuRlRURN3XG5fjeGn/tdjLunySzQh1xL5BThYCZmHvJCpjapvCTcFSrETWqcbMHumhsr
iyPV7meu+gkUyrj1rYFMeKzHEZKVPWtDOWXfQzqO8BmBIthG0zDSZ1DWOdE1hGNrFfVqa6jsn8L8
3g7JS1mHUt0bfSxIuBuW02OEJyaRhjA++Hs44FCgdrXZZqFYT6WvMNPenMp1ZFKK5Nv9X3ewIJKy
OgAWLEqaBq2e6WX9aVgM5HhRUeKFE/k1Z2vI++qZeTuUyP8aLIZG7ktXQnmzCa6Tkkmgcdog9p+F
mpNNWcjsnDetuvdsUShGWFCLJ/amxDVtI7gpWealtaNnw/1+IGFHwEjEiiCoAQdqWSJH3vJex+31
57NaF58IwdVthIycncqNc32wyOgkfq4/so7GqKNUn7Mb/t/ze/KrAU0Wxpfliw2ttHhDgOAJLVeZ
dwIruPzC28Vj7HRRMzItdeXrSBPafopAKIeBeAUPv7gfrvqI/SOjNV2l2cj8zJO7j4lmQNn28xAx
uP52Pd1IZW0tF6vb4vqs8kbbSLEu+O/eEWP5CMZfgGtPP3ANAAEB3bNq+kyuoO4ET1b3abvilhCD
byU7tOYUxGQ/aHWE8IX/45jEeH9e6KaD5kA27D4BdQGSjCTEc4koAYrowDvsunMFsT/cZj9rs2RF
82HHwAoNIGllKzjKp5+YD+pjhOLQxcDN7rZT/Gp3CCUD8/rbQ+7U43cwwc5JMTUCr7yjl4F+uHX+
SL/ucnpFGyghVeuLxGjGkp44/P+1l77hpK7QaVk0YYmDb1uW7biUjVQLtB30YOihm/tqKU3Cg/rO
rd8Ayf7hOSJ1O5Z6SXZX6Z6cmH9lmD3p+idaiBAFnV0+Yj3I2jgensj03RaRrENm64aK+HCHPljt
NNZaPkKWe9x46xS7t2zgcXJOXW+/vTzFBkYd+ApfyR7ZGMvPVJ2XY8LmwRmgxUVUrjJuNPZNd/wq
rDj5WqxhXlGvfcx3Hiv6uq7nJf+/3S4qkUlxb0sQL7jqxAn4Tiv964TMrAAoqWxf50ypV1B8nN30
TScxiiMczjnexrAUGYaSP2QdA8OTOdvQip4PiyEsL3WW7PqSnCU9UV99R/s7LdAWfUcv9fFZtJNU
EpjNKRV331x7X5vt/mNnHTiQz+oCTe8F+nTB85u8trqasoV7HGP+Boiv5c1vFdry0Td73abpVD1z
lkWl2emeKiyzYB+/ra2C+TNEftGReGwvH1uPATL5xH4el94CHWNqKegm9TsbHyyGJA+1CV0tuOsv
uDWsLRWw5LB32xMmEWVwMFUFO7YhPN/EwxAKhoMWOtRHwvO1a9mgQFDQvc5gVVt8Njy4SKQPb36C
xee7KEmYCmPUlYbSrah3Fb1/52Te6T68jCwtHHRHLtAp0Hr3VIRFW98pntlrLBcPjyMVKXpNAfoq
jQO7iew2b/rRyTo53rMq950mdBJX0AAcYdqzU3H30FQqyMDXgWzBJbR5bfa+k4Ah5TqeY9jwF+jf
94Yp4PS/kS4OoeiKtj3DVp8q9fbsH9QektUqDvOqF0+XKJeO1LVI4VijOKF8FMELQ1eIboBIpY3J
scftpoAgXXM9jbrXHf7CONwqI6OU9+DAuZbGfs3//KRO2PAMX3ZkVCwEkKDwxNFIHufiDMH7Q6OD
N8TBCyYjDXKoEKOd5XzO+2VwDaS1EvJqQTgIQioRXjAVHkek1Tb5dN5aZ6L3I3xM+ya7nEX89yQ6
xP6v7wPox9G96EeuksGlhA2V7vcDWenNyd736Cn5HKPybT0wivD49SaufRbHdLfiVY+jY3eK9ufc
I6kGtFn+dqunZeO9D+J9VU+G9au9DdC9rrsz8B+mVSz1zhwQxE0j1IUdmvHVN1pzksKewDEtztZo
MucY0p5kcukSPnEkyw4xe1p+3QBlXRB2IOM86eo+XC+8K/UbAgDPI1yV6pN5WBpOYEQ9vGXaHTzl
V7Q2bb/P3GjcN29kgmA5aag995Ja2/nI/nYbFK993ci4ePOjMYbhxyu3nTQQD+iLzYxPnYtqq9+r
7dr1woEAOxeQMDzO9MYWUsJElK+V11lPSoyXVGOlUDUqiw/EkDyhZqhgwuZ3R5td95q+zd5Ciryw
50+DZ291UmiVZN9YN/wxYj3WIW936LrdJOUNydFe4m5wWZ3spwrygJk94hGRaP7G1zhBzblNp2z/
N7oEgJ2gpeHHwEYjRpW8/0ysf05gK6kiT6cWMaNdCjdisMCXj46Dc6qo1R494lHE9Qm7GgggqqqN
hXRE0YBd0+PSlCPSl25RrAhfeVYiYpBPAvbd3DiRJeuorre7UqVrVN0xUeHJufSumPWuIXVgC5Hu
O39TG8JZVXz6O9IHXGxeAHb0hahwcpz+PFmXxXwWgeNV1/0jSw6oYL/1fkbpx1txv20nTJVrjtNJ
GMlZA2DNuIdq+K7wUusgYlVu50WY54ZYllqESqwCrE97gMBOq4kI1xG2rQbC0HoilCbVkiaiXZ3V
dvYCch3rPIC6oXWA6UC+1Ha++l6eO0BcSCDL10uoaUZMZ+uTwNCfpdGNuzrIi51HzaBCPCUQCtIa
S8ZCE5tqmCTAA9cl/9HB7QWOhEZqa18D2jJ5U1EwM8RWJstt+j/QaeFzZI/NCaVhUyY6G0INnuKx
MWWS/SJBzU/FeFo/8HIQmwhcRvrVIeiJxmS5eM0uOXpPODT0UZ9N+aGj9DTu87/g7mFbrdYTLy4K
sxInuUSK263sJOXUSbTnvhUt4PHUg51XQNueqFy9fDxmlZvoNtB5z7ZRqcDBL+p7Rm6DoIbx9jV0
LEQAVHzt8DL3w6tf95KWIGsQ5kiQsXfILGxRjdjm/IF2EsaQrRjUQwfOO8Zf2NVMq+a+xg7nKl/G
oTe92WNexWVnxabPU7anax688HavQG13tjbi4wsiHVO0O9xLt0djBZL9zDRTlD8O4M2TULOohNHx
/rrY2oeqUnfiFhR6ucAkQZ4s7eU024oxOikCaYvIgfUAQR2AbYc+fyt2h+lvoTm1BVaL6sDdmQpW
HD+kAs/5o+uMDddaodeznUNsfLhvLnlZ9yak2h1I26bEoeHqiXNfmU+TkdY1XhBnp4O48Suuty79
1Lm5pvTajhUMkzuHDPsONYQlvnOC49gvwATyduV0QruLU+QRG2UsOj3zVC6oZN51tTtn/9snTlVv
kmE0j5tAVwJj5XRgysXagS7K01Bds07liHtmVt657Wp5aTbok/vQWsWUmUf9TY/DcyFGNXVU/Z/U
KuAKEjo+v0KU0N4Qu16sqzcH9xyKSHskxCEYJZpgAbAGIaL6E9D257mX225WDHRcK8Wiq/UGXJ+j
R99zmiZvboCf6aFrgyMWrKU4M9XUI2di5diJwUVBRi64DSQCOK4iZmgxr/1dCkBmJ/L8biEyQjcn
TEB8dxWBabLcfnkB4hQtZoE8qiQLOYtk3/QLf2SZFJd4S5oqfDOZ3thdNqAXp7cxL8C3EyimcBOK
qLjS8focof0+FW3ThR1FWGJF+TNtqi5eB994ffvlHzl17rMXtD8iAsvYWaushr6oIUFX0MKyKzzb
yKLo56vUoejw9o/6PWkeU6x8mt+K/bDZXUpX8WO3MihumwksrSzZAl8HieRtXCZNEyFXR2WdCXGT
PvOTbVmYGSOj5hLuwUFPCc7+dmenzlxBnzPycA6DKId+XqluIZ7+Vmc1N6icLaY7oIae/CK4FEM3
C/JjqCoQZydw+ugWBJuYzM+oSqbIF8LsjEsAKALk1O0sJtp6OphMwSHt2Qb/ISPbmGsCYcy60rxH
LvswH/3pSgIyppjSnDmmgn8YZY1dqUZIul+T3q8fME/K8uSSBURILkt5WQ6LMGOynLAoJ3KW2CQj
4weOgVez2Zieapm9vz3aqJ92fXbz+5533GqRdi/4bNlPVcuCDHAHQW6TflXOfVkR4IfQtBEbcQWe
mi0fjftuQnCwbAVqmeenfuKVpVrgm5+JbV3rst+ojb0rnMVWwCxKgOWLkevpUVR8HZ1xPFPUOmRU
NoaegmhVuP8w//PxqXndyCaqJOwWVwlm9K2MYvBGSTQSgcbO283sq36oaOUGEpczC+9zSZv1Sfhj
QlzrjhBT+1bn0cbVarhYnzznORJbHB6mMJFbzL9LjV65hKPvSjWDHQalVWBSi4pKNlRimgBx/rJk
56STXb9To7NGVm9jq/vvuSXmQgADbUnDmQ3aPmRhgbXwoN5+290KTBxqb+1bHal52XCEjIIZ/A+6
uwjUdnCJjSRNCLvFm6CwlvCIxz2O9ZD81zF/7l1/A8keKTUqV1QfB00m6OywdOY62CBPZw+Lu6gb
Duadhbx7lSURxQu5IqmudKQx1ZdIEHBNK/sbxPzGbL5RnK0zj2WWlGkhWQ02OKZCupWICRNQTnMC
I0yEawQeDrfXmlXK/UYOBCGOnPZhjFvQ9K7sYxez3TJO9EXj5FlaRGYds0EuGhEw96DvhFWBstvK
IaGyUh/5lFFqYHLiWgJRemBUfHadlmx52raqcg4/tfmJClyu5OtyTt8bhUHPvGifiQq/BXHv2wG+
EMACE3Df10oX0oZodWEZsnVi1L7mY9OvrWYR2pRJI+htiisNFXejb836pcaR3bzUpXOkdGI6q+kj
+68LlieZJHZRJvrKWBmwKb4DQikEZ2poctuzludrP27HyzL9BcVvaIc+0EdR+PfhUTqIcs/hKjNy
ixKrzttzAl6z85rHAiqOcG3nwQxmB4Jp4C6OOclFtxvRk3ka9vF0SXioIhvh6ddFJg86dGpQHHio
EGZ8jaTUzn38z+gkW7V5PLGHbCo3k8UrAKtNW8S5C9mxd1pyrcAC2ZPPuUxbRWuTe9T3VbzhwiDb
PkwJoRB+Y8b/hJkNHTGiQWvBHETalS5bnE2jN7xZ4saIp/FyWcL9IuM+Y4z51PUK/JVBwmT+fmqz
PcJmdIyjVEas1OeMNyB4RIwr1P5iBQ709xOucOCy8USvchKFmzHHsTG3nneWYhpDirvA1sQAHphi
4chPnW7HXU/nK1Hx9Tep4FVsfL2ww5JAP0hMWI8hjzFUoAY2iQeGIsfqJcUjYyzBg78aGnvucYM7
0YEOOOF6ke152VPuv39mbF6qWwt5/9L7jh8y4JU+4O6o0X0XUDA3HQ3y+i6GaifR7Vdbv8J2nqsX
wljG13Z9k+oYeQ+zuG1xz0TCOMMSOZIzQJ8waHDxY0DNhwQ/qQAGwy8IpVjlMaX0MHF5PUBPZLnR
FLIdfM3uJc99n2k5Zg57X2ihgfgTVULadkyLzagyyJcknGM/USKNPB2f+MVQW8XtezDCp6BEG5Be
NC1qTu01QVaoqmOET9Q0yq0GPNrYlRAz0mgG+S/I2UdK7GtjGbNNt7Llnti5OryLFiT7PmuUDAd4
BARlYyleVEmxg4GaWPy7eDGQ9wTx451VtgSqxtAliRX1MM0DJQMX93OHQUMw1cfKlpWpftGvG1Y5
z9wFDAb+RQCjywgO8OdFEJw6VolnrOclURxPX67tc7fQgSWduwmCG0F4Xv6JcsdnNo9MdFdfEsMT
Tb01O1wxiRdo85cOU6kvmdzOrgBtUCUXJlHlhGOWYmwgXJt5uGAYyjIHjI5y6ptlVk+gaTrt1sEQ
QNRBQT0jP/toyb6IaCfrVq664Iomky8w7SGBXUMtOfEDrBT6e4dx/6moZAubJo/W32HeW+aJBWFx
XPrH2ltZn5Sc1CQABw+NXffLw1EnWCj1zCq23Bogv6PodSgz0+Cn5o8nkiAQc9wQIGOBTiPStMB2
9J0RfXC0iZ/n+c49Z/DReNhEbi/AjPI4yBjQNAwtWxAATCNIm2aXdmYingTQA0qpaqJiWGsVAqt5
Hvlg3sJKBr/CZIJYlIW5BRqXTIFdV7fC/V9GQnuAPJkaNzbzTX+jpbfie9jBgzA9qVjwoWBt7Vfq
ngc/PrBqllb/cFZYrnQ0WR0HmbVr1BoRBJsZ0zA7iwenE9SzElA/m0JQGS0Nppe8f60oJ13/cShJ
H1xtodihpaLFCueWYvQmpvAv9mD3ZiMS0DypFgq35OsbCanrYjogGIEJV2mMgavS0SRMMQE9lYTv
OFHhaMS9nEbfM3ZdCp4AyBTgVd9XojSwkocSnS+QrFEHfwAbA4YSNcXdgMoi50UhEaR7vkI6n44g
wuRL4tjgFi+RPSYS/FUMrDzSZ4nE/Aiqu0JXKb4CGQSIO7EtCnI7wHgp2lkY9USR9F0W8sMDk24b
2kz1UeCyzz5ugxHy5Kc2nNgjCXwiNma5MArWGzX5RaB/qLFC5CHQd6HIzbpSqYs2Y3FQZMAQfRQy
gcLNo0x3VjbtNlF4Zp9D64cYN3e/pHVIZHC1/mXSgz+E29IsxFgfWHqcNnQsG8hlfdO4++VodGyr
aJQJkzO1kJxn/VkanCgHOveiI9+5fpp5ElF6gCQgJfUvawGJp53NxIkEpgjC6S3cqbNchpC4h2Mt
HLUp68cWwSq+A7pEghLWlKSVAuhGH31I56yDfAt9aEuW4CbePFcotZKVwb3UzmDSivT2tBZb1VVT
6T62qOg7use48O3ksH29PZd2EOEkAqc0aWRCz6/rqcwwJngHAIbgf6H4LbFlLkRalNfjHBfy/wlO
/Ooza/HyS4JB35Ncir/dPnOki7Hw/a4gBNiG002MP2210B/6+l7F2MxNMkaMgnmkyXoxJZnxTCOr
/63c9QfOuERalBwqXpaYIIcJGBSt8bpJ6967MB4Sx8E24GnNUss+qE++MASvC90U80pbj1XzdjTN
uVdkgUbOICCkgjXb4VE7brPWm+j6pKKyPGTyVXdabrkE96m/8Z7J8wc/uNFvLGGD2aO9P85+lPms
t+QgM7/UeBlT3m0P/91RzkiydpCaFBn40fnBgMUrfhD9X171TjcSP2ePFYMVgPEydyYCjJQMaqqQ
g4kZ7yyF49D+oHYkFsz7e6oUdCf/BwB/ZRjwMBMtJIhp9UB2PcTLtlnPkN9i+FBPGOv0i766iHE8
yDEWjb2mYYJ4Y8qNl91SF8v+Wgl+ksQs6RW7q93gjlVteSv9LdAsBf7wDUHuQes0GqfTCeiShzx9
IKqM36pyUZwgtCHx5+dnPK8MUeCXxEN+xbXJxh9Ox1+Q9VRW8c3Xlq/azPWDyueB8fJ08ixpjPnD
Wqbanm/NNbkTRZ8Xp95m6SwIsGSvcrRm2HrnwBslZFW1UO0E/VMI94j4hG6WMebC+zDXD0B7kCS5
rJhZBUAR83el6faxTEzI0KOtC4VM/D6j/7Yr+hKjnqswXjxEjGijZiJE7FyqiCu87v+hycRurYkY
xcvLi5lI99fJbxTuUiXq6SD91b/3LllB9K64ovJp0zQNqDzq1ZoWSN/4gQlpYFHHxtEU33UuCG3h
0bbdX4AIT4xMqUlGih6FLYzcuiOMPnpRsxZgyyYoBCnDusWCkCJA5EHBqZbmycieiAXYhhcrAo+e
UwW5jRrLyzC8qBtI5v9tUCZ56IKjOHfnhBL1e2M7PqOaa3/qpjDo148pscDoah41OKd6tGCxp3ro
bD4hAV3wsyHza6t2wAdKXKtX8MWhnyyEHFKsjHtvkDooNJVm0NSq0DnLxTFAMt5bUxT4EcgNhPbc
Zxw9y8ISOAuYzZk/DocIpniLZCvgIenzq6ms30Q2vNIkoxw8tRgpQM0Yq/MUyOSy5uWCe6fWpOSk
Ng4nJFfpomZ9tsUSMnyY/cuXSrVE7RJIuZVidPVbvvbgCgwqwB5DWXHEBMUd4BrYs/mM5xQVDCS8
9bTOjkCw152fje7G2rb5eFY/rzcIkzwYyD/gMPqjbVtg7IhCt6t/v/5kepYnwNJ9O8nIGM/54Li1
5LpW79iJslNRvlYJa5J2KSCIny9TPEzB1sjpD5iUsWUqLTE25Zwd7xLJXxqJg5S6FDVlakCTWMdu
RAb1QbYbWhvh1Ok+/Tv9G4ajwKP675rYq0vmVSJS+vob5abWbUWRXm9yDuOm7cxo+MskFk99fmvl
9OYsKkrV1hAPsm7sBcSg1CFMAkyU96PiXoChrBUEBFzt9cbLFOQcinP1WVAINaMtUND77pzXkFYu
RfoDgTLMToPyDOwUHfvRioNupkXRZwdsSSQG39+lrkpAnIKYa2pGkzuK9/wiUJK21O8B2U8QY7CT
rfqhCZPE7/5tvQ/W/q5GtfqJ2zNOEocRgi0KwyNkl9oUdRp0yUaIz/2v6/YodJ1ylkCz8qp0vZ4i
rKALNWnCyQWjRqAKg3dF8w1FlaGS3JQYbUWkI/qYL4qZeP6LhaJAs9KbaG1cy+DcAjkhnVI0RNYv
txnSsRpvDaMA+Mm4Z19FkSCflgBqIkwApDeAu7KXLPqcUJWQSA6YQ4Ug38JtowBFvYcHrNqYcYGr
3q7xV/sgKGxspTym6kOkdU3JjULSpf+UgDyLIpjZJ/DSGnAbwsmaZ6TEuCs/11kfFSy7tajmwAYQ
vmkEJoXMThT2TzBCXb5M/8gJbIHM+GjuhHW2wX2cIikWZp2gJB4ZgPrLmifTar9mkvzvMvEJ4XcS
mpsU9Y02z4BdTb7dmPZj95KDvWIWS0SBQZP3DD0YZD1aqYE6myCt+JqF7zqC2VHrvl2z8rfN3+7z
YTeLyvWYYLTYOWpkezMYsZBIdsFXsIUQf/yysvqRNEdxoq5v8kAkBnDqtK2xDp1gSVD5rCTScfFI
KHvyQzO0aFjkIhGEEB394kSLnyrv8pICiepOct1J+qXDbtgQsgv64FwCefkdXE7mV3Nw9JrlCnMZ
TOPJMT6rTkOc892yIWNDagZWVz9KD0aKDm2Bszj6SMIotV8TiPTl5XVphbQXje6T26HwFeHm5Bnn
JKH/uX4DM6lkcs2U70YGiwYadiu9CRzrskLp70wnlaWhneRzTZs7Q6VauvcwRBDbVOxb9yenKBIK
L3eZi90XapkNoh4ArqcmY7POTzHw7joz1tU3Unxu0+ewjej/F0+lJl17gsY9e3AKpBzFzYSsOYD0
Xk058s+3lV2NcoAkuNAHbdUM1kqa0Z7ivmEFsfUQhEqkwWgZfbY/7u4zGdKreEsp/88JUpJXVkgR
SywSpgizqXv31cIkhWKoN6pLXCBxUuQcR5qikbuYt9xbUjfCp9cUb1ivsF10vhv9wHIbZXDTofD1
c4S0aN1yr9oeHuconBIVbIjmytJ70M3c/VGbt1mzp9sIweZ+c3keBfyhYyS+9ny/FLyau2BSgAzt
74m+TEeUiwhBSqGanb/ps17NWGCpi/GSdFjPsJozOIQzw1nkXaYzthUd3He2lYm4DP331lA1ooJs
vkQ4Z236vxND6aw2glfn3kibbTPg6b1opwkiRg8mpD5TqvSFee7+MvOumAL3dNUyaECAaf7zyLWz
zAkmyphhyfsrREU11LeiA6jlqfPn724zVsWDeeGuDPP5BnHr5xUf7r136c39ObcFeA5fGfWDj0cW
5nRCpRN0TPbcICizY10amH/zSvwGh05ksStc3wo4aHhU1/Lkh6vg5sBmCq2vanj6nMsrkBgPqQjj
hUavUGzMZTJ5MGvu6cg3Hmk6Db/+v0g0gh3AlBP2Roul/zLKJ1bBy5lx0QTDnX54hmHoG1Gg7HJJ
Lvij/Hgm78EC3KuRhXcSYxvXpeIrKYfnMGns688n2DyKJB6+4Db+gpLKBct4R/m0L2eqbjJLD8XM
lpXaikCGDygAlwzt7ekShtGwJOkb1Aqxz7aTIh9VH/Id9xf2cFGTZzO0djEjuQpn3iEB/sVOOCVk
jw+MJrmKY9hL4cIqcUz6qZGGR7GXQ+3o4xTvcNScBepM7dYT6Z2FGWnNgteIap9khAwLV6YVUnpZ
3EhgSWcY0dmhk5KJ+IABUuOFgDSn5zalEMPsteXkrX/Vpvel4sIQe18Dr6QCjyWrqEbwzWJqgG4a
scHWhCMGayfhhAbgYleYQGXVkvxIC1881I8TtyNHvJvmd57S0ypmMOXFSrhLI5Q06gHLT0PjDGZE
sv1ZsfIz32daU7x9tXbN2REodKpueMSJDVoiCB8jSERHWhZ1TxL4mf6rIcQhzXEAUPgoee/czbr+
gBYCT27irEfvHVu29Z8a9eBF+zGa6W8uAhMV0P3pmFfTMBsBEsHUFtKGJnBCrTLDIOedTeyAmsJh
gBWeoLZon/LRa4O9qUhpBxTmRfloidMrMYzxOkW1eXAR51CBevyzDv+M/aqEF/YYQfkT7YSLNbT9
72H+S4kIIuD3Fj8aKNMPilUlfXaEa0QwYBdHAPjLb3J8tlrX9skrqq7/BkJ+e4cNkWx7cG1/4VKS
yRzbUnG4Uq4Csi4QatkpnR/QkmNvGHG+VOdR9pY6C3ikNkL8CchXHZ9vbD/vL0IB8yszjypOXthK
I5Ltr4KxBGM9+WkBLtvcazJSZaNMt2tUhJcA8jNdVp1J3AoJdP8ENgb8MTpOsxWWTYhorETq30FL
WJuVHlk0g2fcG2o5HHF6jWJlUTH4xlwaTzr8IR1Ke0I2MudmZUrY+erPggKO3r54F5z4S8IbI9AA
fV+/xnR8yQ98V75xh0fOjOT2aT0ue5b2n5hvNkLyMI7/JeCx+kr2qQYKODqCe190r4gqcQib2EZY
CRuoQikmaOXE8pCESmaZzdnaGKqtl2SaoSrATTJigK7sW4hQAEiv5m0005Ca7c7gXwu4R+R4ke+f
wrcCygwBsSxNTrpQYaVEHbgaONhWsWD46XbSbTCahzU05gB0cwPgxvKyecdCDlFxb/OIoQUjWngA
5oLZAxPx/GFD7fGuH7omGp7z/qODHoSeLnmr7tuwKCedYX2MV1YKZ79dxHgIgNiviaMgMcQLAsHn
dGitpl4neGozeMfiXepxKGvg+kJt7VpCusIbc1hdRnqPWDl0/zS+Hc6NmJiCT5GMZs7lcejYrLKr
D0T/f6wJ/R/2SxCZsbnMCHj0r63GNjK+Y62Dsg+JugDfhGZM15bdIEzRQukeAnTmiW1V388jo3gR
XOkf+dZ+Q4XO/tX2+sU4MG0/zcVMEh3ZFxluv3VMFgG1R82/+V7p2DSzkUIFU1gpdh9uHfYdoglZ
Gq32bAGrr1bbNFscStcRQmNHU7pcPdhpJEmYngHZAjLgfVeGkuGwmgiQmcnvKGhWOM/AvqPNTYVg
8KqV5+RhZnG71Is4Lb3bU5E08tBj6hU1SQ1OMorxapJ8k3Nri2TJaGAQWi3JQLRhnp7tzI295bhU
bERfwY/Tr2kM0A9ExPFkPxG7yZjA5Kr8e1kCyVr5AFm5SpAbTFMnIgNcZ6s8/O5Q+cUg4v6EjI0b
byd/Cy36OOFi8QHOdkJBlyuEV6WeLRgoY2DRCl8Rtkts7SNDUT11vo69S4k/IzwMI5lTLLAtxlAJ
BrR47W5JH2XtYXYmZphaL15NRnEjtOLoZWg2dnIAWG2R7YBEsI1cwdyJs49xCUPc0ZfmpsqGACyL
23VirjWO9dp8Yn+F0K6WTuhbsSePhs85OsCx7VDNS3gRM5MWREQA/mCiLmWIDq4F7GMo2gAlipws
j/UIc/a4CoSFV6kbLud5kDhqn4FXuA2lL1q0aHU9AOaj9TyaMlBg4MnCsrMbc79MANJT5g9futiI
OsJCXTgyNTWDkp/OrwlXQ82+wCtWSFFthM5YqVApEZ8XSvlEThhVZWO5TqWS0ddMBYZUk87+8M7H
lJiKnpcRv5IAp6giJJlcFsEdUGJ0ec8hVBkwg0hFwtp18Aj63Ku8G2GoeDF1x5wO1jDtKi32/QOX
Rgy4vi4yEnttcLEoISQNCCx+nzWoBpLg0SahKWZwW5fFG48QUU/eho2ol+fVe3ZN1RlZ1scrddsv
UOEIClW/BCO+7u6AUvravsNf4xVac+uceKR0BkYZIDqSbiydFO9HqiHOfbyyJwv7qZzZIBQUZCWb
d5wvQVPamxWpyb3Km2xWMx9W0tVpUwKkPTXBLTgcap0qnoLVVwhCTSdNReMdYWD6INBecwt6McuS
+Ryo5ogzxq7kzFqkVOchaZVJ5GXzwNAwBdL6Cc89fWXlQZqbZUNV5NVANHoE7wc/z0Lk9kklAEAu
jo8y9kBNIdpmo7Y8qVqR/f41I0r1jJqrxq4asHKN9Y2JItcldHVKpEQSUD27nrMWCb/LIyJdqrvv
9H1kkofK7hE1dte2G/8Q8NF0Vqmm6FpIlZfyyCkZuytYMr1eWv5Ho+w7fPKOK0AvVwQLge6Q5hE/
mzsQfvPR4xrDzmD4rGp9ZqJdDFTXiZJCoHDwO8V909IpGxQB9IF9I7pOLhbwo+lixRIIpeKODh3o
ef3xb6qBcKf5VV8kBPLU8MPTNqAOZXzTWKZU8+fDh5WtocMcXanJO+kHs/YZlNoBHsVJpq3e7IYH
bb1byLMMX5xnocCtpq/nAIimRfLWoYEuHgLny+kq5XUFedb6Mn7XRv1OyUM8/+KKkqcnYO8lX2gp
+SlpmGGNYMLr3ps46y6J4m8T8tZ6VQk8ZfmBIWSI9br99pJzvq5SjlR+weEyuti7DzamD8oQX0HU
vwraGHoISoLfShoxGdgQLQRKt/IL6gg2LLcCIiKtSBwL6aoMMMalVFKIksixeOa2yIRlPRavz9j8
9e51tNOkl79fpql5CaViUF+yBAcR/fLSuMRZkfta5HyE1voxj9cfjjVQri7H/4Zi5sYIkaf/e4Ga
pp+aH3wyrZFXo5LvhZEi+vAUF3ChqU4ng1p+Y6dy2CkwqaXA82vjsNH8Gfjbg15CjkmarmcgJulk
VsXW+E1af+u9FHKECs8rdLGqvPmBKXIUXTscmT1/lJ5LCxdbUS0V6WNPga5I74AhpChleLqf1ziE
a52Rk6Pt6D5BgwGhJIXwNQXj1oeTHOkIRjJ6Z3qqBY9ncs8lj14E5ZouwOO3zPmYYTW39QdCG+ls
kaWiOi+d7VNECFAY+DtWVeOdRKVN6atFJLKBRrIwemYGFHbeaMC+vUw4xUr126al90C/9FUD35H/
5vhffH0K/m6aVO9Q0xkUmIXk2h/4ys8Dd88BWmOlfXwmuj/91CeZKy91gQdKzzVUkCZk+NKrcbWe
rxVDbOH7e/StF6nC17q3T5RPjk5rW3RksX9+qm+FPN5HbJkBNJVxskaS6edWSEniWTcZf/dkxrcm
lhpgIUEtM0d92ryHRnpojQWNkhWA58jRNDrhSv2pPcp21iFIQe+LYRUkvFKsD0Q/+GhLxBq4pStA
o0KykMc0oHtYO70JHto1GRaKGUav8WbY5ANXx1MT99H8dG8a7KmFrOvty9DSssiWcQRRdBeXEUIj
pTpAQ7kx4GL/4tw9JintA48ngeYGL6X6wT25CSqnDnDw8AzbXd+RUUaD2cEVS8fmN24Rq5UpBPq7
AyHEVH5bVU7ZvE6B+csMW1bygQ/2kufCXj2Dhe/Lvlx2qRXvWOLoAaitrvY5aOEMeAqdTSerGc72
BYJg7x64S6BUGN1ShzjxIRqHNEvmorn/qpX7sWYT9mCv+Z3W9wUCHCjoBKJvIw5F2G/V5SGXjMta
MZ/Qb/o0zHVhG0bgij/G78xua/tLhs+07RGr0CklzjJa7UaIX9bP+CXcA9RWLq72++/LCaBxUYAf
hYJ5CRbR3kIdEFo54OummHHDS6XsATUK0E/YSIFmQqjv7nnVUEisTyKRY1QtqZyZmL34c7FnxSad
CEX7kLn/5enhp9Rp6RysLKKZevlBzYg/dLsgP+xtSpVEoPgYt9xHPBSuPyXgUOgxbhgSUaNQiMDo
5V3JKhUtwz+XiAD8pddRwwmfF2Bs0Mwv95l26sGB+ZhOMth/WLW2/OXUpHySf34wdULexrNrJ9Fk
8iTa+lI0m02ZJ+N1van+k/PcJ+UKN2l6EpJ5HPQ8rrQ6Ge2zLAGs+kdAHThpkRenLEAdLEPLrl/5
3/amd0LZNKSB+mJVoZGLjV/UhVMlTlAFsWBoabmY4FWPMPcXHw1CY0zNPoRHxaFuwSDPzZFQ9m67
vqp058Lql4fEcxTFbJaXGZIpnJ0KQSCPWIsR9z9W48UMwA/Q+jStTDreYghoLVAhY5BsEr0yHRmQ
CCA4VQ5SbE8QpbTaYRSpLiipBBVV0CTqcRtKafu/SWnmSgLIQOWSW6I4FVZXQX17/g+/xflzIGWR
MeHXnKvpww/OLKHef+h7EM3ywQE2pVE+AytxZPSYRy3qMhXzKiv2zjmjp30bb5r6JVLTOhNFOpJ2
Mup7uMQzfduJuQFnNATp8OOTuK04XNG73/5zKJv9zgDtUMFjmnZFNCgKkgz5gmymXqYQ4FVl7hBe
FalmaObQ3WAU/7vPkXOl87S0f2kiK7QtluYqM8P8Pv4fKhC+sN3g30je6qrcdTLtZaROsoNrsf7v
QO1fHLfd2j04s3VGDgKYpS662wm99xJz5Q4Zq1JzI+eODYMpZxiWyi45l1DyWTB5tzdEW11mx+HE
tEINqIyocqzycyA2qrYcBGMsoLcUGNUYbyClqw7l81NgdoBqp4sVxBzCq9p4GjZxMSyNIGmmIfKB
DmC+qIo2bEG3pXvommisovS694rOKvHobx3Kiai5vd3zLqqbrX17UVtumkZlDbI0etvDkIbGP49V
2l1Tap1KYaR/6aRUqhkyDMic+z6d3gACJTKsvEXwVIP2o2dkAnXrEZLy+nKQrZ+oEzB7bFN0ZJKb
HIkFqvltj5rIDRX7ODo4FR+qMadb/ui0wYOnUfqG0A8rmUWfkN2YCEnEab7wFjBT+KOzNefBnxgK
Av1mXkwt1KU2rWeMy4CcFl3aq1TCaL6kXHxH0gwnXaEOZmAVZGs/uH3CETgBH3PjvHFYxbVD6oh4
ipfGKrxAmiJB/RPhWfzGX2MRf8rB9oEC05oxm+LojY237zI5r5ToN0aLH7DcwErswurQZ5UAhb+6
LlgI1r3UK97Z20Hw7Dpu64uN7d01HE8IdJH9ldxtZbRVgJMX4a4UUtnwuFJV5jDwf2YPfP5cZi0P
d+Uj0ozMOMwYh5waxvTFUkSelhHi/Kcy/KYY57w9/kqFUaDIETsCJ/nyL0XS71q+GbpjZ5QFxnj2
3s/+BBwktIBjhrFBWWK6dOuhlpzXmlBeVawUHlBHRsxwAgr4RdejzcCBg69qctoIN8aSkqMdfK+L
GrpxD3EQEXMDsbUezvsQmVZFQhI4ZJsEDBoY3hXx22zyzNn2VE8yTthnLSDA5w1jTFgak3KcVvGl
+RqV82DnEMhIFRj/ojPvKCfaGjlk3dgUsJtLxAhlqIQus2/WivuX7lf/jQfWeGSjJEEVzN9P0sUB
vx5rREIE/q711rgrreP8M7yIeJyt4gOe+eYjeE9+Zwgd1B1W60uCimgd8h697Mg/oDa3Tb7PpFdO
EHdcAiFJNiYHc1fP7wup4q6k/X34uyyHEZFKlkbgjOY51Hkom7a24TUAt8FBJPmSY53mGd9GjWxR
nV1tmhcxSQx4kaOh3rIjDeph4V+PX4yIPdZxxLDEhQZzGKzr6PXeDk0UmYjXbcRUDBYRXo5JgDYR
xShEtkf6gGx+E8JKfiQ+YsloVMI+9Y/QQQYzw1ABqdByhm98mGIGTZeYL676QnWlpvNecy5yAewk
cyaoXv/xGnN/NY6WMxzqP5n8mFT7d6e0/ChPqE3k1W08/60tiFClPjWyX87cSFRIH7Qhztpyavt5
YIW3IQ6oxKYzBcHTPeQjVBS9GwWeU9Z16egiJoW+wbxyiF8q43DUrIhLm9ezIg3iyRzgOd2Y984i
v6wW/KkHkt6L/gz/NV/aPvkeYnxBETkoFx4q40KneY0cJAuYHULA3EpedvNmHNSKjLS+xje+6Sov
ROb5nIOHLZOj8PQOV1s5TXiUfya6ztUOMAl6z1xXt92firsA6vn7qyyABf35jXVw3MZIb0UWGAy7
KOA98ghSb7S8xupqu9KwvPUpGwRhwyVIcYbVGvYJNSENH6yiUL/XcWMTo5+R49GxPQrr3Hu1ELj+
fCHHGrzb0esKPhosEfbJNGOY8HgnGS5gf8OuCaeT44cZcaud4tphgRSJ4/oYPO2Rl2CHOApl4fGK
iSI4Ppgy6QraGJzyAgpSgMzur+fNUerlp6tXLrKRYCAilxllyS5meEPwP7uJ5GbBqKxi27vIFgG9
CNfpp6W70NDnpyAVv50a/7aNtxbhFC5pER/FtntlVTTDuRcsZGNxpDgC+Sy9AFviJ+EJ4WICiAi9
/uhEit+TdMWeQsDBnnFuR5coq6D2NuwjsSPK++wSoriHbmM8KxWTev10KE4Tghjps5ZSsoJ2lfsS
z9fJpZ5TwxXQvmLltGoAmB9mWA8/3unuB4/HLqTKzQ4YMO/NWJd7X9RgxEB5fhgtlS09LSzGLPft
dA9fI8DBXmReaMG3NfqBAirrnunlvm6AvtS+JDK8oiGJOr9/KMEp9KsN8elfwTahXjjTIrO55x6Q
/P7+36W4qAPD1y/hc0xW0JcchPgFAUf5SmIsebyqsK623XtfaxZvKi3DfpdjGUsQ0hSqvHuUgcG0
wewEuHY6aSR/yuilh18AHgBMZIO7lunWwNCfZcfzp//BNSJnytGn/kgVFDmTIEQK313TNVHm6Nr8
RlRb1xlyq21xMENW7aJ22hkg47p4OP76//Dia/2VuvHCgywXQwYmQ6bDQZlN+e2z/T/mcPxYgrwk
sAlQp3vyR4JyWmQ9v/joarHhh29KQDbDl3szZV9KG3AfSHk4gQy2o/h4o7yM06VT31EbfBeJ+LKm
Pfe8dsm18xT+zJHDEVTbhpDHBdt5FfDHit87NLkQwUnwO7aCNvyF9Y7blO94cEZgHF2Ghc6mWa0M
vG0O2YqB2Z2Sryn4ZeLPpkcGKcKakU5FdC6bW+9Kpjlj7jpmp9D3PQDgejwT2x49sTNcFtQPnd5F
QQMFkpVe+KzRHpeLb4bpSxc+nfYViffMduNmP4jGs84b62Mvju+5EaJ5eP16cdfqqcASNV6ch8We
UMp6GsYKPvXAFSfNU9Oe5zxQ9LjT7i7MjGYg6P4zfCJ6fp9vOPI8Mj0ElxgM30UC9bFipBe9eEUV
aKsP3LJpHopPtmhziTRrYtBIyiqxBvd0seScETG6+ZgSRHdRNxmbZN3nLqOyn1uX+5asK2DattPo
nTA4ac3d/mXFVVR5hjnOUTQe+DqNHm49/t+M6E9cbAGbxaovYKsLil6XH3gi4f9PdUzBRJTG9Jdj
ofFIPHH9It6wRToRJjemwMZ827HKk7OUU2u7Q6vcMtatwqzL4I31c8MXUpp6F1fGlwFBGaTWKhqO
9DBpJE7k2ka6DXflr7IuUIn+KKGlVtfguq332wppx8+izSh3wSEx6ni35uO3X0dtetiGsORG+OBU
YLnujES0XIYn3YyL1LpASuqu+9y6ZpcGrcfzZz9qGqraOKnzO0ch39NKtdxix4xiGs0OZNL1Iy9O
yldMhmQ1ibhTKRY/YTQ5+SrfZHR639PeDwQRUEEBFMMNS24PhZ4zb9YnaigGyVd4WPDcPwU9R++H
b2FWAmltBnYMTuqW0RDZaEXjz+Jt0luFbQstpra6LOCc9Djp+zzB662zBtXWpYN/ZxV0XueppY7O
rYXnAi71+eGHYtDvV1xeRbMNa/aDjQPYeUmZymGQkNl9UA3EQTgbxFBROYOXaOLsWThv94twc+7E
O9b8jmx3pWew2Op8/QZURCRcZKJVrazMxdEwq9tua5gBWgXcgwVBp9k3xCMrE05nDk9w2dhie4CC
7qFxDOVikw5XdtBw/LNs4Sz27L+eerZJsjv8oql8gvRqfmhjquZesIKklPbMdJ/N9+YRgh1CjUkO
OJ7yqOv3KSrPby8EiGYydAuUc9DtfXpYGMqnLQX4ueIgQu/2Rfc8C92SyxCX8Bd8GVb48qdOBumc
tejuo9P8CXFKYpe9C73+U8NzE/+Q3A8Qt7I+DI8K+r0WTNu2axhxDlr2gH1F8QdlB7Xw11yvPcxC
8FimKzIdbIdZGofAeUX/ByfhmkmTpJaB8U3/BspI0St58YvhPFIJD8z67HCOFMAzfVTK+zLiKC96
B8Fn5Xk5kjqRJk6ufa7OdGM4OZGPH9k1ojiWSm3/tCphjykLnAWH9CIc07O7/L4K22u+5N0G1fx9
HNK4rChl+oPN3VEArbBN64e7pSblbG6ZIAeUAoEPqCZKSHk1P+El09z0e5ykY9UL5F+f25zoiJ0r
yA5bHMg2LjWPu7Q3uzYn6gvcw3bZgTl6DqIV8azMfZvWyUjIG8TQTYDMY43uzkJbZ5Faxv1EWlGE
J3fynWz3pIhW3IFm+Fjt/0lOXyUjHhbJpl5ayZUW3AnpZjdh4GaljWr5pWmhnzfbQTMPF920Dp1P
QfX1b7HG0T6TYbPjlBqlqu+I4RotWIegc39KIxbKmlCZv2pnoKakokfLuzrpmwz02DrzwoTkzv6o
7aXJto6BmzKs5ijFVbc9kgyUof1lNkAjWdge3oeSiGMUVvj7Bcg+hLa75ZZCKmzZNI4BS1D2Km2y
gX2+xycL4Qbs2loTf4uaiN+Ptur4p1CdJbjY1efQFpNWCFM6oxO0bvXLduSlxy6vofk/+nFv60rZ
UDADdCusRwuEdJoAgooLKVtz1RUed9qDUs+DQVT/4s3qhig1bbvgGZn+gZONSofGUbS0YzCt3Hja
OoloXKwU5UMkfpouduReDCigU0Kt4HaOFt8n4Q1td6dIlcjkAHrJxGqY13exCdZ4NGPf7XQUwKvf
PZgPVvPBskyz98yqboB+CZiCCZe79NSmuzbC5b+okzhp9hrm2xyw9+Wg6KMDAJhq7m4Thkg6Ei4y
zKmMQ2drmeWyTgjQYbltU2LhBSI0ZeTsN4QK8B+XQOzHDObXiQKYb0Vp+zZBobMAcJPKOwQ4DMMw
0q1YbVFOzaIIqLSOOs970v8Rq6ZE2lkmTqgjwEgJcvMYMyqjsiiL7pXyPcHzYbk9fSKZyzacBQ+f
ucnt2XwzVBUG6QoBGUjHgfRQdBH/YGiyCOUJOGMtt837B76M6GuKPsr7bBishsyB94ZnHMuDfmIh
GRkjKKMBgpl76ZTovvrFMFOWWYFHVh9aZM5UDOjnhs0gb2O52khovDTZbiMjw8I16ikqTiMaCVhu
n7JChRFJ521HKBSjoJjIUAk244olPiYUJ54w0wbWXxS8S94EVUqgvwigdologynPW9t+paMoqa/Z
OPFlV7fgUHCIdQt9dNUKfmJa3cJn54rjRQe5/AYZ82GJNpPhEPIL5mao7vsHIdLtgruOFO+KfXFz
b8W1J2+ScLfQ19PEc5lOunuXIjrVBoCJaFx/l9K8+oWCt/7uoRez0KFxry3PyUbQ9s4vBuJ40P+V
aUYC3hvsWDhIDjKE6pv5UNbgLgogeIn8w/h8LdC99ODMDaiINmziU7CGmJCPSR8uHtOHLTyzyJg/
EOMw68185IugS+GnKYIEcyj1rME++gGQBn68HhhVWojO1Wd+aI0BDleH1rjl2SxuOh8ziVkZngQh
IMEirrtKEjc1l6L3d6ctxfO2+sqZ96nGL74ni+UwTv9JGNRueKsMGR3UHqmAnotGVlFguhx/iTTa
3OVFZYnfq9cujlJR1CdKant3ik6bCILhsJtl+oGqTWKjBL79IqkuXAhW+/iVeLzm9eFJoekpW65G
ypN7oGuePufdMtkJVTntppK3rG7qTIU59ssy2f20VMS65R7I+ZQV6f3mCStnZ7GpfUMzOHnR3K07
jaI7YeXwJpmgjKR8T7L5MJCet0KjEfv9g6vO32pjLHd4+mbxsrhXlqyydqrRF2wRuplDl2FweimB
3/DsiIxhoXCAi8XKoXz/H/NlzyaWyKHbZEWrnXRDVXi51qzjI9teON3G466DXuA7z7Pv+44LZpT2
6v2xqrciYErccp6R1NmxmlVYRLSRu3gjDPSJdQyUusHe0yQsCB4pTmrf9q6FNBVrL0PCRDNxm/zl
Syl9+IAg+Qd+LcorXUlfjV8Nhes0x7xfEeMC+Dr9Q7nFPp7oDQZssvq24JdmbVdajpmZA4bPjpXk
q7aKT8EE9IfSHUiopdaZ1PP6XbaZgBblyPH1sh4mloMHz5zGyrHpeAJiK3vrKGzFriLIj5A+V+sv
i9K5M47aaE6jplRshfIEgA4fU6+mS4dJ0TwkPFhqmBzXMKW+CgmUgAyq6Uky+sWEEC/JP8E1suwx
NpirsyCIxTvoUgtH0w2gXcqkdyWNvP9Hl2VdnYK/MuClZRodsQ0V+JZblhdQsbUSIwK8V3wXx0iC
A2JFPU2LGz09jOURiDm1Y9N+jBnYX3pyMxKydOGHVobumt0AwN5y5iO8OOnH62hV9iWsmVQBP16a
R3jN4Y9iT1T2OKLFrVxItIVd8gM+hROS/xyvon61DOH8kAewF9rW+YEHC0zUV+EcRaWp3cmC67gS
tQp6gGep3d63l1pNfniCJm0yXm+Vvfhz5tJZBVJOa7mOeem72fWpDM28cRwy4BUr/3BrE7mIA9DI
RnvOUm1zZjZ4zBrK55lcqUFnmmwajDaY/mQA0cLHqZMDJGirN2RGIzMCnoRdwISiCD3p2hS6MSoF
2sb6nqsrSg1pvJKVhg9GRuYS+n4L9j++KgAc+1SFzdcp3uaJJOv/1dD2tBadUAUjm8JgmnX+oNsc
wO8xoLhplSEllcsQEJ43CIpmrWW1E9xI4+0P6chJebJBzLzlx/kI2Jib36kzaaDvaLj+3+ORziOB
NrI+UFtUWtUb/9CSsVwC9sIXwTV9oRgYdMRhTk0wogIdm/xdcgO5Wt+ISfOiys0NwdatpZ1W/Tc0
MdkrYJm4jwI5C/oMz4DE/I4ZXk8yw5V/lilFwK8Gph4QyXnipt9RxhoGUKS/c6+E12tCFfg9wWWl
qJZsIw06rYF4jI88wslOtzU7fld0ENVfxc2p+Pltws27umT6umJwgByZNH1c8pCQzPWMX8/db0i3
oF0ocLGODZwXhRYNNk2T5G+p7Nz9YCHcN7eFwaXTnFu+bl+729+V4TfoysXgjWnYe/SDL4TfZsLf
VuPqOuOGyRNNMZIkfA//MiiH8PqUuFGu2ydvpBIDtvzEUPfIL+Z3Zn4ge+9pphhmxyP4j4SSYzg1
gU2jyAGbBnkG3ClnHZhxQcVqya2MWh+Z0d8dgNoIDWZOYrq+QfLe1nSoZ68X+vz3UAD5tG9UK7zf
vPOWmclS9chmSQYYyBdMTsSjh7JGx2VG+E7Q3KeFGDyd0HZhfsMXB5fBUxBnfD97k9thRZZlMbKO
c0RX4tc6WF8w5X6Qz2unoyl5pFXrzlSjqgsLKuebDiPrEeTX7NwfQooLHKXYKm39/TCVDAN6nEIP
0NX3ShdB1O32M6Qlj2XkrownyBHvg2qruFb1OI7iarjflgG/E5nPVFpYcun7ahie7bcrHDQbDO9j
c8apwCh6TiRnt9ERZE+ra76R20Co0ljOzpIeSxRir908eMQR2enSERNxFPmCNoXoC/BIJ4wrb5sb
SX/6WzR1tq5FGwHCvnT0/3fKqt9b/IDrufZT7HQ9IruDtBIpJpZhWItw1E8mGFTVcMkKwDjxgNwR
Jm6p4KEDEy6XWlW/4+z80wBpEgwKMDkFaZcLSLGgEfgjQI0jKhb3AozuBLbFYm3KS6ieJjC92mGG
5uiIG1OlcQ9MtpEJsACXxn/XzJGXB8xglh46bEUxc3V4eUznNYCWCwkeskabbPf6igoM18+RrrBP
AiDtGMlJpLizT6qntQfgi6GLMxqbnD7kU3B1p7f4K4T3FnmR2ZsWpZBQtYQKqAUnvf4ueEYtv/7F
m21sNr4OvgQx87AAVPIwdYxS5UrJtXgPW+gKapOlHDCRwFgiEEAKbImdW53jK6AdLKHyOKUgxN/V
Bd5IPZbAI1QS825aHT6RaTct9ZJnFglifGxL6rcOH4WcJ0UNn/SECs7OQkK6fABtSBJVNiKol19m
6mXcBrnrMDgog+BPksxe6YooJ+kSuAxb5d5ibwbqnk2wKGf57F1bC4ueKWVz3yAVrzUceZF/mLfj
gEvdVlRk4KIvTD56e2zKTETq5kjWEwx2etbejAtXVnYmcS2oGXdYcWBWfn1JgBVd3xFMfxlN67GX
M+Pl9/zIvvcmZJMnwJWgbY5n4441MSxW+1KdrCRXk+jQng5IeV6Oxi5/YjcGUoHFfE3EGu63OCr3
rATpJXBK2dNsRAuQf1v8nd8hoAm6iT45y+VnyWyEmlN/s8Q+v+iAkZ4tAj5op/12UMxe8bK6/TEU
xfm8N2Zz4M0uNC7T3BndxOr2dpvv1e/76V7zg70XWVrXfTsYy9IvK1joA9kcuOUxzNvILGlyywQ9
CYsQQajAD4k44EXXtaIcX7Xr+Xnr9ywXmjEO4v0MgOsZL1Zj6jCDebgMqV3hQ0U8d+3mee8l+Gdm
k3IOV7Bx6CZFaDZE5jQ0zno6+ck7ZgW21AtC4fNz+w1ZhVDgrG+yORTnAjtL0bC8f51K1oiTVgS9
wOKkSGP7VMMMqLg5kmPBlXCkHkOErfSbh/U/2mfHv1qHdk9F3Koj+K0MqHXNkJ1oF1xi8YFG7yfg
G7Gurd1JmVx666WIuA2P3QJCMfsb/8XTilMsIkyzfa5kubOjtQGDBba7hneC5gOGZPm8k56F0rJC
AhUErMXMzB6qANt1+Kto1CF8e1g2cP61mGDX/DJqwlIScHvtXUZtXlowZlcRwhPt68YY7hRSIzhl
1gIDXb+KyjjCz1xG37G2KamR0CC4QNA2ui6TNrs/1EfvTO4Mk1N1ObJVjanf2LOVSsKeVenUjV4o
/zFrJG1+b6EWY3zNFhmnjsHidcAky8upHWZy4mPbxmDaK8imcpgBnSgfwFVS068BzUVq0Z4Emz91
EPJIeK7WEIHad50SeG9WrKaL6mzWdeGj4rtXKYwYkrnQnyOuy+TFDlUNVzPGCn5jB7usQi3Wc2QJ
dpMM3cZrl9UjxXtNZL8R1qDG36Fp2PiVr/mUmYgB3x1190IRz/+xtTHi+ejw8xoa4rBZIXHdPzST
bC29P7oI9hOskqNbi8YMM7WEezT6Jpep53iSZNN8KPJEKHhQ70JMonyQ0qGU0kPptHAUcX9P88Ss
V5fG/FcGmGZ4DM5dWnPMwgRQ5jTPkaomta2fD3iU8xFna+xK4blXa2xZq/tZ8WvIlDjHRgIOVMxS
4cVIq7OaPUXuI6b7QYPK6WN+EeEnFkApGvzq8d4Jr8fxZf1R2KmQTrEs9dGhY9wpJmujJFfDsKEz
MDJI1V6aWu2vkNsqrtJgkcQsK4LP/G7g6x4HqTiuM8ASfnRSS4CTmCFpY+dsgyELHspTTZTHrYHb
n4h2rwhhJXGvma1Ym2TfhJ8F4ymqzsfV3YTFlZG/yORO+XowoDGrbaxpdu+h6W6twXZsYM458DyM
MJZ8eIoDQEkIYdU5bRdfDVjFy3oGjEbXbd/faq52XcM95Gmdz/U+v70OlOc65LxM6yrRGLa4Fscs
vObSt4T/76ZF6Px9Qm9FoNB02Ja9ZqsbxtNYepH7pA+zx+zV7RBdoPXFUA22jSW8kBAHfXp9tKC5
7cMNSAX/ciMeGJIQ1nyzn1crWDC8GvwUew/lZD2MUiqt857XljMi3o29QccNOeQJlSZ5jUCkyj7k
Gipsvb9aBE4sbaDGAB7L7nPXXvmosbx9IVwLx4U30kifzmftMgVqJOxCQj6xHUNyjlW5dvYz1f3s
FVhfBvCezDxTBfU8fhwY9UE1jkgOBVTK9SZFS864spj2CKJAt/hIRI+S33MiB6uGZuuKdc72NNKd
L8USbYOQf+YrWR2x8owWtiM8MFCwndYbG3I/coJGTUsLqCnZwQmRW73aBg7g3x5qLPAcntkCbkFH
cyAAmRjSgdcdy+lcnRoxFqYxBc3xECgluOh/0YBJ3RMFj4Qi5Ad5/Qr319rUIuORq0qCCJ0P0nF/
SpydzISqWP4cf9Wkz5NjsyIQdNBLrub5lABIcpJUTIclAIVGg/ptJ//uYHvz/6vVW9n6VdYW6otP
Kifz3YQYQOMO4rhD8JFeP8Urvuh/r/n6X5giDrOr5uU0E2R5AsSeBcpgNzj7VMto0cLYU5mPBZ7i
3qOB1p5QaWcIcU7sqjqCP07WitkKMODF22clGhVPKKJjvVAC6GPVErJGnncn5QbFeI7u6mILGNAJ
cHVA//k8QinIM2dzek5PiMoLpNnAzUb7ZV+PR8aQxjBEJ1aubgeaE9eUZnRk08y1GC5cSzmaDID8
k9ITJ+2wqNVmStOD9xoIVP8MHPPcw1a701tGK+Y11uVozbeiO5OZCd71Cn3gL/0TWVqbeP/GQFWg
5dXEdnygGi0ms/LLA7mzce0i0ejp6i0Jdq8BpMzRzXqrOXBaUj1buAE0UogY2bAkWhdITS27ObTk
OK7Qz4XuQ95zgpqne2Tt6eQIvF8uYnblZV0kB+c7pcX9XL+lqL3fbl6iH2Y2hcZ66RRCgBYlkT0d
srR0q7kklthvPXuoPkauDoWGOnV6yo1So6m5xKOWP48B89OI63ASQbEY0Jw4w7oE2x9QBAAoaWcb
xzF/i8rlhtv5UAiW4DNgzQaUsy2jJ30BtZn75CX6n2BUQ4WgNtVzll6JZ/xWKKZwuH65RI+0bnNS
p3fHVPc1W0AeLLATtJDCDQiQj683fmQxznHaQEKz54TfmSsUq4fVP17zKqoP1odP7UN36lzyFnyk
bPyZWKv5iys5KDunJTEiEKHz0n8ODJJktb1sUqZDJ9cQ3HmVBDRfzJgYXbAMjxYZCSyZ8KOlKnI1
Tn+2JSntQ/XevPji/ckYXtZ681spJB5FQxebDtjCpFvnNHSI4w5dURjywxap3ip9sqWJDwIsFpNZ
38ckeADUN1asWhKWqevsIaWGCMveRnszslQLhMjpUmPeaq+Nv+F93jEQdmpl5WyWQaNqugyiFtsc
G3QeSAKxGE1DxNmLxKpfpeVs68kaI+oKUTYF4xTYs9SeL3lNfZC1VBICjR06HDp5GxdzxGslYgrs
F4rnf4BOGGkN91vg16ZRvkSWZgemTvQLjQ5iRLGSltTbWx+21vkNDNfcQzytqxSNnc/1RIhb87c7
gctTeSUKO/ESqD3E7/4dNVQvR9oaArZ537h+wa191QH5fHSPDieoY3MDqkzpI6lrCboUNyBb/1iX
iodQLyW+BcVyUmCahfk3rYwPtdOj0qa+FKAfYVn1heWcZzDLIWYttz2+CY17A5y/0hdFSUKqj2o4
VmvSBbx4vZwYdtDGolDK0GoCyjX1bzcRwKWthD9d7kDTd8K+EZiBNR3L11r+t9l30TGFf3qfW7py
CaOcNbciO5fVAuY1dVmyek7+V0mowP+bI7BwL+LWyIKUxiLL5ft7MI1Ghved59hjfF49KP7rOYpw
mt5Kv1WYvn1MXgzIykWie4+8CBZXIpAzzCYnU/jurrGNqolPxcIQ0CVcBUAj0qy5bYc7ip1xF/1q
GhTMGKwJca8pDWVSyXWcfMFEsE+mUFDc9wJ7489KBpKvEmzzTeEjq+C1FF0FpaeCWfarqiixtZma
JUcR1a7gF/RdH8bjikOeJxpzyMR2HPw7tbhvUiQrSQcZfr/auGiST5cQA5MiPUM7zKQcLKb6Rqq9
VwSq1lpkCeGgROa9cEfs3QrLWqCabvFdi4ZaL8RZ8LRC8JFjuAH2UzmzqYzGP+V75vgyhhF9R5cQ
j/ZbAcxODd7eDAbaaWotWuHCwexp2n99Hm0ygr/8wHB1C9Bn5/3nde8/mlcddW6sPj4xIRFJE2JD
cNsmhiBnn/Gnoy6OhT1BIgDHMcAopKsZhEHUUW7wLFTbMOH3XekBPIZtDqGEFxrB5lhuQ8KWxHps
Kaw82YQQyMei+MA50Gjx1TIFoJqeawS8Tk2fY/0l+iwyXrd3XpJ5hJf+HKkLupiKkc4+7tROQtBX
BQS463F80RERThAmk5NmsuEEQTKOaxEF6mqRDUlvTfW8+sf1Iu068TfSlYFAwOhLFf5WRdmB4Lo/
izGAdxIqGmPbDZZ9JJeb0+3s8WNKGzfuR0JWwllyWtS3SOqfeNIe3fyKK6OmwZN06TXRUShV/L+u
vc7LFdMbutVoloJTObI5BcGCyZtDEIxaMBVs2R+p7yJq080HNHnSjVouoFDrI/KFn0plSf7TS9i5
+hEkrC+p85utcFXrvL5+H+ZAYbil7p2aB7p8DzrZReKncWGPSoLJMy7g4KssTLb+gvZTw8/PvEyI
nN7p3rmwxnSeMyDd1vIb8JQJQ+nhq9sR0TYLBzq8PyM/Hr6o41Tbn6A8PCRc5ofG4cdhxxcEr7hx
X08zaEFAyKmPlTOOuDa4NDNX/JVMqjKNP6SUjeUQTUTbXA8GADUTTvQjPf+AS44dlUmUj202bK0X
6nl+Y37jTA1vQqRE37Br6w70FZPVjGD25zoYE/EJRs+dWnmtnXJaoV7loER+qSCVYPS2GRJfgrVO
BfHL5wnTSKpkYl8UblZWzNKrhP62U/fz7ZG96ipyTehS8PDY5vp5CpSNsvzlWmpeEKxIZi3aE9Si
WlZ/8oGGC47+/5TXX2W31AufiyiqpEVP2l6dIk+Smb7A01bh1V/2ybvl413w98U4eQeKTE0tZqJF
oFnqAgxfyKoC7aihyz5fvo93WfbWljIaYh5G4farqN/f7BKjdQMRsvuMgam79JbE5nvH1SuniLnk
FvvpdJzSBidAUc/pX6OP0dB/llhEThgcvq4nHGd5mg2TQtRY0ukOYEIdvNBgb0cqcb3P1zyVuWSZ
MH3ArB92/FOs/q/fUig8TRPHNmz33QkFkogaoNrBu1Ns2lmcd6/7wnap5X8nmelKVNy6FXEEMqu6
/f0D0fKgK0u5enC9DH/9WSROzZLVV4I13VJ1i8UcaCZXmBk/RBKobCBLH/DpXOpf/bM76xI7QDIx
weNb1WnKP3w/zYVNGufJvrnSLFAJfRpjJ4Yu5LQ627dyUYndErdWDZn2sJj2rVpDyjnlRl/yDeoI
kyzgdbiVdZPo3rxUTkjqTFQzeLxfRAfNy7AB7EObEgSFZ9yaH4CEIYluIIrXcj54d5TdiBCLKrcP
gjwwS+USNKBry74wvFNn1VSXnkR/Lqg6BAx0WvFRCl027mDE9DrUuvEMRmuXnm1yKb8fuOpTrWtx
26RfafzkmF0/jx5qANAMngoiyecRgGQSjPW+mTLUF88NPaV3F2Ydm4Y7/obcoHChufYWgeFKgcPp
4tmbWsaO+nFAApHJXyiY9o+G5+go1kSJ8TQEcTWmLDm7J60S4nfl6L3jdZpGvNwixjNiruvuLbu+
/84UjdOOLxCpRsQQ8A52imHlaNe51INBxiR0xs2i1kTyNGtdJplm4Tq8zMz2ZapJKh8KR/XtB18k
4VBL+QI6pWjOvYno+2lJXBUyBRWvWTXLqXRxtk9o49XlRZ6vNu+MNaOSW4JUNlWcoKHY0UmSRuy3
FYFlvKxYmF8C9G178lTxqfuI6AscQwMZm+Jr5kizXOdUjSwrRcngTACTt8gjkJjmzhdp+vebuMIo
jX28YiasA4hfG42QNXTU/BO97WQE8tH7k54xdC+xErddHN9VrbZTSpR0Ui1AN8n5wABlF/XaxblV
n4YAKb+Bpmy3MuHS03v1emlER4AHjoC4c1IO+yPtWlpsc1MdqkqQmhlePCF1AAYhtGLT1LHd9Gvb
Kqd9G7FZngFz73Qf/d+7L3NflwMYeO2g2yEibSLoIVEaSVyXl/sLS4qSYh9IeFWqY8tg5ZXhk/p+
css7c3vNVDU15STJbpmYMDJYvsDsn6c63ygZOm1iNdOo8lmIXho9J5Tt99hAgT6J9tzw3kDVnuVJ
n+I28lm9yerG3BxdbQLhM0VwlC54QrBtjw1/L042T2O9qaBqpyONtWLiNGRRVSCr8PVAY08D+MCZ
sNf/TNP0chEPJl4IgNp1FIimNXmD+oruY+7ct8t/4Lu40e/h+P8uDu3W9dUoxHtk4uilfREAMdUm
eeF1MpNMPJBIvus1LS2f60UFgbv9fmVE6nyvHSB2oSH4DyImp/m5MncEINWR+94Y8Secy9vCiGxZ
aC4hdFiOtqWjJP/YNXhbjF5ELfrso+0n5DkbtiIZkTNR+4DiOQo1bcjro8zpcEfyQioybRHgQY/O
tBcay0Pjlx5+9oHTkIxNgl+3F+XPh9m0eceCYkZSBE5hnxav6cAGz/mF8/lTu+qa6KhL36CVJ+R3
6GYWvXVHV4KY9eue/jCgXi8jezVtGdRH/pYNLsXgXVMKCOraZ551WKCoCHv2eco40AZkpItOjIez
sNYwm6W2v7BldcOQb9fMjCmMOQVVvG/f4EvHWk/8soI93r6DFUe/kyoGXJgarOqn09/Olrioft0I
0vGk/WwyFRsqvWe0KkVbgwqt0hmEZBF8pWPT0wjZ0QxDqxak1UN/0Fm3Z2G5c0Oa6OhijALiNtg3
SbG1fAwqawlY+ymZXNWmPYeXLo0lDZoNty8+n3K3ngv409HV5HKtMOgGu7QJUO5/erd/EsWLVJ0q
AC64VlIKHuq08iKNcdRSBBjNivKoqQAUb1EzXWMB4CyKJWx4fuBz/ID2SRA3atj08xwxH4x5+oXM
s5cC9PKnCu6ElWnjhjwqZFIffypM86KrtBpr1QRvBdROdtuuItW+6oKhKzQ3xoofAMLnevRPYJ+Y
npJqoBT9D6+as5/4pNp7ZYdiGOaZ86ZyXSoCkp5Q70WpVIcNOsL94jSUTBRN9qsykTcjaH7ATqVd
Ik5Bylk3ebPEDzm82xGAlEVCbkfrHCKYoiNBMQkMqsY9wLqn+3HBNqKXHxpcRLeB142NnaeIcRVI
Za4H1i2n6YVH/oPKQDgbH2gLMZXtUCP7jDySLur9Ti07/Ix97BP8WQXHVB8CEWsdIPZ8S15qNuEn
NQTq4u1hCnYxGwug+SZTROZ17Qb4/cOzgJ/XWwP+OPd/1maNb0hLHcRG/JSmNNT+os3d+MuTnuio
R65Yko5cbLbwf/NUgg/X7oQP/X4b4/3Amh9A9wFrPBZbX8vWmKWbJVVm8SCsvQt3kJblWVi1pWHt
CaXP7LgVMgTG75DuCR3/WNizO7RWj8qHpI6fxKy4AaZCbTfvdJKYvBPaBr7pUos4IsGKL5z6bESQ
IzSdXWbcmTwbkHj3Zs0FF3QCtZ9dH4uKsTUmbBz1gz9+1uLK18qbuKpkFJ9ziXvARX1zepGUqVF+
jIY7tsPShqOuImKXtmppNJebzRltNIw6IP5N7X1W6wzPxIEv/1ajNSdi/bqMarII3r4pOmg3KOfN
pH94vgl/MuWkrM61Ct0PlM/gxnqirfkn0amx+rKY26UXfy2suhAGpgaacel+5KHEWXUchBAMHecV
lRI46V68JNPiyIVCuwrJzffo/t6Aqf8VfraP5pmSj1nRpM0q71j28xGWnx0LJ1Rs0nOINGTQesWn
2+m+RjI0AYbtXGhu30IlQP7epsJiLt/p+ZM6zuWFz1938IBCRuiQSoEIQi0nkaBR/6hjAwhfqY/0
d7eYuelNMUQtDadOi5VrWO2hWHIioQFbqd1myZUIRJHrKc35WfDN1yLH3XdxomuK4br6AOcE7eEi
G6NPtlpJr46ZHTf92Uy3ueJ9fltwSbmBstAokaNAg3D0XWDHxAjDsewfwUhqkyLEP3zlpUN0zk//
hUSKpKMksQU/q5l/76TiwoaO+d7UD6wK/+jdqDrk7ttmXMYL+4G2F5wiZW+K/ndUNp4V6/LMjgNl
sJQ4cw5itdZPhJkHO8qPbqWR18oTPKklDEWpnnJMOfMIo1XnkAGGdpQPwoSllyg8YK0IBA/pGGwA
OaAN8l29dYiy4b328XgKMjD9Bmib9PN4QyAyCvmIaiOiQIy5erzZG04o/exrVCYMifVHLv6EhvQM
I0Q8KUvgF+iaMeWhTVx0r3+DP6EJb5lAkpl20um3BE4LvJMjoM5JgDIq4g30mnPB3KXcjtwk7QXY
wM5ESqGH5J7gdwUPX8+s81VCYJ9AtIXIPsrE6llOlgoS7xr2ByxTHlbwh/Q4XFm5/UWii8MjD5t6
/TSXel8Un08Hv7INh5cEpEUwEj4H0tIgbRv53BrQUA9LAKy7LoxJfEdbnEjDTUrR3zHBeSI8qbLS
FiAIr6O0R0ahwyHPzwNyxlKSWeFoqjmomHpf3tLIsNtLpv7Tf2Atjo2hfTKW42GAwo3TNn8RHI4D
0uRWhIug1MTTs+iBojhnJXZYUWMuefQQSZWCjMsHkPMO0F/FI8Bx5Pgu5HVrmbIWiAxdt9ha9XG8
Prw1cvPDpz+eVi1hIfMIcDGYwuYLg+yCtmcnj9OJ4gEEM+ZxMdgrGK5Gt6OBWotYgkDcsNam/tU/
7gPUaov+G4H6NFwz/jN8R9PbbYFXqi0aP0YpMZrIr62u8u7CoIyn3/ZVOrcu4XvISdpArZoYowoJ
XT53f4XQyVWNNNRGWLjt/Bbp//Wz0KaxaPFU5LKEr4pc+ZuhZXGv15AF6M3VBgB0ELBdK6bxfphs
lqEXe1DVF6hJCKj5YWeZW/MaG3fOdL4TAfnO3FKxLj5q++vWo6r4vTu5dG09gG3SEb2Fme8fb/TM
KMSm4q1dv8OqEn3kYNEBW8lO0Ue4392NsyenqHn8nzxUXUH+xAhUWr5ReBDQNjcse2brctkfiD/p
XAVRT2CJkAVzZvUn2rQ5Re92IkOQQuGwXN95pN728f/UxOCkHja5UsyEPJf0X/pyxNe7OR0nQPpq
qniZ7C6R3v19we87FtVG14gx7841OKLJcLR5mW/lruNKRZjCXXOw+9FBDUMfiKbvGrdLQZC41R6y
AfWVaTOI+P+ye5kFmcoM80dQj6NwoC5fSi9uFYDHCOFhxMbUql0KfXpshW1Qej1iCi1uqji+tn7B
7bDRK9uI3W1Nmp6c41vSNLF6gMNYszDmSwt3/uZYgKtdj34/0BdQuL+pnT97ZRmlJREG+ZuoqPBk
PGSZFkQcqjZysfbz/lKdaBt6aAMs1Mho47Oj6ZpBFwKgR0jn9dZttnMnFhitaj+sMrGRKqeN3LAd
O0a6SRxFJY5rWFFKY0FBDLG7Dret5PYEFaHskEIKZWi0XT4cylKAWaWWoaVXkm1oVbWObMnv6dBF
7uiGNj6Y/I+h7LHJ+8lyfQhAKRitcMPyDvseeNqgNCVFP6VDPJHdRac6vAWFAH30IPbMEi2PtSbm
1dqLxgCn/lZ82Ft+rB1O5leNcczhKJ9JEMQH5jY+XSy6prRHBNPvaw8j+jwj7CGcYin9cSkGjzNZ
eUOEhKRoHMBRF1W8028P8c72sjOF3W+4XwvIFa/gwmUk+RKjHJHFWgJ4YXTQd9iFHEGSDZTFLW3a
rMSkeEDkm+QhXJhLlfdb2zufyYnnkwVKZiMNrZD8zTelH7tOHZAnha4rKPJv2kSMI2X4X84LDrPt
KlBiLtUWTsUUyTd4wvgypmKG+sn2KvBYQqIVRJzYm5QLCI4SzT7AY9YvDHpY6AEGZ6Dzq/1NgtJA
kEYUBnekKjqqVytUotStcsv/N4rWbnb8SW/T0WWkdWKyfS7nCDKylChSZAfKRMQXmtlctGS8dcxW
hs4eIO6qNKbh1FpvU5ES+Dlm8pAJH15MWY0KOEdXE4717T4CkuY7YF3IoyV+oRJn2PuDEpCHB1JG
JTLmH4+puT8QmVI8GyA6zvO22sOEE9O4YtTIjfKbm9q1KndpjBSxuqr9clhvgLVXHlW3uZVF8vzF
zzmYgCWZn67/K3KMYE+RzZGxiC0UHFqGO9OCYbK7ezfIrYXJkPx6/Yu/TUx3bBBWBcctVvooC/Xs
nBSP6GKExCWglHs0ilcykgsb0QKDQJPMnnTeyTbDzu5LmJaJW/7Bk/zS5C+gqTlf21A2Fd9Q6zOx
MxpmxP/obrSyqNH8/zIALTfzIma9d4a0e5VOpf2t0GsJ2USotxyLUDCmk1HlmibFa9pMCgS3/ul2
pkVGCgCeRQaFsbRuCQGEGHAEW9KzijWoBSIqikGNdvcanRAUY9qyzgtBM1nOEgWn5dLzPCrh9e73
V+F+YXuNGfmtY0AKhJYpOPQ8aUL7SqXr1Ad29NlnxZMEvKW3kWV547NB4rqxgvC8VMBVWY/Ocs5K
yUCEKhRTWy2u4LvtewvMBeuc552wVOSH4OapvgeEEDuSyBynZg6fmhejimYH0NUVE2P/rUw096Mt
5A4zG/qBDMWZaiM01U0YCdVyfvQVuf5ccmRFzu0zjv+7dRblorV3M2w4almAtgMIl11nG59i1UVU
TqpElSrIpRF16tpdj1TTzMyLTsD09mUzDjO/icBMcxOdvzSs9ydpl9KJsFbPRi+f8/xA1JTyMqhC
qf7xV1JnexEHCMe2oleQNk1OPpAyK67Lq7iLpR+VlHjoDPsP+hJPRgHkkP81F1IAl3lxwGJylSQx
hLzBLAl6fZdm/SRSkQwqP/uu1F16/UAXCCekElKUpFPpO5Kg/vzA/xZzF5tPcoVHIpJAZe+Mf20H
rF9z1W/KjmAgiCVK/iDBcLJskb3l/54rdQk84HM6aiNJy+hWIoC+rWwE/B3EJ8s+arwdDNtFuDbd
lyf8s/GCdVE9U0f+CVZD+p/DY8UAdg0sr/2AQNKynJdTdCaLeekwhsUWT7nlczkYwCkHy4rUVMJE
Mu7kieZCCVq388JPahgZYJXVIDc6uK1Zkm7EKKJZ7ed2Zi5yYg4Sj9OOO1g/9skc8zpuiTXcbTb9
6S9QTknPQKf/CimNIf+cL98prgM5+wjfc0V0gO9g0+7bp7bN2Ue6IWnq/V6GZzfck1qiObbM6FJh
5PIv04OS1ufo4ARoxVEkYSijZJDSnwMgEshPGME8VWbjhjzxu6GvmLuoqzvYZUqkihYIpXfLcENv
ovKDhwhKgt+1lFYBmLrUF97V/XmaRvWm1uCVT6uApfQyCj64HqPHF3oVgPTz/92NktQchTiuSdAG
klKBA5dsgxqrIFcg6x4iFRK+Q3lzXSfjzgmP440MqzhvR0nE8xdg9ltockEkf20w0IC/uQlKLWiT
UVjsa40mi19OkLpKlO9vG+I8KQIx0v5aYmw3oTk7QrUq08gwowpueUZVkqIbHto36Pjh/pYD0U+D
NODSY51T3vV92NumWjmrBNm4BaJHQkhNSik4HFmsHjmMd3FJh5qt88viQJn92hOSQJCA/8TrQ6dS
KoxXubjjuaq982qfJ0Q5Gdf4/YkcNqWh/AbO3EF7r8iasQUCY1Jq9KJIBVppxD5ooq2phymZTPYE
LThuOMhb9YOkPk4ESx7xWtk4LNjy8YPY6zJ0rAMrUDbWJ8LUPSicuIpNFL/NA0pARHzOkFX5oGVv
XXUnkR38Fs4dEeoc2a8Pu8wZytDuJEftCNC/be+akiZZuPB92L9NBprRWZNQtVQUpYsCiySJXDEW
59NxqJ/3lBGUxDIMUMHOfuaHHwJNe3hweWg5Dsi6Sd2fMEwoPatLKxRDntZvarroFlgyVrGnmQxh
ekIqQppVWrbNa0mDzb4uAWV6dEa3uK0jrWVD1D9PMPhhNmqg+vHnOHiZiT6D/w7KQA2c2ILhpKwE
bcSFwnbX2+Iu/KCMeIeCW0XcSuAW38VKAobhXoYquzCST7cKvspRqnHq4lM4zczU0XLviC5wChGi
hJ+JkI84/pqkMGFEnBj7/2z9Y2aPb9fL9B0yKd/E/k2n0vvblixGNUAIiXoqlu7H8eF7M4MZEEAP
o8b7AwsRagzRKw68NhjAQ93UtsFYGJ/dA+Dd3chm/wplUlzFf9JvxR0P8GXLNgxF9mSBodonj4ma
pjnpAHoOWd2RLSvPLjbB/MwZERgYiwTh6qZsW45dvPagDGPrwSL+t8+nX4hhs/RfyucuwPG75inQ
WFW0gwh+xtP+ZyJ1DTcDilnsy9ACi3h3XB+hyAsm2vHJN768ksu3CPaiRvnlWzcB34oUi53t6TRY
tGlsQHM17VHPIeUCOQxDLrkg1CsawF5ca3TKR2LBGAB3BaalpX++4F7MIkhrHvfJwDtKswDvVMc6
TgwrV8gcdJpnTfNYNo3jkPVJxa3cLrRsxCEGPRQja8KbMqo6vH9HPvOTlmjBgsucmD3P0xcE8e9S
VblhwrgT+1BfIpKdv7S8D3h0BnxiNrmkPqkQK9jXLBrcquPGbXcDHzWKJf+9j9QmvnElDSeBom33
av+0yjaD3nqrpqR2LnaGHi5hyhA+NFrmnaX8YxjIQqPmAL6zl3PZcOW/Xy9HfasSVk+PcM6wps/s
Va4pk9ogf7c/Ut233Xl+gqU3x2pX8HPcgEj4UCk9FnS+SslXMmrLhKckN2HykNKh/Mb6RLUy07Wi
Io1jNAyIB1mS/infv3/HdlSRcINYSrx7J9bi2A2NjEgdF+OWt8tiy/t9/B8beS+ZLGdY+8jjVBm7
WewWY1BUFU+RWib5teTaTKM6yCxMWo9o4k3KHJ+Lyv8v9WivGktbC8FieA+VG9ih+NQQsHerU/SH
fxiBrMVke+owdQM7Ll4ZbQh7Jf6dhNbs3/O0EU7HCbx45Uoja52qpEdqT4Z+LW96JFTYz/hJ0WZE
uA0SPFfexyOgepzaUDC2b5WmhluzVynxUtZhR/rpA1UqhRLQ9Jjv1LzO5PXGbc9C1xWAPs4+VkyB
pmlTGaCPp2z47WQOtXdbDZAzl1yd1g3YqAHBu58gE6MZ/iDP7cE7aftX1ulWGmbtILZ+sWvtT/OA
V6POvKyOKNDr004Bb+4v48X59qnLFm8eFzEMgTI62t4PFQisq1NAiO+8WaKoVYvT8hsQ1rFL1aEW
uzkESnNZv1QL4rcgI4A1aSoSBObTYrBQ4ukFhSDj32R+B1O0mc0fU+7EDwDXUvwNA9MVqPCvnpXm
2pEbSHVaC+jQs1uGzkvr1iRkJ4ueUin8RjERYic/dr6/7O7f1E6/21UJtMWUTdo5/8m4GzkGMmwz
lxsLfQsW+Qa7dHFRt418ZluqNHULT76ga12+swfA9QmM/c2JbPFykSugR+MlxT3PWLwIhk0IujP3
YVw3QS6sipICk1YYenjLq/yE95cWWJnzfpsJzOScgs9PrC5B/G1/rTUs0fRCRR8yobU2vbaKZjHl
1C3MBpgKswlBbY8mOA/YV98BgfNidf54mxtadlIAoSFqee1lwgD7RVjVSK3kaYj/9W6ynrGqD7ZZ
IYP9r7setCapI7/IRpgWx+V20DizHKr75WIEE7K4vRClHZ5kiK7rTRDuwDVDiDIv9cNNE+932m+w
n/v+UoErYNBK0s4whj5D4N/FNLFpq/Jo6iNA7F6EdHXpoAFe142xF4M1jY3r1b/McvTp9dcbGO90
XyGuuIovx9w4nvU4B1HscX7o+Qk68QHnBJZ1m54Bk0UDlojNAAnmG6oRxfta3w47gLCVtvLywf2c
votMHPFNtmg6HBErLbKvI3w6xEK27NuFi5h4YJYymy5jPjhsafIWr9LqusNLtK6eMfWmDoc0D6s7
h800dw2gg0mG/fN815khJp6VbCuaX4+fp9zxTHs9i8NGgs9oE+N2T0o5pBFL0CTHctbXb9sc3e+7
51WT6IEhnnTiUiOQOIhmskV770eMnQnrsumHfsYoUroD4nL/U09iz99vjpkA+Jgpl5eWxUeUmOqo
NE6fUjMRsQJq58BQR58Wj6ob5lQSRhbbJMMSg6z03qIT+pZiGEj1L+usH1EEf9mbp8CeUul1OlNa
bUUOBoaNRSzbxgHPkNv0tHm1rXa5CqO1iDRz8howcPozVEERl/swS4cHFxsv6rn3BL6I7l5DPYoi
4Tdf/jX/DHSV+67Q77GiPxpYylhzkWo6lluvbYjHzar571/itL0Gnn/Z2PGDuLs8oyhd1G2jNiqd
rK4aDh1U6aaJnYJZr65gbz6k2Eu7gyEKhkOa5ID3znKo7oT7EFsBy3aIcqjYQhIBs6+DEZ/twg7X
AiQlUNhbXhwYAwP7IxH4YN2FIgtc31XbB0F9Sei1Ja0T7CVCpRdNSGlFNkhktZKUL+veoEVY+n2d
AJ9t5QJeVUsrOiwcGdBUF+uW+RxtFdEU3fcRW8OKW2alETPHqcApnTeYfIpDEAGjc7yG5PqpGlwX
qqXu6K0VnTN4a7WuJ8HIHbWQ/eMGwpNevTtwYT8B/Kx69TdpXemX3oADKcSWQrpEEAfYjc+RruPK
CV9i5IE9VP4ZX7QHbsQltHegl4AA86t7dRicj6zXS6QKl5LbYm3Y0cmWJ2UP5HQKLr6iFctNXC9B
v7+SyYbGgIES30ksvT5Xzr5q+w7h1TV5yWiadrBxnvDVJUXKumyhFYCjZfR0geHKFI6OeyynS6m9
66Wpos/iIz2bDMMoItvBWYvbeptJyosSS0Rxmmtknf6L058sqN5h92/ifkk0FKvrHH5GhCr+qGou
Bo4YSXAnj8xi8OjR7hgAPVXz7qDUIpDQPX3s+CzBzFDg1kI9jZ/4OMQCfttliffubxQngUExBDvJ
GKSOw+LPy9gzO2//2BlptvnvAW57giGrfIu5NpbFiU8i7x4hEBCGpKOIDNTZ/fo/vf+/6sOubd9r
miePhTZ/2KOQX/DXwb3QFrCEGxaK1kan3zcHMsffAiq3C0r036HNDNQX9xSAtjvEVT5PDzdicz7Z
EO+LDCIIRK3uxJ9TBJYCb4rVzo4uGg3+Zk0GrKFzYOpwmbwK9pcKFhSK5CoHjSzkDVdpa+ouOKrx
4ArAgp9rAyrDm79Lgz7OZkfidddd/ryz98A2bYJmARzo3y8Zi2RFGSJlYPtaofabJx2rJdwrGAsr
iwMd7xitSxR3EoJq194kZJBPvwZFU+V62BlJ12ufWRzVp0IPwQy58Tp8eIhXI6CpDHz/6rrJG/ky
b4z2wUk653x++TiyW4Lyqt6HkLnDAxXuvN3P7YBSrp5F8Fp5pxwRLzxEFhvt/JkLDt7HlG8d5AmC
6bLY+cWmXVkaNSqdVih9woqY3/yrVHyicuILoN1AmgrtXodHVsPLyleHjblXtl4oijal+Ird85yg
Frsc4BZ48BgfWwEnHVKUnEXUEfaZdUJjhJloJPoBunXiT95njAFEwfBIfqXINaR0EEIwniRHYWwh
kj1LoUlzfAMRVL5D8o/RlhPda72yfhL2AlYK79hG/1UthtcM94vtmEU4Lbbbnc9nmXz9PGVCRAfx
bQIEtyhdjAGPd3qw7g9o3MzhGbX+Gm6O91qtSfAdmN5qU7IAt+47KVkZWErd/hn4Ebos6cKbGiDN
JJ20p+UquXTPHo7NhiZGSBSibVoGtvqbBxRohXU90RGEQGfbT3QT2zWokrc9OIfVzqLpYfZfgHab
alM8v5RuKlnWPQfaFG5XRTwL9TGexJwXOPdnCj2lUu/NHe83u4DoODl1u0oJWTidG6lDIe+FLNeK
Mt9n/0ghjsAM2sRct+svd7dSfqrcUcYlFjT3WwUz3osKg882lfEoqUpyBTikCmUzWlQwcARjxjWt
YN5SnhzEGRMlgdJVW2iaPhOjlvKeO1XsqI8MyaQJm91CmM7BLSUdq75YJT6qA6kmtRyHzYYt9YkA
7COeVuV1OWuwpPs7suwKQXMC4Czyc6pD/2PaYa0mSkXDhcM/2w17z7XZJIho1mpoDbAbZxbctVpD
SiUT24tXrZUk3FD0W6HFisZiSTzLW/BiO5pudMN+Qm20hAhIznXhyY/Rv2AR/I5/CxNlFq1YrHpp
rJQvb5rCmlqHh2KraUY+a33c+Fp8UE07ca1WQoBiLJ3gu8dfq1NEdsi+Tf+ksceSPSu7U1kZX+Mb
DaKOcP0Qg1BnNdmQF5QnDY3N/UkTIP+5V1m1RlE6IZ2XI18iMBjlTjPgMGxUTsHZ3nLFhuEGB6Ff
Mo6SCrjKYAvKsYIU+G7J/MeYu/cpnmS4mr/giqZPGyfQe5UpS4MlooF5EyxXUUXvuV5BbiYc5RZ2
YSiDQHlDMuLhMkxasFHmnOCBtbI7nSA556Qai0LB0nOOt9730kchncYzEwdU1+xgbKNciX7uNKbH
XxPN+y7IogQpL4jVJ0FOd3Iw0/88pjYSPKBjrml2P6Vh86bBf5lF8jwkfKC/KIuaFWDSmDZTw/vL
6gCjABNKJnD8IM0S9jc9zcJoN3x46vSF4eYU0jTfN26Y9XXgcGB3f8f+y6/ULuL0wspML6nvyZiN
sJzWNbpFOh7qDTei8HCqNzXBcEtf7zKlCmmxaNZB172LeRTkRnRkwm8zaqTv7pHACa7gA3Ol83aa
yn2fkB7RoT37ARR9W10TXogcdMPQ5o6IqcXWCCPyPed43ijkJBCzblcGyaonuy0re9HmRDSDCX2i
iimdY7MPxQKW90fkgs6WM9knbu4n2nUT7WN0Etgy3JWCk5Yjr1crS2Ua7w+yZzk/dA/QjydjIM5E
fRSABdeQCy1Rptshplgse2DJIL+aAlaaGlLukiFEXwoAvOLs1kqCcfWZAYWGc66wmyMgkf8vICqr
vrBhV0cOetwFL4xrMJZqTw5N6lXjyDzmU040HC4sGhu2k3tZOsURjfVMDXSzcLeW0BwvK2xwaFHp
7drMtpUVeR//JHcBp6xqo2zYl3AnBcu8fd8ZRYI6CnBE+6YCph7Tt8ezIM2vqfpoxLpe4vRoAHig
Xz/VV74eUvihXRJKzQaSAVXXZmgZJ6JVGERKe4g2umoOdzyIRrjmtKD2SU49Urn7yNvn700D3ZTj
al6ix1y/+eyq1iqqZNHabyLcjSlBkElYiCemq8pcpLeJoHTbUtWDQjz2rZEesOSo3D5gI/XOoUmo
A2wvL32zk6/OXt/bjJIhn2VLcPOVWPDqDgZbTiPUKmxVCb0TgV4jK4CnwcJi1QTfvQoThTHM0jyZ
EuqIGj6A6KM7D9oslZGKiTedm36mgcKh5T5qngCGW+6Rz+0pcud5A8yEge8F8OlUUIFiiKGm8hbg
XBxsUdAf/w3Bz3qnGzZNeNJ1QRx2n952FxbOxD7H/SzFCtEdruOyZjF9EqtkSS0sT5se0A79CM/B
0sEQVOKfDbHtE8B/OFq18aPi0AnzvG4DCpPUAi5DjNODONSnd7HDXHsaPGtkcnRSzI7Q5FKhFhLP
s1iPRNdp5/cujMnuPoseI5orvyvYMH5mIUVwfyyEMJOBwJzWXjV1viAhffADYmSvjYsFeAldcemp
WlHucnonSxhAhfdwvoMHrEZ1V/Tbhp/T7HCQMzGkWWzXTr/k3uWY4AjZ8JehRVo+tXlAbEa5YdzB
wap/iJ8bcLq4v7nNerrI85oSPrn13mO9X4PViC+L3GZaOSssQh3k0WRipG375MxalmJsImtGbsGf
wTCrt/vUH8xx7L+9Iunkum4kQzB2XnBNtofsDs+NqVMaNeetPsLp9zsPold2L9XaMexF9JsvGDuP
S5elzzHECcKatauR/sz0T2pq4BS88Ug4hHjbLgcOUY5liMbH2s0cj0am0AmyVWBrYdk/Ld3Gl0ZI
KEYJlc6aMIQSPeAgSKKiB+OB3ERsp6Ggzb4mWZrPwOH7DxvggLRWlYBFrqUeQuo2ewx/XV7Jjs6V
2ne14F8wsMx3/k2D8QXSZl5xRPwrR/LwZ0StFoj53vm302KNx6i85LOaAnMILxVmJogPedouhbcj
Wm8UiY560w2s3XOVTxTkZnT5Lk5XTCxrP0KmGPdz38jf1EAZn3WHTfbm7ZcegDUvhpZDxMTj9+1K
UPQyskIh9GlUrqGqCfKqR0P9ZRj7FV0/mIGBtvzGSaoRUpAAFGuTnRVFP2Y5JZyC2fPRkAZ563EB
vqKW3tzWHaQceCCxJhKocFTmLYibSmIr1iYRZ9Z4VuKJbzAn9KDpnCcaW1DentQPcRvptly+rr1U
FUErdVPo1VH6MpFh8F9ZG1O2cLOLwAlHLWwfeFPMaXkURWa5BNiYH32QjovCjNAJQd3IYSx/ACvF
effEMj6917mEWZ7qq/CLAMkJL3b+ArGll13sHA7Mc04ckuYnhyK8YTkZJF1ykYUy4Rj272FXz5Oj
zOpekuQKF8R9Y9ocro/KOezCb2JRW7RMsf5r13RC8N3uJuazOgqLC4YliFrduisf9w0BtmB7Wa+4
KVrVBwrbwm1JpKFhanF33iRJKT0Li3g6TiOb17QahifoIIULRgPbl5F7wYzJYHcabhtcxOnT2/H+
FaSTjpb0LFlej15cRu7TeDStSeztPnB3XXMe+HkbDZOht4tksCADCrXhAe99fwFKAUTXgSGraHHE
dK87MLv6PpTXYdm/sBG5FTuK6+76aRmY7bLW08KM5Lf+cXa/josKxLeIWVujH15U0dafG1n/t69X
eUeq6bmJchSd7BOA9GUyawt6/vFLZ8XGVMQJj65d30z2x0toNVpBYDDClT2c5e5csP9RCM1Cv3ia
2Y8j++L8nSVb+uh9e81c/Xpc1Xuy+rsZMiLevTMkIw6iFD1Sm0jKx9NToak9mC3tkj80JLALATHT
1+Hpw4LlktHKnOY72xkIYip6ZBeRDDLHSVij2hXY3qEK6qICx1L4w4bsfevhEcBQF1PQizUAY6KJ
u8qg4KG3sbLnV1c6YCkybhL7XyMqYeuCxskI2mtJG83rMNXN8k02exAE0Jukfcg71c6jaADFL5Tq
CUuQ9LxxtZXP4ke3cCYEFrUgykgkqVJoY95xgh6wEYCleMT6T30BAwq9FxK+YrvUmw2cuFCpnWHH
zAA8PrzWCFjmjt6FWmxGimS7GBrEDVlhYTYwFoVqSj2Fb+NL5DUHhePi/oL/amNdd+fL0V8k7CSn
WaUDdQBTg7fppge3Ai8cUXDbHOGLS4nGh4C+HV1NR9fmX+YR0a9JXN11wRFl5A5gwxakCfelC9sY
ZhBqgg9LoB95+8a4Vg3zNW3ecTzdkAp0KwX5qwJ33nzA6vseA5EJq19P+VKmIa8JJMj6uKs5vEww
mjYSknZFUpopNqR1I3xgOWvOsDlPYUwOgak/odI7AsG8YxpYYbhLF9qYQnknyBaqvqfPT4Wc8lXR
IouC+GA+V8VZykO11DwtozomN5bAbqv3tiUVHdsEwy7XB3lv4UAVfPXqFI7zC/Se8/8Ph35mNGcs
dbi4FMJKOySPInWsqEMZt+vkmBIGMtK49dn0tHofCF1OWJbbwwL0dx3xVnAX5Ma1d9+28Fap+ibk
iC33cYwqWdqwAveyyOzb2Nh6q8vP8rrEF71ej+3UDrAmF3seBnYRvypHcwPBQwa2YCUfFLo5aVG8
wrrDmcqBX802KIpNhr6RyDAPJpoFJ3HbnsYRKfyYax3g/qSP/uS8EZ7F1SBsiuplX54qD25rjPrC
BO/5kE9U6Ua1yT/NzRvf7LgQhxbxD2UWjA9hExDjRBrmxuj0XnZurMM8DANEkXT9sktAhGoBAgAP
rWhQZoJaxMji9KreFOncUy0DdE/HK5o2hjFrqnz67+aNq2SGAE7gHxWAuDGk4yUf6TqGfq+mOrXh
xqHyH7z3ho/1C0U2SrpJr4BV23jf1RGbse3t1UGSnhlvezWIQBMysZd9PeQtwmUWL7E5lMKwbfg8
04ri9eJKt46603SGDCYJSPMnDqvV3/yW/LA00QS18Lk1zD0mdMTCKMA8iqBFb1HH2wRyA2gDtuJG
DEoMRgyRjmfOyUccbWuHrwhPGPr+4I1/e39Q8FScMYtVBJHGrZODYtI7E8WIZ6llr1AmrS5qi2/7
I0q9AkrAESO2oDPJEa2CLUxHVoFyUfPIrMKHY4K3k2W4QSuVEmOZo1WYIep4/+Bh/SPN8Sqf9Hoz
LXfz7cVTLav/hJvU1a/lxEfjK4nVlCbeheVMT1hDWgnP2FklcL6ZNM1j4bRgnAuVAps1O+KZMGx/
WSXgluybxGR4uxv5RZgBmsIDKjEZiMPpIwu+TpSLfFs+CE9cWlYpXj6I7f0T6MYWMC4IdwHlQt56
of/t/hApm42nfYEY6AZgwWDfUqlWGrHin1OO6jI5/zc8OfplE1VxF07Eqs99MPET8tQrGBaFgrge
9QDhdAvWxq1BNWdjVk0Uz3QfV4mFNBxakR58tmLc/5WiQTI+ojNnHl73dJGPtVFXI+nqOWTnYvzW
y+aJ7W6awhR5ES+tsjntN8RBjELyTgQeoV0l7IIPWCOovxJObzm52Gn6YqyeXVlEClmSdbEg88q6
stqeLI1R+P4CjavKaH6gjkGL2Hy6fz1NY9+rJU1gsi5RJ0m2iVZBYvDTOTHdFfQb+XhRxsPpJ4SY
XQCFsOcDcDhYZkX0Pa9fP/uFmpgKtQqV9D/x5Wx4I5k0vqdUzM/UfH+JUc84YLtpTbebSu34ChFM
EfGUT8KC2v4hC+fEVuE1yfwFfKDBCMSonSJ3jVjUwWMmSOfUf3qOChdLygrz58PF5G7yp8ZfnddD
Zcop8x7FqJ39aiM1rOaQLPiFArElYQhLUCn861KDVbYQq2hxLQdwGbwlWl0/nwaIHcKU8gNX6gIo
oQ6Nh8+uK+TcPPHhjCzxhRNUDVVvhKjkDEnMFBt5+w8hbsgLtIXLAiuy6e+BhPGzkR3PnZSRgXb2
n2r5K454SBG+k3U+RPHrRyvtlnmPCI3Nikkne2Wu4af06fMlc0+RZHUGSIvJAaGzJGx/GifJ8+Hs
qBdf+KB9F2ugvLI4vuWZ6HWMvg3fn3KE+Q0EOeJREWXLWp6p8wGQV8zwEa+mGzafqjPSaSLdPQ8z
HXx3SybtQlD2pENTI8hmWOT7kYMrUzNxtaRDhQWtSWJVIXEi11DOyxwP7QIaiWEjxJ01yvrbv5Pj
ogZgdcwGkoNN8ptDAtjqr9mMCldpnbH+oYpraOklsAF2SCPs4ZZHhe1ks0wjpNbwiGXHv409ztqB
H4T0fsgZXANlTtpEGxdi3AvwzwWmVzp0SIzzBcMULDjF8cnEyMA/Qz1LFj13cBfu85wSwcQcfl+D
A5aSWZDvFNH4/wJhP1eLJg2IPj6/2KEn8O92llGHkEkODbHP0gDv4z1aeimwV4E3rmHRI7N3wziC
EET79/5HyPn0fd1fBGFkoMM+MDFIe8YJn4NaficqjpZ4M3zUoZQ5IBebURA+JWeFQhug41reAUlw
uaZTRwn7b0zB/I2mdz+lyDfpEPyO7YidFuCyYUXqoK6Jtk5a1/vxBkKsun7NEExHT/fN1qOyOeHk
IMjJwYra4g5RVdMYVuUVWGbulPKn11Wlj8WJN1LSbH51APrHDkg2IJomfjzy5gIj9fvDfRNZeAsV
a257Pziz9h4+HW8qgpqRnHlfHw3P5qHwy3RO0i/J6oo1slm91UDYTpr1y26YDjeEULx1fR14Rggr
AAQgnKFZ4WeTW5V/1qlBV2r8y9jclSSIeY4ul1OJ6BtE0cyqskUcFyMoNcXT2YhRYypDFI269Uxy
5kHT11h6cGd5vltSbBDNuCdLuBbK01xOoPSId5fEevtLVikZ+QO/3uImEsMWDksE5sfYVW69OipL
OAJ7FH8P5nkD3Dqedyqex/Nz/z708qC4fllTof+T26CF2DClJUCIvFiA5XerUWByCJOOLPIZQzdS
ApgdjFb3yRnxmDU70EGALC5iqhF65G+iXCDoarNuQH512uF67dIRCpoTBSLG2UKT3c6VEz/RSU5M
qT7Cc3FHhpxcNTYVk1Gh8ELcctAQH5lKxP90hRWB/luxjyf80Zwsa/eBE2ZjOCwvi1TkHs0yCCCu
gUvzPHN5GE0UwVpmvi+LX7yG1fC/fzvQZ9Bxn9mHuEmmiVlCEcztV1sTQU2oRZNe4o18E5VXiZpo
M/hSVhOWULKfL46U6oul5OBjccNKZansn8LMtJEdyxuMVLjVxgDdHJn41erm2o5N87Dni9qpe8qd
b9FMesI5UZzi57Uva9wvIR9crl5/eD0narnNlP/qYyuiDnNq515e4GIjEuIa5s0CiO2JWLAsIO+g
WVk7XPd/o4TCMwE9mInsQsCNc7VG/jo2q5+NIBAnYF6nnx/3zyYGupuMCfHa9dn8oKPBiZxkaRIW
hdP2KmnLMJgQWB1jLJhJ9bgHnhmBbTpaCWMecAkhTQsqyEz70wh4ormm0eQHNW6/DpisQj1WlERp
nQbiV++ghOC9nsH0ICwPA2hke5D0ta85Ea6JQfVtmC3iAfQlG/NwTp1G6lJ2XcUbPxxWiiB/dlQg
SBmODkkQ+gS2uN34nBbuRhgFLFDj0TPBTPYf9Z+RGge5S8W/YUkqXlw6u/xiLvIT2Trsqo3FI7Yi
bNUNR2XmPk2FeeMwAAFgEpLd447s7rkHhN2HlpF47usYb8aEe4NyTqEoc0Fos0O2jgD1PsX6ttnm
EfHOtZkn2r5etuz1ie5OrBTiuWSYoK9xrx/ihYq3ZzOyf300y9m3YnA42KwaQadwqeiVgBI2P0z4
/ZRi7A91ZNbpWxYWGGPAO/Aoa3jMNnR2eL8F+TnrAyBlxGLMQ6Wkh8zi1kMnofqI77Xh7GFKJ/hg
J4CdegMrr6y7LHIay/ll3YI8wcoIMvLRmjzD+4aR+gD8ZPqvJ2zPslgXAly/5dfdqjnGNvLbdtfT
/96yNgdHegF0wkkmwQCph1xziudOOSmCnxgI466Qd4q+V0xwBoo2N1M1QlJ6LJcVRn7+8nZR5tWR
ePnEdFU3NckhIwu7uCoYIqozfcsNuEXSVwwD7ULztngbdAfXgrD0jNrIrNmP/M4ICKoQkRI0tHvp
LR+QGYqtanzvqR8XEcrpSTCUqE1ZZYWlhaZNsPi6jLX4e/awWcB0QothT0DsktmiYAsjCheUK3UM
I0J3ISuTcibvjMPkH5QtT0sqY0XJM+r+qpD3+WH0Tv+p3JP4ga7IrsMbYc1cBy7XjDKSA4SaMvRi
pj1wu2XKrK1qiNqPYLPjRlfFp8NEvf0KRX+kV9HJcHYhm4rwfnMGoed6WiLepctVuMVwF1ceyux4
uHGv2cHpnmHwlzJH23DmPNG7nzSVbBN7hsAikOj9cpFyahmQTaLjKhNLlzH+27+rw6sGxg7j0iKU
ruc0t6OKzKYuU4OJLqQgmE/ewSRmxh3NCeUrG9mjLXLPH/mMhir/ZXF9sY9b34/CKwui14ILIKLt
gawHNC0Iro+p0Lzpg+f9dklPfbCDZZClIhcTwnvuO8JMCfILG3FJWTF715+DG7f2T9D/ToeHy6gD
9MVRe/ux/A+b4rkWEKktkNaNw2bLEMh6Ll1IwCeWBNtSgkbJj3Fb4WT6an8LSYaZz1RfYJjiOhRW
7X+kwTprew31lHcmd7XvxrOqg0RGSOxysTamPiDfhgrQdK6WR+6jjvfdWSPtF2PDhvAMix1Ijh7N
IhF/kAdZV4q9dkI2wN5mh9BGBhlfce+puSkweHEKOrIZ7ZgtRpy2NvrE0rzt78FmBc3ARiSkH3B0
iTxGQaTW9NHVmxwueFXg38zKY6FDGGZZ/sUMvDJMMGf3CiF2nrnIkX+XyZ6JrlslEwtpWVCkwJvs
raGD8/kam4jjBJCg+cBtl0d0SqYwWiMoJfglOUUvAIa2k6t7o/UfTTxLY5bgyMHTpvDiasV6QRWr
7Zldpyx0ECUj+fyBZluhDUS1nTR42qKlZAMGMZMNFnZx3tzgefQ6DkhKqxAqqd8VD4obZ3bWUG7h
pFnURg0mdm4DGPv2Vz7dp3+6QFASU+M6hXCAHjr4MgQ8DNG9xPHJsTpqmJWnqb0BemlH/jgkZTJO
L6Fni9KbxoVBS9zCzHMbrlqUo5v12lhw9fJ2T99H2Kv62aTpLCEETM/1r347xQnF3Tkn/NVMjLwg
/Po+ku0iOAwF6TkXIhi4wDVwT5qMqKw02SKxYplnK3YofIeNAgJ+FbyRvJN8Qf7aq1d2RAKolk68
D9wlgbCzv8cCrNBuK6emkyZ9bdTkTNQdRaBfhKy4LSdZ5Pt2MZEBBcKI7G8GMEXPNdaoUozN2IYu
B0KCRt1M3ikPuJtjNv0hRPC4JsVecMJUsbSYvHBqvGaCqHZEspmhvT3wgmDWsA0ah7Do1tCi1ZAq
gkClgvlRijCX7xTllGym19WE9KsaWEmK0+UqcRrut+pcDwg2LbXgsQ2lmdk9AwT7kptzCfZg3rsR
GaRnEowD8/vlDoZuaRqqLBwvIdm5lOQ1nV80LGBZRk0xycDUJNHziFWHXIu7PsfibGkmyuYqAdlP
QkFR9GMvQjWshiWja4r2PuiSsRpt3THgRKwVD1N+JT8arwuTjdfNCeVOL67QceWmUYInOC++8di9
TKb/sqcI48Mjs+QZiRNIc7XIyhLNqNNVvFOFH3394NBCkdtNIe4rwK8n8JchgfQuYsldxwh+j6uj
5l0KWD47WcCufjgWuR/R48QtF2Hj0zXDqE94XJyz4ZGH0LdXnJOZO8jeOOqpFKceMvzXG2i8FFjC
xt40PXr3qcBNVNJH62ScTUofgrQSNwWi4+hKATUiDVYjE2ryoigWg5px9l4sz1cei175hDRbp6hH
vqEKuIO5uMfshrwUUHlLk6zCXN0cHAFmgU5MLgY+uyxguxb1d7ZQo9le2qgyQTEz5hDjjIbNjdog
omZQwmsNQHjOuw+7+lQyrvBnJ1EwZA4g8A+QQZqPzZW/u/U6aC3bt/AVtE6Wq34poy2sdhzYdQB8
FHKyGR+aY8V4FaLARqIzsGz9egDfi2IMyg7TNA0fU5u7s+gki2InBt6ZVAtcdfscRc1P+62zGKqy
9J41AKXcHmnSgZdf4ZcSgstEhSV6cJoAH5qH8OpS/+KGxqTXGhUGts349RBNUs9NInfI+HcauuO0
4uL9hQ8tb4vF8AwfkEu5uFiunwUmTva4TFK0e/jtcEHAHoXI1LV5cLU8d6sUDkC/qm7OdGT/V6DU
U46y9XMBx4PVztxz5oacSGbKmXCCAEMhsqq18yPY3gvuHWhFCMg5zfyyFgW/+p/FqEsCkgeJVfdK
BW+G9RLxWP6N5r1V0yMjWrP3xkjwpXXdXxouwC9biTlUOLGbLz8NTP0sdm/G0IIswurJFpHpC7/Y
XXe96B1Gfc4TsWpyTC/56DDTt7pjv5ilTsJcckMRRIkLjFBF+NWkE7rNwkGWaOcCTvVl/+5rc3Bo
U5wC2NPfxuET8Fh4LkZrM7CrAdYKzWBYJskENkqaKlCW+n3itoFy48II7YSe0l0Q32udU2M+uf5m
MtVaAuCwOv1jjmI6wwxFHdqGxyZDIYZl2AIY9lTMB9rFHantangDfx33gY2Ocjr4RcS6y39QTTsF
cPjzYYVKta1cfHMchcDYhxQ1+591vdE0aVyRASgJAjTbvm1WT4Ksf9TEpG9yD/29HecvOuL5jBur
KIcu28K7lk9laSeKKmuSgPH94JDGX4LDC9uOF0lnSYu3kFOaU+IjB8TDi1AyuVsAmRdKs3aKpK87
OwnZ6McYusGpdMVLpUbsXH8CZmyWP0QYTUi45fPW3gNwCDBiB4U+qq1kQ3DATEJNhANOYYXOwHOm
gXaV1sUFhgRFWZH/zq9I4UFY/0WylgOmPXFoKmhXc/3eNHTCDQ8yHwURGu6m6TDWEcb/KVaa6tn8
Goqo0nYYcQiRGwwQ9Q6MaZyhviWKyVkMe8idkXtAHVV4ZKxKsUJbbyCTd2l8V8o6IBL8mLNUlQau
lsCPKRS3t0a0Xb13zO2TUwZkF8GiefsVLqqcFFXjuqRW+hllBSfIOVH/8NgnT9GJqowAn58rTAd+
AGhCQ0SLQPXvyYtJsz4PBi0CtJvBKGBYdTXv+EM/zQSHsXlMbncaFhT7Imy5djBFhp1jl5k1EL8S
soBvLvJutFtN7g83SWIqLgE+JHnn/lxbgZBsIPVLCBv4aZEW/ox2H52O25zFqZCDk5h6btqd6cVM
YEjibYBJsid0l99kKm3vljzmmUzkSjbK0sxBG7BhKur3RukTSZj0qmrNY3BflUNwenvnDrYYV5OH
HQyXual7e6MoBc+xRuUxKNeNocAyazWPEjVT6hYfy+hE2lY4Rbj2A9ttQBhii8y0YnQKIV4PSLIt
zWLLW0cTaDPOh3S8ZeXxQZcxmMA+9GN2/ifl9KIaTjXb9oPxVTc002Xg842aR8acypM5ws0yrm5M
9+cIAelal3y/5tpDVNGjxsskJ++UpyvXBHlAVxQSzCLnlmdjsn4AOgDoCdF6AILQw+NRRMPCv0Um
WgE8pGVnOT4bFGeqxxc/4vQoFRDcmBdmygaHe7yn4D67U+SesBy37XkkK23LTPb29Xl9IqU9FBxZ
OCp3azaD+GYAEOEjlm83bizQtQJwEYbNL9Hq3YOjV4dUklnsyB+h1OxkxhNCX3QyuYeEdZFfZJcX
wEqzHRLqqURphq0MEDxl9tr1ZFODPgiceTUEiP8qyi0rJv0e162eSV7T9EJLRe0mdGnbTK/GC2MP
kmkLSc3eLpJjyMAg2D9mcUIsKPMEgFJ/bthDv95BGr4JGSoPZxJisAaA7dWjVc77T/UYfeFGUjOX
u0K6SBcOQ7QDQCwypiH2j7tgsFnm0wqdDRpobTor3Nx33C76/lgOP8rVzWS+WdaajIcurzSg17Nq
l2beGfK9JoalXnYDL2fUBRwzR302C0//EEz7QSHvCkI9x0kcpnQtunfEgKH0V3MoG9VaiOmo7DVe
EBzSd1NsQLmUIEjXKY43tnzzpcsExFZwQWH08fbZ8u6TaA6KZ/L7LBXBiKzLub07viB7AMJPxTAF
RHTuLPvgJCryA1dSggyjGx9huOnv4tI1aPY97bNsZBBeDfUshnekJYCV2uDJ79waS9QhXd8BeiUz
GYRUN5CpF2Op/4Td8LzVD3SYilyMAO+ghjt0jfBsnoYXpYXXN5OvGYCIhvL+Y2o4nfQqYRrqPYsr
5eVWEgiw3AXIfMyJp+ddzqwbFED1teXdD31yV2/poGwRZKqeoWfvR9blx8n0si1+aur12iqJ/P6U
efKMHttQ75smqgkwH2e6PngsjoCcyp4VjXhB4/5GFlEs00/KHPbIBn6WgrzH0b8YiRjYut5NUeYx
HHzVjXtV2hODubgQ2ml0MTeuP+sXZmF5rw4UlNPUS5u2RiGssVX7x9JyMJnWHxac1yCaCEhp5moM
HTLl7REfth8+037QdQSSTXOa6qF096YbqkwpoXfLgDwxECabg2XqhwHqp3c+G3A71pP7kf+MEe0o
bTUj9hmbJXCCj+bsSw91O6BO9nIpMnounJ7zyVtrrfewoPmS0i+6onz/pMz54r8kAwyJWWCKF6l/
XFQegdZba+PrMMlQoUQsOBbH1s7ufGOrtOpPtcfOIIZXhXI6IGnLBeGL2TZcJAMjS9J6NBXPehR3
QEr7ouAq71ru+z6GfFJ/K6rJdRrg9ZLMX/oPBWFSDQ30WdKvv0GbGNyMXMjDGAHk2rTrppHRpmVb
JgQbLrl3eHjnYn0xNknbhU7MxMi9EtyIqjQwETcXCKPt/hRXvYDyg+Vxjn+kEKh2mR9cKj1C39kR
+IEfk5v65e03UVoeYea1jrog5gBMlmErvtiEPlbjLxnhINF+Qs69DF/v+iZmClFOONVtnvAUT6uR
F0HKP1Uoeuo9AZqa0KFh6AxLbJc8IFfVA2pws5yKmlLp3y5cs1OEyC35ANlK0daGfrgkGG6oMA8o
hX2X1yA4avL0u/U9kn9SUb5x0zD4z9THKu+uyjtugyS3Zx4t9/KL/rOhgDIVtoLZo7gvnwrrv1hm
m2U9X/yt5qJQnvumkyaCFv34uwe036EQeAZKBza3i0vYhrHxjRr9/Dfxc9Z7Z1v4rwWTYxHoKt3V
47z5v3FzbigU7xp/sScOMVz0HINm9NeEC3c3wNhESrjTkSWXF2qigxQRY0ii6qDFW0IBxHGzyQYo
M7vrphAD83wDef6ZWfMaZkTF23c8b8GBh6Giz44bLtCekZhwqUw6Zm3FO4StwuEW5lJeSGkcNzPv
D9n+tGJA+0v7eLp5dlfv1MJRCkeBHDjmZkbUtzVeYE5dNmHpGnwcMHHoPlsopYEIfd9Lbc1+f/qe
a1FNYbz3s62n8X9+B+gMh2eJN7VRfLBzrMry4UQ6Osv1vzLKSLaQq9/uaiRhxzCRv6Dvc98nTrh5
t/r8oHOinEi5sJAHGS18M6s0PhvORQt+PXny7GS+zoEfbCo4qqRPdQXUr5/uQcwa0w5A5co1MzHp
8f4pgyAwCkCUDWjeAGRz42y23g2+KXO45uvB2qy+fHsd0NJ9GnhYetRToHun04JM+sh0N36ss1od
UdOZG2yNAM9H5Zj8vcU95pxJ5sE/Fb4wOCapUBCa0a7n1NTSO9Oa939LkOPK1LfxtlpNRBjm3wUe
/CgvbRNfpOwZB/cn4X9Vwg3d4M+1MXscxyw8RtxmhLJ2XxbpmHO40GKRtTYacaA2zHQO3keat6v6
hoGsZOhuITTvYwi5O+uD6PLNaSMvch8oNst7e1Sc+RxJoL1csn1EtR2nWZWLFPciibcP+G5HjL6l
JMGJyStLJAVxPCmCSzMe7MmqIe+IYg3oFtxciA/p6040+W9TftGL4ybpeoV1iF75kIv5snXPyxIQ
vIHBZWQRvhJHKWFWKOETYpNpPJmw4iUTxZ/T7zwZOwTJVkfqWF/b1bdkC5N25BdlpujpPlt9+tsf
faf1MR0qfd6RkN8uz7A60wVyUfCZlbzZpNAfrraHjdaqNx0L0jW6zg8xvsb1X13fGpMWYHrESYG9
yvkri0XixJbfzWUaod7UKY7NZ1zFTV0DAGo15VMi5smj8+d0RqPt6LtZS8TEHlUbIpkxV6RxXDKi
JZ78VXq0HfAztM8Cnm/M4F6tlZG9VdYRGo6HVQAYtxjaEvKTqO8EJAwpFIS3IsfJq1ABcO5L76/Y
3t2bnRQp+sB9AcmK1uZY4NjLPtGNrHAVYf2gtCSHoO3q9Mwl9hooNFyEm8miudQiJF/Bfd32T+ES
0IdFM9j9GU73XJkrQmQNHKQDeENxnqF9uuHv0EewZmZ5GpDIX88HYbVCM4aCR0P0E9Vb0g8sfcaF
DIvgaPL0XHl60hbmSPWFHMFNAdtuhQdEfIWEdZTjRl6ZBd2n9qZEjvvtBThxWwXzQYwf6w8Ol/wg
s1izh3sk3QOh3qBCWlMej5GeabvyoLXIy7YxmfUsOlpHoawau1ytYrKg1feMfzfLXusLYgEt499z
vTRaswSCqObCeK7d9vDMoC1U7+zKYWUfn70ihfnq9oSX6AtvpfH85lsCBvv2F1Kydu9j5iLwCRYZ
9mAx2z5rOJXSTX1yVmRLWt1kFxFR0vPcxVj+YZk3U6ijdzyRzzzBUCBR7yzLIxBzIQLcAn1VPmmf
mOQEDi0k7pKX+BwhD4hE2D6jw0EDQmZUKnRWtUk/Mx1MTSNYm+FRrFJE0G3WJM1rmdXp5O2Y+sFt
Dg+jSrwhYWY4AKUN1sTnTYMH8WctwNmAokQUqOE2rROzpVgY6sBHX/DUFbI1FO2p2sTh8+znh+xX
i8Y4v8hj3gkT8FiXP9eUriTlM6kcbIVPvGiMdLzqDvlNlyDnx0M6eZlpLTYQX9OjxL0k8Zzq2Rvw
D6CkHGJMisQXkM52fnLntUHrANj7POcWVew+gq4a1b9AuSHIWstXWFnCTW06HbW1h+EyAPTr6uAw
WIfMy2R0KLnvL9qjg0j192meWxEdMKtyvaOfHuyZHjXQOINwkG1Q8cpSnlpa5PozkgKvYVZe9UDH
VCsNWOhyIlmB5xixJN9JKZsZwV+PnVsZXYxQ2DWMTme6B/T+vhDayGtNHR4OjreWVI8i1JvTWTMM
7Iq3ToeuUaXhoWAPzr8QagQN0UT4howYC4CY4svALokpUDPkqoFUkee7MCsu2pZZGxW+KwVMOFWy
EZfgTqmc1rbHyG9GOICBuASrfhSc1afLGdp/fRfy3PJjgBU2Dk/Vmjy6i9ybgtwD4R7yEBsq62zp
NWqFCnDCnlqvxNY+21LuERYFT0k3ovWKi1uRuDwe1yPS2siI7vNDTSbZziHtLC71j0K5TOLW/Ez/
hguDnQ0kdgUV0FXQk4Tbv35qXrhDfXb0u1wTxxeVcS/7WrcM+k39TcBKrOZ2IrDVNiIXrPBq2aeh
V4AkoAyz1fgg1Z4DGxObHs37dpCypMzR0/cGv+mrdm+EEihe0UeJC0wS644xspTcqfbIoug84DI+
Ep14HB3piY4Lgp5EUwbRTe9tqvwyEfDER7O+3AYeBt9DfMtVhCU3yTsCUk7mh3JsqbI7ZE/XR2dZ
R0XQ5/HZd4ca0r8KsNza8CoYoIwKnEpfKR/rPv+xbrkL2H2baEkmM74Dny6fQXZ9y14pF86y85Z7
K/bn4980oySkvuDkn/s97inyH2g5ibULA1GtZBpYTUQRasnUytNUu0bU3utaXTWTYZySs+mvYPPN
A8z+Pb8JmVCeHRx082Q4m6DPxJhThvxqBlQLBQT3V7kkrvofny1HhPFTKbz5NEzsp5LaCwmjpsFr
RnUrdLFyAgE7aDWHd42Nii1mUcBJnBTEQ0+eIo6mFnGuWuFnllUz8x+jTCoKvVv/h+4rTfv6y8Zh
9pg/zzhEG0g+XYG5s2u1Rc+MdyxfQe2ln8rJr6XJt86sQd2NA6SzCygtUft3h9bw9lHd+0MgqfZG
K+d0fm6w+6Q4KQnnh1lTBOiZvLaDOJ+twFYpLtscu+AJJMPUOq3PYI1kvv0g8ak/CDSv4aDKqgwC
AsG+JiZHVj6ayCtFkY2NSQqADVksjLNhhPnKw7X4UCTBDAfo1qXTUt53VnwVTFjpCHBzcMtEeC2o
tGRiO29cnYchLvxURiwmJcCtVSYP1sgR7o1t0XBLPU1Zx9heyN0iswMJxoq9f/0KWGfWhJAoBIKt
9gN2qo21upWfZ3iEudm15gVlkiWk3NfOY/9OLO7TMQxwx5t0ADvwQUgz+KeeCumKXQAjDN7ONRSM
MlixTS1gP0px2HFCaNEfk49NejU1JSdh2DcJvZk7YwW4z6GFHVAXneCTlf23jhaI0aTBcMNBuOnQ
8EdjVR6cLJUhr7dtAcLZ0y1ypBynbgf11dGEUu0YAQWSwepezlVOlB34v8ckAyk6UZqKpHgAeGwJ
efBhIEDCs9oAk6ma39twyyH5BrCB9YeiPWLzMWGaKBMycKPfVMoz4Rbe3fjwsW+ik+6Rgp98871E
RSmSGI0U/TvdeACmYimHEgtSzWEZgO0Ib9TtanZgAXV/6XA1N0wJ++m4Xhvh2hmKI/JPhZcH4RxH
nymVvTFvWhZ3G8B/Gqcv3zlgyqu/m/b26U3A5qHihepepumafZSmIfIBz39PS0q6I8hVRasEUKrH
LoRNyumLW75kUiRnjfR7m7kgCAgmsYC+DxOrrymZQmZdbL/ervDKHnkvhBvzVyKJ9cUvKb74N7L+
auJzv00WPryDTXWda1L6S2j1m3FjcNwfI+vHBNislD2wgh8FkPSFwMYCca2TPewJTytpfj1w7OOG
IR0ZJ4IUwt/W/+DEhSdZKXI6YB2mYMgOiqjTc4VvgMtBMhGFwJ8hOXDDCKvLp6EPSMHiDpiD+5vQ
u26EjDJDxZD1ofaY69WUgcah9XAB3j/rhD5nK9E6p66kFVt4Ql4EOjldZjLtjuSjSWCfnS/jBYqr
SyZYOWx82tnRdlJCTPpLiNKlhhH00cMbTBPWfzndbkHFZ0gs2nUa1/Ma4G8B9sm45K618Udvikkh
IH3weHyboWS+qU5AcuY3OV4F/Ac1gkOBqrKCnWewAuvXAx+qn2EngrHvdQZKT3FTIbZFDokI8EPJ
Bt7SY6ZW3wfzGn/CjNIzrdbm1PCvw/xm2HGUeAuC4edP6LJOCvtGJdH1Q4OQOCQnJ/RJfyUSPSDF
vHNLwVaRZXh0/G7gET0sLREMZKAOPUuGP8W6imXjVeNMmo2IrMA/7lHN1bAFVspTQnkBXwyJwpJ8
SPByW77zGDlll3ozEdQ6HdDDUmg0E+y5lvQZbU7LCajJ2drTdn7eYMqtskBlw8vx5thEf/OpjN4U
eeeDMn59mJxRRkhLlrguoDW9qzMTaYbqzh8aTiZ1SZweT5suO2P0goUS/Dbv2cjbVtFNkiqE0fNE
LfEcqeojHjEzokgsibNPr954W4XjqF4G4h37zEjwnds3G0Eufd4P+HvqUfnEXcZe6kdl+G6iITJX
beOCObAS00UIgoclMPEs0SdMeHtkgcjcULBYi8uEtD66+0ocuDV5/PA5pwh0VsPSsud8QHRFbdyw
EoTerbZdW7Z0ucX2wn+Y9eM/QJS3bKqp0p7FVDN8a5Y+wNHS5xZ8yeukW6fKQk5opvGhDlkc59dV
qcMOUOiVV9apbe3ZRyJIlQavf3656Gcuo5KDZ1SRAhNUGqvnvE7+bAWULzOQaqec47Zx4rnyum2V
WKQSW90uVSa42GDvtzBOR1yeWz/C69OC1mMwFzyLtjwdk7JrONkqaP9soivGPwqqpD9l1gvLTHSz
RmeWcpzycA+mPZK8N21PK50HyypYy1Qrd82Ru0ytyocuhJadFsd7JW+vhPHwy9L1KmObmxWYr08X
oUMTM9AljH+m1v61e7eOsNrJZPViR4YWGceH3oIMt7+WsRHm6kPVBocQP3rewW+dHi9LcQAyiIq7
o8fxstI2uNZlLUDaMO882h2rQiU5tEOsbZlCyAeMUF2gkTpEZ1joQtQG3aK/ws1dgvgbq8aeEDz2
8Sm61eZgr3vwhd/SidMlLmTzPaXmEOlCrJAlT17tqRLxdJT9tHI5Fr7lcGCOGChoMrcj6uEN1Zc3
0XCdV+vMQhwYQfjVkqugN+UYJhPsx4cTCTXQk8wQp4x8D6Jt+v30iViCA0lrUvKGP6EBrdlm8aNa
U+85jeWNFNz1KbAip8tvdtiGwcMn8Cm3T0kgUwQlqkBmJpkgj2DX2uIqJiIVNs5l2afk7i0jf8pJ
P0B4kmEHQdjgTML45Xxvrn3ERl5aTSRKiw+tQopxhxn3g3SUYdLrdnTTrkBeVmYOx6k1jOz8UB2Y
SPro3lNBrZoIvYqv+NOjKGDyLL7qLgsfXQzL4OfDhLbl81yjpw4SSjKo9wQBwAqQnvFGIqTbpAsf
CogpgYeWLWXgOqyTeShzqUOX4NVklckURWoPuomINlgsDlQCGmTA+OeCdm97DNOy7Ug/GrfxRzJ6
8onOkmSi1IBMDgJ0WR8YPCe1bKDwROhuarlRrNYjPcgiQNjBhNZTvguRXPOOiIInhaka1IxtW307
4zm6uUiMalWIHguEvnh2rAxb22ULZetHe6hHDgIQ9HI35hiq71y+NE2bu0HmdpHpAihHq+bH5LdV
qKiUPCf+FJaePFIiiRPfrDNv59QL9UDuBdpany2IsJ8gJecrc0tlXXZ4CoA3Bf4XUx84Mw0Qj6zd
G0lQNiMiixv8EgL+JpZdG56D2l0IkHJipUlvyR5+txyDgUCmj1Tx01td5YusYwyxaxEt67Dc02Kh
GZHRRzUX9xRc4v5UriAxjYm6+Yt4kOlLAQSQTTkSotGeN7qLpxfqOf7GdgNYCF5XcAFLRdfD+ynq
qI4vZONRP3+4muP1M8WcfX9fGgCbx3Nza/Ou53EOT2q3Q76QEBYvlX61GPrYmL5YMP3UtZITqutQ
pkoJT1yzsx5cYav07cr/aYBv8JdtvIX84ifWDmrqERzluOBcE14SKI2qT3oOdEjO6PJ+fsflptIv
01AaDSoUySgOjjYVOTOGJabCJPDwoZCCvZZZ6cbsrW5xnOgInUvgIr+jK3YBwb6PfWrlAqdFSSj5
a1VhAYIoluQUMkNJJRqFqry0H9es80UebBu3SZDm0ZkOJrfmT6OvrzqN+BwkXtegBUWtECy3LZ1Q
bHrpO0NML+qHcExVyM7w54iPSjsGZrS9RL4SOfJsGwjyn2duclZu/a7+GqP2PxbWBqmYLMUwLIyE
Qk+YG8duv4dgRvWKAsDlZv8P+4LL3zFLTpVrRJWVckwymXLWke3+RYLbuv+q1H2ihoRKka3QD7/H
955PMkND9iAh/vpn2Bg5TkXyCFOiqFWEZP8vtl1k6aLxtGGxyC7mMagQPpX68/scTcRowPm68Zay
rVdKjV/X+gBmPSRDTIsZnVaqysQMC8s1Be3UJVzL59DfbXi6msnrYbQBPtGG7SwpTQ3869i4bf+G
O7hGPAc+ghz/25l1ntNIuvlK2lMDDfC+m5tAm7LMrvd8k6MaWku8fQVuRp6mrvXCWt/ALZ/pO2Bl
NVmHSkOvaL3uSqdQH1wHdnt3+6vvLE3St1WaSOuGHJEn1FOrdsyexHOfY/s/n6wD026b0zay9vz3
gF/PGWQ7bjPPZDCN4by/ckWQPGWGSFRVBN4BWKAVVuw6RDtFVFi0C9zpPtq8z9TOj4NwMJKJCsIS
Aut6Rn9dhJXxl8t7RLqJq0LqRnX0biHoc6d71ovwAJ2UMINlArboafwKIWGHgFahrnSfyInRH1Ie
bT4BZ4vqDjPWi+xRqBXzQc2k/pXU8qRJPS8rkFy5CXwgCYeRe+oLqjZ7b3+uCgvfZdz8hnohg5t3
D11fQw6FrlNinrbDPfHzMcGE/Nt7K8rV44Ew2WjFWgoP2c/DLvUeYDwqu7TsoezTuutMLXFapxFw
1Q4X33MZ+1XeFyw/yDJQ9S43R2qJE9RAmjEVZnbhMOF6ZMO75fvxWaL2fEy1FnhpZ5zqQ8qa/2w8
rf1kZfKBm12b7t2zcsYwaQ+8Qgb98TNrFCaGLyDtVxQP/kUNUBn4OzSmEqXBA3MeqZocZux4y7Tc
8QLsNF250HpaDOFlLQVa/9JB0D3AE33/qh46XREcmg9cR2gKYhnPkOm0jMzgu4JeamhjwsjK7L8/
bGaJ9VHwYeCkCyK0tqxG1lOVwYMC5lPLZGr2yyeWSDsjWX7WCGnATaWAJs4EfHPJ1HDmcvzagVkl
GypK7u83OOSX6DyFneurlrergA6y93XdhIRwLjCCmyIkQhtktgIsTWNDM7EoIAWAE/SEv0e9jnxT
IMzrOBetxVJDqRPHJcPpOl3tTiZm/P7c3d4o16/8Bphn5fxRwPZ1SdTBjMf1u1hpadxryh0eLSKy
gM4FL3ciGlBlbzFfwt91CW8K9eak7Ue0mvORXHQSQfwgVO1ERRlGn1BoRTLHy28Gj7qdd00vDSNm
9q8MHn3vfyhjAcC1jImb8Mtd3RBJ6goFTUCT+O3pT3ZwIImKrzw0q9Rh92Geqr/nEk1W1/1eoS7L
tyZuP/KWsKHbd+eRHKRtkk4Ovo3khHz0eN9Si2pGS7UZuHl/ebnVXmNVGRFGMVENa/o8wRy7vR85
v31O4qVpcFD0CF+edA+uBaLLApdf7deNSD/qtoklcOKWDdDXPXC19QHBa6gg09n1jpaeiIOSBkhH
NIjTGncQvnxO1gicnHvxYLrpWHskA4qMFYp4ceG9KhuF7plWaBChNpxxql34IBZVWxa484BnWKbK
FEwhxkSb0VKW2P4q2QtFCGFH/4+IEL6cXRW8BeAofFEv9csfzCB7YPIbvUAqQbRAlGNLGzlsngSy
cCjhu5x1C8Bl0rLH+AgxRVSWzxrYLbP5KX6y/qrJ/blUjYZ2RCYxRU1hMZO2JVOpzm51r8f6fHPn
M6C4lZ6PHQ3fuwRjdgVXBCWnF9jV8W0CboKqmeSp6rkXFglw6nLGiHTDrpca0ENCQxBr2JkKgzd9
bXSqYHatxMwMY4TwHBn3xg6Ssay+o7DOOhANLCfDPcFtG4sHyYaONyvliFIMBwGlf8TS6b+kDcuS
AdDfhPOkc4b3k2ZxFFzjMJV9Xi36ErtMxOKU5xBOAfeEQUAcIZuBPJJVp5Kuv2yjQbNsSS9tUpnH
N9tgVv4T+mQDcXJQyMBy1NPwBFaQ8Z8Qe3k8+eGOH81Cb/Vj3nWe1I8MVUnHs0h1aWju+yAAQyvB
ArqsWZCGgxJw+1JaLDRr7k8L4s3/rVC9HM9fBOskrrCBovonS1TAzz/PVaiff4QMCStbQfu8NVKa
+8IPB1Wzim8kPlgQKXt8cFw9HAD7gi6RHGBCSlc/zxyRpi3WnOSnHW/56UXKp0gG1iixxVxmUIcK
yLcF9HIf4LVqKqxgPl5sBDv+7hd5rdcoUveBqCoF8yEzzpjRYNaRhDd3uxFPZRWIkXLsK8BCk9P9
VlKPrVoa6We86K6BUpE6cXdE7nRr3EIHKvUqJ6FTHR8+zilJa0blJDLrOZkMbyzdHF8umTfiwtTe
8ahMTI3b3J+CFadOJDHqtkc8ucfZ/UGIwNQu++hkDSFpQSAz9alxPMDKhZ37kxs5Nt3W6pcZRgNP
Mw/lrXTjG4MZoPwZPPU1MsXqTjG0QxskdsIFad+7ISBI1SVo7YZp2gEJCDCcszXzrg391QTfuo9S
+Ouf9Kps2s+6/olPonZ/52zvdehHsE3yqR8YQoK3ifh7ftxjiuMvy+k+vXQDI3vw4I0HcfSMk0cw
2oLTXUxYkmvJ/sGWj3gTGQVPC+TBCjUf/WnFfoYYpmnzHXoregZaYmdYdiPFsa8xxy32EmDXIVGN
V0URz9gzIVrxP5eg30gnRNPoBTnzmdg7HHmNZae/S/y+vQyqULdgYenmBmVhf+4i3Zb/zsK1Wusc
+9gWhnLufXR4Y8SlguILCP8X68trcbhbcb81w1dc8hVFhKHekJBGrk1ibmn4HA6/wvSAumUyzhIy
cNsDrTbnP9YURc6g+IVdaod2wmyRyIlI1w306xDyCmu8X7oQD70nLlXZk08+XiH9PbVt9Qq4o8uB
4jgCsXHjfcAMlSKIEHsHriKI5i+k8urJvaa6DYbjh5dQBpF8ohUCz94HDmVZawDJKpveOEmCA54m
mfNsszvDchDKs2ut4CYr8dyOuge7DK0NXzOzym8FPqRfeV+c10DGxTMvT+sg4oR2Z9MahzNSkp67
HrIJwSsZwAzVtxhHjlOhrJM9+MK61jZsPOTZjTX3eY2iwq4KVYaNPo+3XDABgC8PAK5ZIooRwd4v
PBOIU8IYxffq3+nDZt5XMPYyG4DRTieaqv96CShi0pnOxwjusfuobPVV0rYfWHOy9zD9y7ZFtUaL
rritIvFPoERm4uf4io/8GE9jOnsNs3FTUhf1LQsAzSTXceyMTz/ItursX7banoi5ZR40cY5XIX+o
9EXLO93OzWdtX68/kcTUAeUd3Aj45mxaBcBJICree0s6D535lMnQApwNvQp3m+FsVUh5cqUeV8IO
QBhO09V/ppCarElb+mpClZq79+aip3KhDYbzQZlAaWTiaCsPn4pXPx550pzqCL5FXZDutbtMnyl3
tCswvGXwgGDY5bKffKp9sSY1TgLrl9jtj9ClA8sAhCxZuSaSsSlag1YJuf7x0+NecFeb/mt9C6Ld
SuFRLYM3s1jW3YuwC3JpM9Y1Bz/lZJBwXH/lCkZwAGOt/yNv5q9ZWrtvC5B+LD/uvmj+j1aCFxIJ
/eEc9udis6yjNW90nDBny+L8Tin49aGNEFZuE13eXhF9va4AgpDOhipTGRy8/bRDQjvrMl5b06BM
m8O256sB3QmU7q514qR2c1MdA67zkYi9qR51H2It4nYjGCzXDgsaCu6KY34lixKTK9KYP2nutw1p
s1uDrDKuJwO35gtcuhXeAd61fQhQbquN738IItm97wRsqgkfsHlDFYPe7ks33A28FgcShNGBt09q
9qD5ZzgQvnn2gAoauSFFalwTcMFLyKcpNWuTl58lpljyo46erlu0MYs/pg7Z8+Rb9Hy8ZTZXrgfj
+7lTbX0iRd7w8eMLW3ggqC35vaSz3tW+Qx0kW/3K1n7MLoOVTEPqo5bjqWNadGz4en7dCrU5nBEH
t7HelSJ4duvtM74YKkB1r9odp8P+KPpv+SJJFJt3mIzUTyZZuhlXQOu/xHMj+w+tJQDODXxJF9Gp
xQcmkA+Zv5q2SFxwrdpsVpVEhmX2VwTVEEFoqUWsqnTKIePuB6Jm7RkZm46wcz928Lcgj6iIQFJQ
w2hyJKhAJ22WfKE6V9uGInD0MEjVHYlwL8M7ej3KEJB0PKCYhGC15S5WfbbOTUxBWEuBIwSInAZd
IiD2RuvQXoR6TxWSuw11OykE0/QZJ10ir10BreiCdDN6y0JzlfpgucmwcOPO8gbAOegwnjy0Ph2X
tBLkDSZIHYzcDvD3tGXeNixwxgTq2xJuy7DrrXFN2sdc/HLltAZ5RxBC5X0eQ+vDbI83aPNCQNTa
4IOuEwmDoDOZk8RsSEju9vEiH5WwWWJpOzmvzphkSiPwq9KfXTMKP7yl7TzcO7LtlhKYlPezbeG8
xoLslyOoGfK8Se1vGgk4cNUgCuVBZgmCl0uDSLUXeeW5L4OAxnkLEZTz98kMqvYILbstfI9JbaZ9
I15n+SwP5HOWwJ1ZmuDKyc7IP0KRNNgvDxw/r8F0nLaPTHVeDy2mFygTmJnNe8c7MDyqEY25Tcd6
23wGHyqn2LLdhvL+9rMwpvGhMNLZ9aQI4yklOXtyyV6xmOET2Ec8p72EQKL+O3e5rFMfrPxPxiZQ
+bkHwtKec3joWPpY7yP9vxZLomqmhmWDdcNbJ/aqRO5JvPdurQjoJReQ49mXSlvJ08GL7+AV1PDU
W2hUGVO2nc4epCQyu8Q/EekYLVppiaB8J86YiOxqnFb6FzE5186XI/TC3c/KWGitkJBZAO2P4iHG
zYPLjoM9KKwNkn1+LijBe/JjS5YTzDPLy4FzTMtOAusTG3JsODlbw2s8s9CDBgSh0QBBFbHVKGAO
ttn7p1vjFFK/oNYpfZK+OKRdLTZTcRfI4IRWZsVojMChAFIbtdp1QPfMsmT06iDuv3wZibuVeNvV
xjVY0RGVeR+NJXX82+I58iYmf/luByPbg9iLm0Hxx22NC9RZuYIadLQSvdDvY0WOFGuaenTzoNUh
6MDC0mdclgXyAAwqA1VOQ1xYleOwCoMOaV6SUxQDwx5otluQsRUlFLSYnQ3OioQjSQJeQZTo+XJv
ITbbDWnwOKNYJCZq11e5I5XURZp84ggqgp+VdRDHEHQFpLDLzg4hgFtPJBbRmUCSwoY3ReyWbEME
RVAcP0Sg1grLbhznUxkEjiBEKuGLNExwqtO0K0fRhT7zoi+eU0kHCVU0+F/yFl1AFo6CHWKrARbC
mZa/j0ltKrkO3SdzbrBGWhx4CtvmzdnpCffE7WnAj+38FSk0ILpsy8V45UkmyEo8P60XqbZFtN/i
tMyG+A53ZmyPI4t1ahGH9MpphBOemyHf++7VY8lx0RXEbqrdpP84A0NH7XdqWUU38qHqux85TY5B
CD2lT4FFk96ZOofHdr4VDmshFT3TGOlP5IDEqq9LutDlRXe4VTj4vlSOHPvc7FUYHPQR49SfpGbr
CuN4Y/Foo1qhqlXh+oXdHP+gmUW9nM6YBNz4yV/m184+oHQFM2Y5vuo64TTSZhu0Oat/a4Cjk/iO
bU61xNOiDf00xoijfqMYUsAl0xldmzkmDcLcGsns2tMDEo02lIO7Lt96lfofSDvsoRooGZUlq4b1
z+mMq9l4SBbN5JAJNf4kzbFxRTTDVdskYIynUmughb9/D75/6As3iuCHqV1bMSdgAY56m0Stq0jE
eTrP7K4Y+Zv0rD0LV8qWu38sRnOyBP6nCzv+8hU84p4sfjn+/eZ09FNkRsAObG60ay8R8LCAiTCu
+iCcDLcUn751zwWwE8H2XneKWf+nyh6aihFyLJ//mE6jVud51/obgR1BZQsTQXekO+hXqFOtJqSX
h3cP3QpA8AmJFmzjz5DC266sa2dJtu6c8ehPrUWMNqjieIzEwETXekEwOtSnhWMghJsqJA5+Kq5L
wz9HxCyxtvs/SU+0Y9h/3xoYD5rVurYTfQI86pg7vtpoArB0oDIJi1dHq2NhG46JMj2Ow004HiM2
GW3GkF8Zf5qsZN6GFjQ5KEoEQ6pFvm/9Ve7kWA+B2vVBGIhS370FAFG12n3THOgxydfkaQMa4ewz
HGZCijJpCPJuo5Y+8aRwOwVygjNdGMkEM5kAsikKI/s48OJg38MGu7yIl40CKQARa5QZCBEBnFIG
naU7tCB1mjS3xdkmyGrk4HmflEc7L4Wdv+eLy73BMFYxudZWBPsbTMRhRR4SrxtEHkNgYNzuAMxG
T/G6Hh4mMNEGe/XsVMjaxTN/1cwilAolWAnAfW4gh6QDu5cW0SPjlgPfNxi/3vqZCJK0+aC4igtd
+svTOF53DoyhEXvqST/spYrbX3HN+u0r5DyOSMvCPfG9GswfaX2VNE9gR38buLVKZtZ5hHowhhId
5wBgqXydvKNEymJIJg2piORGmAgFffcIBtDy8jihPGKudlvqo7iMs8XZlh0JVqYfpMIYUoPkttie
snN6XeF4Iswl20id0FwZcL8ylegWcjwcEdZUszM34xpsdrQdmCDQDvqViaJsVeqPqAKDxZNDgIsi
nElfy5wINboenW+BQr6vglhb1eqOkxrJaZZeV5ShOMTS76lL5LNY7e1yRLgI3RLFmhA143kDFCc7
zVqcnDcvew9bNho4TB6eBOmn1rFjIMt1tfuiuLErXb4VhAc+ItLXHaSM9g48nxBTJOs2LS4de5zN
tm6XaLSc3FhxK3f+yOWXrkZdGtgHYY25DGLiOZKmpBRk+YlIKcqHzctOcfXc5DWmXTrLIw+UbBBK
vN744k9nqtRtdD7tTRvh3eYtGzuljdJosRHguCehY1+8d9245gnfkXahdstlNZSXWbonCqP0m6st
3RX0eYOErJijt/A8ieB3Luy4g2feGXkHnpGDHsXnPZkZpPPZN3ADt9mBQfLn/6GKzP5GeItpRt1p
Unh/x3jP2VsZPohFWa3V+KSyq91+k0BXgdGJzYg9v7R8kGzgDuIHWsyotxY2pClLdHyAU0ltIyWc
y2jQ6gfqe3XFjY6eHuq8Qh2v2q9eVf4fdrGM/C5X0nTq9cZZPjY8SMNs+bFz26vCPPWuuP+vu992
HYbvXPv45EdlVQPpKTUd1GN2JJ/GGzymxpR86CS+IiVpK696BTbBluCMiwy7guaIm++kNgxsDUkl
PUZPc+G1oI1a4SlJlDcZyFdL0v5m2xOanWMkdWNcIxUArEJQoBqv6g2oeKAnQBH74Sx3jJ1Sc7Ze
jLDLqlhVV+JXyWq33QIivaOkZejZHiqcUvwlM23sxMvGbvDogSZD3xwmnZ+uRIktU8mSXk82bgDP
Eq5Yagcxj0jJKtDT9VElxZKHGqojcD6R/l0EJgV8yD8KtMWUaHm65P9cLu3/Cn7GjohFPnZZUdbD
/6ZkKr14ZTmvQ6g60Izb1STBbNsPBeaPIbbMQFVBVQuqYzdy3LNPOdibLRbf8G/PMW9RR7AANYrJ
jskWak5ORpzhACgbdco6NaU1waHDj8EoHvt0cNX8Ru6qT15Zig8s0+KaUQkHxm+h0rifPn7wIqLb
yXlIsbgF/X0gDkP6s+l4xqUEyJzTE4bhvcb54x+YJTkRvr7cNTiXtZTeRQpTS5/flFlj6dDfE9cl
FM4i03Cu7glasP+nwlpb2yYJKk35kdxrH1zjh2kxfae3FkFR7m7QlVHTme7hWdeN//9F0iW1QW9c
Enj5jPj41Qo3DXWtw2NAyyHq/0+ydboCb8SCM+7RLWgwiRmshLkDVPF5gf55H9DaLB4y0clWQAKY
57cY7hUVsS3/m/DJLeuZkRtcENVHjskpFTG7+km4qMFwuw5JxI+aqsXZyahFUOSi6w6rNN5isSXw
qCly/xD7uMirCWe6x3yUgXQlF7p574hbnGa8XsdOj1hVsy4gCKopcoHbnT9xFj5yIkgdCODokc0A
gS3LV32v68qdzI+HOA/k3N6hyLvitIq1+gM8oM9EAuCZ6Hrh7yqeC0p7Q/rKCVpUMMSebw0x/s5x
TLIrSLmx5XJ6jvOIMPv8u7UWW88/XTbofgpeO2aTVIy5tBFK2IDU/LnkotjZ/QYRj7ClZFvyOLLM
r9iInvFCHOw0iqIDRQOgA7bNNXzvJDiEYKbJpeGORgQ4S9Xl8JKaTy2V1jZz+OU13Uye1+E5kFQF
BIDewa5Gg/9+/6x/Fy41e6nBSRRr93aHX5nDxkTxORutTs3KPl2V1ftr89ytfdcUBwHZmxj66kMd
l6sFOpHpqTL9L1/mRrMWq2pMge8HRyEVs3rYkOxW277QtebD09x2PT01lFbA8q5pY/tyCHth2dOL
JBtAgMUHq30DanjLhT9nJNQeGqDqdLjpQXBi5xIDXI2EmwxEI+vrjJjc4FpFnJqQ/EmpgxMc+9Fc
o2zlFcq+uOhaMFrIvIXbG3RrxaFFJnp23CTmuFYzRM6uvOtxEP7jtfjWXQuaeDTEsiIhI3ZAR4eA
5XmGD6r1BeIi0gpKyaUvO5Bo2YT8NvVefFq3SBD1CxuCn3tP3Mc3x1HnXOfQ4FWV2Se96iME3ZaG
5kEUqrP8le/31bDFKBQav4L+qxQJBMiZWj94TSweTYrFHE0QrJMjX2SCb0uG4qaDKbgqTCtzV7cc
7zZeHPVcBPN1HrUIjd5anRdztohmAxY2ybi6ZkVOj0+ul1nf8+RH6TC3SjkSQ9v1gVrOAikiL4UD
VMyoWsCVfpYt565w44+y/12+UGxkCD1viY1eyLlraYX8EJNROBZZ3e35XTDmaYF8JS/J5zk6Mkqf
1poXvU9T8HFrlHI0poKik1Jbk2CdC8HJuiHzkJRiGqjjalfk2+xbZz2COmQJ5Yq3kOPxIe+T8DzW
yQ2OCNtru4z4ql6APxjACKFr6fR6YYO2mupdYXtFS+rrLJj9rbAwhmnBf5polUBpsaorgrytB6M9
Md/QYY5Xr7Jq99xIB1DcbBCPBvAX2jkoYW5NatzObRPWBuwooLD5AXbWeDvUPRTGZNuH4B6FJkHN
kdT0GYf/pxn/z3AgzqPJvpAXRJpSwqm3cQMLwEhcTAHngypyzlglMErSoRsSCQQBAV4pbNDt9MX1
HKHkKCd6oYRn6+wHqmvdciBFwETAGtgGk8nHQrjHrhkPFqhi3evwo8pK6DKwteGsOQBYkxL8o5IH
Mi90ZtjpbvFpwmYd+c3k5bLdUgl36RIn3lxYxavbtoPe/pgC2MAC5PXnPFwvWjDFpkEPV3VN6ejw
y03MypjQCByOAcTA6+cpHYzgmW0sobiWk1vBzshS0ZK67MhYhygiZXnvccI83UMZmDGTJB5jsO+w
DjWpux62kCy5QAEyCZ7GgkSYenLF2K6uAQAdX469lcm6x8zZnL2kfOA9+HthoY5uDr04cpG/vH1L
19eAPJyxhR6LabWrnVnPZ4f5N/8HcyaM55zvp7Xruhxfy8dNSuNEVjomIwwRA8mqemhGRGvfhSbF
FypNZc+qi4LydJpaY7FuzfvrZAsiNT49g6Rk/RXZsQVU7kZ/xelgPTlihGxR5cWT6sB1GqTqtF+U
Do2gK6JONfp3rb6FxmI9IJ3l/HOku1zCpsNbejG/ZKQowk5RoN7NSWRuW+IZqCKGE9B0G2ZCsZIT
vpGrWlLGV4iiqa1eDvddwJWYgkJnvUsL/gsBeuZRmym94IKCkic30ajEGCB3sNPtWPBPQLhkyyoL
wfGpEfTe1W4Z9ZlgoCh88+SU5VyqffuSXp3TcS34TvRdTsN+uPkip5tAR5faJrVJwMfF7F8SipdG
ZabNyrRiHdBnx6Nx75NJ3fSAnAjBrKST2pEAS14w9n60tjPHpvc+r/RBy7RCzGrhEGIiHNB94QA2
RkAK10ukznjUAkj6Y681yqfYzbGZs7faqXTT/rjgw/RG+iYPc7YSg+Ip43vZVapzghLk1p07rDf1
jV/fqC11U9YsI/xto48IZIhFrKsnkpR8hEtkRAA0NpN+poyRgJBYiy1pZ+7/821E3Tr5ig1bY3EU
JEzxYzYMVmtjm/qE+yOU2HjOo8MmcucopomS0Mb8RNHz+2lphN0r81HldKvrwdAyUJJmTbudxChm
fawV67mjcgB8JugyUC7UM+neSbu5P2LvR/5QbRyn4d7Ivt9OoBZCh7FtNXi57Q0VLMUT7mokd44L
tt+U5dS7S7RrPiOxLqwd9RtVubiNyvJ5vt3rftnNLU7wmUyhc4+pp42ezZNb6AnmSJePvIkM3G00
DV6wZ3X3tVeVjCcohmy2U2L/0iVKJC6p+H5mgXfFoV1+vIgOYq8/fdc2/Zc3KMbJYraAewLb2uIU
EHA2TNtFRTGDISNNioNTB8LhmN1IItJgyn15Vzb7itV1JUwj0c4kSEHQXnG0g6Jrl6PB03B1SHLu
f8VK/zeVPZU4sgypP1HJhk1mz82z7Xp81qXsbLH5jn6GSqcxzIoMv98mVDiK78xPwLappgAwlYXR
g8VwnWBN9C7Nj+O9Cv+GQKgtW95Lqkv9wn/5NwBRtJ54ejX4/7925Zx1oZrOSWkUkE/jcTV1VmUM
KNIjP89LxDUm1s7rwAl4UaVOF2diBSiJRLza3AYiOMpHtfatxu1lQhfQWxPhZyzTLBaE9koxEk7B
m2lAictR1KrBYBHD5DVljIR6wwrZdQX6Zywh6dcp3ptUSeXxTwKev9GJ8cXBLnERz/pnE1F4PQWK
cf3wrov2oWAGzNZVRIvkAi6y6SAwhfie6Jmma+KMovIFt6OEpaMtq+rIsWXsgFmDYYuh1OQz7UsB
QjL0HAzH/eR2KCw04K0yG9s0EGQ+CmpVGYaoJneIxdu4+Y81qyd8LlehFiEiL+y5Ux96LKQFqvVA
T1xPZGM94tYI9I319msW1u0NtBs4emp/hMxzFw2jLFBjd4QdlNLIC03p6WX1ZUIX6C/K+TAwV6l2
aFwQDzdyPPSD2kYkVs042bgfDfn5BeWfsVd9+TwzPXygIhKUWX4FNgwrHaVUQDwDHJzDXj70Nyjb
UkgxCi6eheNJOvPdBNO7UuAPjn4w21ViwU4A1LspddkdOZptV0XY78+ra9Pc906Nn6Gp9W1Rq21P
N1t32sJAXq0qERmxNm6r4SaUP28IAhsADyxcSDJJUoTEkQY8VyTG24wJ8zCDSdE+CCh4KpqFp4/S
FL0DkEBW8SM6cRkjKkV0NOxyHplFRgMiTSuiRGsAXsfLwspaIt1blF6Ma1QR66yvBOKBdNeKnItW
RV2NfkP8lz+poIdIpxDqLLTgoyq5tIDnudgerTQxBhSYQNiKYBf/ZCUIDY0o39ZpHSIKxFshEObd
LFAXX3vEPGTrKjfYYXDkiekZYK7sUgRVMQoNBvNLl8nDxWRV+yh2xMFWWdlu9xDeha7HgonUc2kc
nL8RxXhvtS1bjkAVSu2303E9lo6dVb5qkdsEp6PQ69eGFf1kCPzNORiGY1EpXLUtVdEaVmzC0pwH
Rv0evtE6pPiSIJ3hTGWxqsdH1JqU73pTRdwJe7ePCcmLzoFCTgpHk5ll7rCcFEi5FTJjzVvhEK9q
xlhiTTTNc0qsWFuGEbf+1xwCg+mxl/YXCYam7Hq94VlJlCDKzlt9bdCE/KtFnpmWX7TUqtE0c7cP
FGWb4psJFUVzimZ7w8GrsOk94pXz1kgImTOvIfsb5SbEgtgQBjslSLXpjQRnhO4FtCK0imbTGaRD
U9te8IrMB3vxigEHc1vl/mvLhJimQlEx83kF4d7kK1t3oBx2cTKGhIqJeI5ktWXqlGJxdbCPvtcx
1Q+efwhMEhE5xqdDtlcDTn2UVLtuNthxG3cQ9PBzuObX9KSRXYOPnTpriJ+o/f2jz8T+VXRgU5Vw
HtUWd3L3bNE78o6eXRGdXAQFniiCdfLjKOWCsG/3ai0SAyDyE3x2Uk6HmRXHiDXXyS4Ek4AGHqFc
c0t3F76V9qCyPhozh+wQruqBIU8jEDl6Uz/HweHE70kS17Qz17NSw1XpxV1zZpgxVbqfGfvh6bk+
Fg8oIYDKZ8RZCuw2qPTZbwnxSmh9Ofcy+uVyMI4QwwJdiagi5On2s7hndnzfEDb88Mb1vyMP1IBO
so63rJ+koZor7kPwpylFEV0fux56+2W0T3QaGBzfQXNcSR9tFQXe22gBiHvZX9MLRbMF4Hpwv9r3
PT6SXUMb8i+00Roqplmcds9Z1RIQ4OKNBp41yHdPnMq8zyLNPmr8IPLnWg1MKraAKyWyK6B4L2X0
YXfagH6T8VI/vNNpySLzxsivjCXMeokSWQdRorwAYMyV65HsH6EpFrlTJl5dKYLbLhKPwV8omt2u
3Qsn0RgTyr9kBPQQDvZ5TEvxq0EOmvWi/0aF8TVkwEqToBKOalxIfcRnevwwC1ZJozUCguE3eDGs
FzYjG8ed7UrJPim5+tcE5v5ocmTyWltTQ9vO7WGgGkOVuqHjIgGpJxUFUtTGxsY2smoeGKmw7WLe
ZteGCZ01x4h/6wWLch/AY05Eu179CLfCLoZJAxB9hH5tCx/BGN2aiAnNEh1/2UgbdD9gJJiH+I3c
4/3Fmq+pPaGxSSj5WB+do0UWt7Tav4t4XEUwfiyqpSSZtSCp6h8k9O8s7bBbWJcA3KwHuyqXAVJg
64bAMXAchj6NV3RDKkuoAv7CeYpP4/VhxQ52ldFxQC/bYVn3zafOvnSJ3TENn1KM4chwaVhpBVKf
fPEzrMFEdoDzl7ik9uU0nR1FZo6wfG4q6CGTr7q6E64BMQpsAoPcFMp5p79xPdO/GIQBggDN7sVA
74F3BDNyMqbluVGK7LfZGZV+yHT9fZXfnGRfoEfCZ0dOa0BN4674VqFP+7Ip1pjAtIJGa8uXIwWr
BWfmKqhyJng907dJzf1VXeq91S26Yntc4rZEV+5rS6V/g7i92Vuc5X8j1NqEwdYK8/OxziNjrir7
lguqAeZJRNe2wyUvQ84kvSMujMAuooKO5LJurf/1vWO1PfKOj5GaH74bhYQ2qxNoWnbq7vKg6mni
YV/j6hVeDzqGLco2qZTxYFWCCYKX5gmysxI6ri5dy0LgD1GeoSolrZVIfyJao6yViNPAbHi9FD1b
LvgG1bsQtsgoE+tj71vVQp87901QCHdkInG8Cm6SkFa/a1uSLFEbT6Fw5lsGv8fXsiKL15r5/FVC
QRIzMMsw2Mq6orGNlfdl9I3WR+rf3OtuipugF8sHioCb/k9SKmuhV7iqHCliK08lq5PiTmHYbO7+
WZHvjoWFCN3LGMlL+SNmzpu1wVPseKy1+hnTYeIonmIV1UmNqHFcygytnYs9KJWwL5r3XesYnGol
uOXfwDqpHcqP2ZkIzsY/dsW+tOqiQjtb63lizI7CevaX6IxP4nA3cIdf994bC7NMcjlUZslgKPuH
MxZYhSHurDefww6WUePsEOMYEtTulBwsqPuqEFY3cXBhdqFCOdGaDnK/OnKmlzBJgyZQsEukdT0a
ia9ZEpVQSklN+XCWjpCKwq5LjMgMwAt0sUKLv8jJdSjFLM4n0dXyW31q3ldfB9ST7xaqWJg1+Qft
rbhXlAcPWmnhR/EACXq6kip1+0vmScVzZQlSQQvSVWRXnC8Xh/dQhy+cxCaLe59r4QwcEugk36Jr
o6fAto/2f6F9yxsfeBo5uvLXHeqs7le77KAqFD9ejv0JtVW/xoSfgFMQByD6BNIVO3WJrdgJRPPE
xnAs0SiopF0Rrf/2N97KCaBo2seZMplwyXKoRBoWhtu+1gDFCr7wE1E337J5AND4EWJS2mhaJSYu
+AwZ+SNmHJs//8HAgk8WfeOwGtFtZswcOp5g7atrIro9JuHokP3gQQhy01e/wHtZ22EuCfmIJUhq
EfQ3eawJ6qOiXtz1qmbXC6mD6owhf7f2NDhNZJvE+FlPUI0cJSj56mrW3aWRm2wSsq7u/yJNtwzD
DQl8YitN8LIY1g1OpF9+epJVvBCaZPJxONDq+evDbMPDSyKrI4MyjbtZc42P7qGsifvXOq2jr05H
rGPLkarkRZT9pl4G3tStX5Mavs5wHoEGzx2xawQVT8KZwLJRD9g1q1nXO11U+vVgoLz4aZe0h5YD
GvZRfbPCu3gDMksgj39HtXdgTpttG+XxynR4C4aBi2Q60sRU9yDrim8dXX/mXSptNIhZzuZJSlZC
87VKYLqvucbK8gGTS5Fog82VefeF5i4Ispb3i+gqfcBZ/bzckrCaDGO+bXT3fawtzGTeh9vD1k76
iJRnXqJJYsqT7Y4C9NGwSfC12+/MFdKBIHOby3IdKZwYPr3d87VjEZ5T+zpL1HJKL3ZymnqRWnih
Jqr4nnBRKS/8Jg+dlvC3BAl8ICzf7zbxnnEEBZuwvVto3so3U8d8Ad4/Vd5XQXReOMuOV+urXe9n
LP+/ReJNNusIb9U16s1XYcBQ5KhmM4bul5Mkbze5cmhXFu+bfjTrZoY2wzTppRvcsjoW77V/VWqt
J6YMpq4XMbnwyzT+vS4phHHpyeDQGsV1MLmQf4zFXdqpO7cUcBENiIs05XHLxbx+c1rHbkwBYdiY
J64V92hrWpnT03xaU+qKKKMy6T1WiEJU+IbZ9wvU5hW9/BoYjCgqjikI7JiHfGjriB4uf5eD60d/
mQcJ1srd3SCQdvb9dLBDy0KC7VqLAQOdnaGRjQ33FCAWSOkPV5ZwHEpyRbr7ZDZWQWsXIvc2HL0a
0+CyvcSoxVi9lSQEsG2TUHN3dKceiQ12Km/kvMm36STH+GYWcfQH8ttgRa/SYl8q+48kSxFfEC4w
IKXRfwKAfmWCwqi+DVK1Ataqb/jy/A7RRIUPgpdIFqrlHYQv2a7vrGWL5THVo5B7ruKDOXXSWibt
5Uol0Mma5ZnRYCmJdBBO7qbGnNuVExGo4YdYgBilS7zpfCmQ6huP1u/oIlkX/VXUeiGNK1IzvYiq
lbJhxHAIdCY7UGxnXmga8gbg4wgQeMZMQ1SfECPxoFmgB1EBKRGLDaohKotKhYNGP92HTnS3Jh8O
fBRyZocByuyia6SJ2AdMd4Jr4rzv+oOlsdZbddP74/wc7xA5K6Esqkloz1FrYbh86MHE8omF4MRd
zH10Z9ruSo6WUu2D7T63bf/+UPc7LrdPHprpJCZnSWiBpGdFRY5AnVOX5EeCKLd4vFGC8gLQTa1P
YICnsXscCasKNjPx9ZjXQHVplTESxRU02WrjjRkwX3D06bjgdsQNkIQlAX+ifcoL5tjIOlVTue7V
BVreVqLoY13nV4tEAr5Iw330TYm8wxjX6che9ZFZ5VMPP72ML52LSPv8lz68nAGGSFAU9aPS7sZJ
lSErE7lag0ArG11QMGs/sKYw5c8iMEaWvTs/3Jh1Y5lFNuoT8DoegOxgF9TqGkC07yqCjZCdrLbY
120TvDpoBeIbGIIXD7VYrN0doIEwuRvy4XYhQ3NcqToQ4Etv9/Ph9vyHk27s99z+3TFiZ9v61F8Z
PiqFcqVhFYhdreeW7cZr02bcAY/rfPumYAkNrgfK8Bdz822hVZls0jjBnIHBV62MX5zzRP2jO5dc
HzP+x3+0oDLj+eD/M/Kc7PLSUpac54XLzAfEZxoOFTgV0ZVNRBJIJXcoz9VmWvgxf9bKLrJ+R1AF
QQIPlE08q9HtrUP2S/+XIa5EY9dUfVe+bmad7KcMmbj8WwAzcdNUW/ImEO8WJD8PPlQ+iJqE5zIG
cimQ6itlOi7h517Grn3EkUnTncFfUByQOft/iptT34chiMTwnJ59+UFabh9RRz0fYa04uxOP9yuW
eaRXF68JbmCr+bkoNkMlqpIoJKk0PoKCxY+LStBg8CREu78gsMARrze/IgUVv7gMcTKahCH7JEtU
eX41qD8MNRqGj5qoc6yjHGIsBxG0TCqy4gdEcObrxgI76GjR8hzcWI9oYtJV9mcOIxfCWk8LmwmT
TnfUACvMZl7nmJClA/KwOypwWew1bUsDTgjjTHGVpwjuGrjt1RrK3V+4GEmDvTIY0ix69/wI68tu
XtpynrwMWuKM+HNba0YJp4GusUHR9Rpl8OomCPWsZoKCATt9NIuczSnelac4xHE/48JhweFtLsLe
Dl96gyBI+Ykgq74kmlLQv8sUY7MuHvmbLkEA1NX7t1Giq+qfKvZ8XNdX+5IWdzCDvSxJQBlbf+Xh
hIEE1mvp6jdF85Dcbr95v6teRNYuCowdjmsDR2Z6cidUsOYavX41rcl8kP1tMiXPp27cHwLDGNbT
gOGiL0H4PazO5mL7F/spuZN3Y/oEEOIEkJYc8a6mPfi0IQ1vHRhtEiDDDQe20n6IQl8yHv/Iz2MB
jD++wrXNVL+lTUOkQKlr4aBqmr5WP4HKgQ+m3m+Api5aIJxYccwcOf162IMpemw5wNBAe/RiGaaV
CPtAJ2mGyoW8vMrFl33Di1j7B4J2uECef2GEcLwDTYmLvgH/K/HUpHheqHDlIADftpAy81ElS1Nm
1ndU8yD2WpoTVDOYy+rv40uzlA9o1l1DJdkeXYacvVPyhto3P7grw+aCIyZlqEOr+cGmULsjIeMp
aZlTARb2ckvklNcbI5o2UJ+k/PcwYFw88mQFO821kwni6xn5IVswW2/NCiHPkCW7pUJPcCU8xRjH
02jUGnyLakpfkxKJFSmYia5H6TXCbiIS2FAm4q2KFe7QbKp4BxZPB10VTFMhGUPG3BrEQpq8D/K8
NsHYClTRYtf46+JDk/J0Zb42GOHYaNvSLR+Uswb87ieiszolQbFOkD2iWGjCg9KwSafBqbx5QH+Q
01r27fxbYh5jukSKeLT3G1PbyX1T61/rpyOf15kn5jrM/+oVIyOxSQ33ZOvXoByes1M5CfuXXgh2
0FnHoHcN66W0vulIZOTKJOupbKnERZ/OFNQqh3D8BiuQ7V1SwObsYooCx5Qjq5LsUf0ULrABCZjY
8mmGzvwyNgDoKiE0ZAjh0DxCcL6YjijfX/jgSPMyPwVGv5VmmjMA4S953rE2Ws+W8n8EGMkYO17R
Nq+QTWqqynhS91IJAHqd+146psTwg10GMF4lmKbGiVhoEN7RIaVKUC8TNopIF767bM3fPIgM5JvL
4vNvjQxHCgryMakGohhkrGPVS/0nCkjzu1aHmBr0LlKaDsHJJ0jFwZiKtEnd2yAddegEY6GOiuE6
pe+CMpT4fmk2kJ4a9lbGo4L+f+zvQnWfwXGNrx17HpkfQ0xgAXPCzQT38RrKV5LzU2mPXj+46YQ8
3PErl4AuzZXUfqcNhE73Cg9S4Nd6+GKoCUuN9N+yOGYVKkmn84o1Ko9kzSX5TDY8I+XqBkWtw2XL
ChfB23PinotseK8n1CbajJQ+5rZ0li9mENP1eY+P1sIX8QvyQ6/bswJCZ/kEwLZc7dSnQaSNyEuX
MKEJt63i+woeLLD6yHNB/s/9Lcj8xQDCujByNq/WMNs5zxikUGuStUBaVgtIlsncNz8G4GTI+m8N
eleO16fQ/r1HmUC83UgEzHRf1poovNzqzlTy499irpzJTNeovJ1FHG39KEsJqk0qgk93hCW7jYzg
CJLjSRxjkS/1stL4hmVlZ3J6fK0FuNWdMgA7Yrdy1pixnhm44+JPbQ/RYvxa9PqTHI/CB9CVvZR3
tN2Embm5TYQ+qOcv5MvvJ3nVi/1l4PZUb/UjQ4TX56KOyRO79vNilntNRqxWqYkTZoNmW9pjqgxf
Uav5YmZWn3XdbMJvN9UlXzj3+zJpPO++SHWNpjNc32U1vvoi/R4OY++wd6A3Z7RU3GvdKmlYPc3M
76h3h/DXjVmSxImzJ95ujFBWMVJ7K9DGMBoa11rRWd8Q6WCmkKp8eS48g+J5+GsPSIkjzhWu+W8o
rglrj7SS/UNE6FpdwywXAG8fstYL4yb8oqZFAWptDJxG086IciJI87QXp5GA5bgyf3J3mGe1J35u
jqAI2uSRBcEWOJCcahu6o2QXFhdsmH6AXuWjFy6tZ2tUdOdBj9PNglDSI54npSWJUVpeK0hEwAEw
HFimGNf8Mo5hQR1Fvl4wT5QJTkgRTZHkrgdx8WvdiyP4xwG05A+Clnzt5A8e10iNCl0FT3k0B1oJ
wabi94y0r4875uIEPpbAr1Gz9UHtmJVrbhGSM7W1iHuHTtRFlDWUDaWU/vgN6wLF7/rxyAYQ7+68
yw6kMR4RPSpjDSmZEWV8abyrAMSnCuMbNLQgoSiRZLoV6LHSQimuwFHXa6PAcpYnQOnBPn1CnxBq
Kk1ofu04yFb9k7Wzw1s/L2YQi6ES6lbnffOyjA1tieYAECw32WFDx/RqN6o0PaLqhFRFKSFzDg6y
S7kITmRquOy/WAi3uDYA33BQa3vyOvQOiCCsNqNLs3zVnTE5b1jOxpEqxoWJFm3GoPbbMTFOxqu+
U4yCbu6JFHsMdxiTwKD0PF5dHufvD0gz7rNM0fBplILxvLqiT0Wr+hI6J40JF4Vmewxd5OnEqL5q
r7H6pZv06+p0eBhCC9FpZSnxwEpHJ9G0kH9/Q6tAZ9Wi7KdIfugwZV4ewaokxmkBP0HK6wRc7xrN
g1yGI9W4pllGr4flRhiu12jVEzeHQa1s5bHUDYrgEOJnSuQ01JJ7W+Vzscke6NFY3iyNPBLLesEi
H22UbIrVxwWgjNVWSNGNPJwLw7cMR1pUyFoUK41BXVh6ym/RdwjGh5s2nYXArh4kQhOkW3LgWUHk
9EqSOq+WuZgfEzp2/vaELDDEVWT6scYuOv+t9g3Bv16nI4lzFWeX5TXd7z7MEMNwmCunZfzWtDXz
Nq2z+PK/QXuTyO+jF/vQpbBbkH2MsDoij7XjyFmiyi8CBvw7z0jcUmhO0Veby2JVtBVQ4+CxshNB
bigRl1ST/5udutiK99bn2bjOLlhVYfpWMs6xMHfBf1ZcXog4E3mOyHZlQxnVikCSXD2Pv0xHAYH0
iMY+EME81KCJm4cZTaXNlAUg9pFvZaYYgQaD6tfPWCbZTUxEIV3hPjpaiL8c1UFgiMOCsqS5REEC
13si14Nc9i6XZVPS7FaPGAkXUIsAwhilMYZh6Y2rjte/mahoktl4sjSpKNKlwUbE0Qhsl2ZH8TkG
wFzmvNInLkPjpClw7bgfAAhKftXOPDfjox9BbruOH95FOwmcfAL16U/za1K5FE6HuwU9Po7mIX8Y
2/G20J9VqmhAVs1M/+MIN8YmjVuNC4upeuIRA6NK6XYgn8q/WfGiOnqJCsG7SFs+66HXXQwhWdaB
tKWS04moc6I9m2dI2qCBFSJd9DFS1DfbopLWeQZTtxwP68lsTxliEGaczihFMgF7hCWyGTzqS/vM
LH/dRzQV2PxRt0erlKuLn/7HGTPhUvMqXQmnmFAo0fWgFf5pkXokVfnpKRmh5e61qzzBMd3Wm2Ts
sGE6PJLDIjAFfotQsOE8IxlmlUSAxXtx+nruoIbjM0+MsNX+LXxnZQXYDirb2RJTkjgsOimJWpjX
QyfhWBn0iXtwO3ll3ppqirI+gKxdHkvNMaREtKUxuPexbg62i1Bhim9FJc380g9GhyyXg9fhrXaZ
QFdHXpPm77w+lXnwx3pL7iTomKoEPbUSED9q5Bq+f/0PXghAeeDHJFNTlEC/r/AqbWrC1fdszpLt
aKxQGqBkoqbWZejFbgmkc55rGcmrgZmNdQUwNffe/FAfID/W/iqeAtrlR9S9avjBbKQymIx5EAiX
d2Xhw+4xJIGcvrhQTtGLtgulyOAIwNBMRFdb0KbDUNMdkBerU65f3mJ+QChI2Ahr++NDt5UJy6hh
uS+8fvTlmo7CyD4/xQWJfzwIWGHuoBNOvvMu6z80W0udrnyQr70bD3WIppcqb7n8HIZ9I1k1SD8Z
SuponeIOvU7+0ql56nQQTLVaKM2zlXOM5gIk9ePFW5FqvvWzCSpCI0hafIWS+r9xovPsDmwmvk6U
V9Z6YFmdjZylU3uqqnzeUa8emsGX00i3PmaEkaYIAo87TMldXrjUEH+bChUsUT0UzhjIelJwzAwr
o/klUblTcZA0wx6qsIeXOvZOeoE6YMjOeDtCNOvdBbyz4igfFPpld5DydrgT3en1gOjbtSxgShrV
9xe8YNhZFvO+kqswyzzKmQDmyFTGoDosSKIJFYBBGdL4idQLdd+wFb1WBdFoRVs2+W2dZm7hVelt
Izp1DVxqi/HdJPEgmshMzV4E6LUhQbIEKnUnjONCeh1AhO7z41aUhfdiFjpj1l0Hm08L4iex22k5
1d+4Th79BsNaQgsO4KYuNgo/BGO5Qj39mUezmlo559ZdnNEqL8lme01lQnFBfBiQZphxnZfBl7+6
C3CRwyae60IS1ioMzLAtIG7PtIymBFrfx/CXEHlSl1/5mRFhodx5Nbke2p1RVyO4n9w7DuD6BUUE
u4YiZh2GY70CAztFyXtG+PaVOSo/y1p8TzNQhxj0zs3YVyYc3PyoHWADQS1d/pASg8QwPjKMRcQp
9WuePN753XRXHQQzBRcSOPVfH5t+olVDgR3XldLGVIpcagNj8lTp0BYufIJ3qAJn6kbJwEIRy7HA
1/XKbOzDTfRG5g4lKPfZFSPEDFQ0D0aaqbaCBD5QE5A5ZcmG4Qops6+es57cDoBrp/nwvKm7/KjF
FysNdjqx5mPNE066KuaiC/DNQCeoAuLsdO33mdmhkzuq+iqGAZbBmijdXvqS2KfZpT0ALUs+MmdS
H/YOWKgy5lqQvgDmTUtf6ACJ3AqZDrV2FO5l517o+E7jZa9e9yJdl0waVbZJoLJOVfM4aeJ6WHYe
gb1YyfINXUhJbKomzl97N+4msoCNnzPAW0bz42J9FD3aAhh8UgFTVhtgV6uxAn3cyrUTb7HaDRdt
JTQ6KPDkY7+JG5zBl5+abfJZ2E/77/JZ+/VUWK4STAM34SWpo4Y/P4FWNlydrXiDZDgbXF3sJGIH
8vNVk5Xmfhcl9XOAlb83NT/+2OJDHoTc9mgwuZHaFTJL5jSqo1Uv3qShzqBZh6reGOjI9no7zOQ5
BFomuBs0x+S2SFP/g7KD/wWDPRmYN6TD6sbM+oBU5YcAWHx8+oLy5pd0gu3+gfhmc/csbeiLrZ53
vl9uhUixpPADwUyUX8BJuH0DzLXvsV/bheXvhy3Mue6qhXaAiFhLP6O7NIe5GDrWuX0yCSBfZHjQ
OFyvKMmDhBS/dpYUm89Rr0o9/Zv7sW0p5X2DKIhNhdOZb9gEsUEJnRzUfNqkPNWTsotPjeQyrpbF
1F4irp7TAOgJWo0GPwHZt2UdH0uGoKJG+LE4fn8kmTOtbdJu+NkBUp3ArIrYX5iSgzCT/Kz52Z56
jUXRMv6rz5zCSqtVTEItAvQgrZQ6d2R1EKXX+YIijIXjQZSoV+1iAgVpR3rcMXvr4jJFi+by5ox2
SDizoA2s6JByUhgzagJDEMEVTFD+0dvQ6F8CK5M8+DYpDG0YMrjFR4SpkkxwDLZzotjy+DtS3P7l
I9lcmM5txAOtZ7PjKAAA04J2IQBWn2NYdtMVQ7Jtb9TyJ7DwSi+xrVw76xSijNePDLPG5QgLIvH5
B4xr6VwDnrIa0zx3PuygI0nPLM2tFrF1Zj8uEZBDejDJBnMvWQ2H2/aIpmGYwRJjqxLpAu1M16em
25nU0djZ5LY1eDaVxXJYhYBpuT4dYznMcpfkXb6Vat8eMuAext/fjr9BAgqHU7wlbvzluqHHJYrW
tvbKikL4NGtGa5SapdwSAbQaRluzEdNdg2Uum0zhZ9kSBT7llUIiIPPGG2gJaoQq+lpTFfXW/yAq
hLMetdSHJeAYiYHPsnerRROfikf+TKzGJ1z3qNJ8jOY1MuhMJtInvZZCAGZaCZpuxN/QhCk4y/9e
1iiL7kk4pogQ1mf9KDB0Lpx4RW8HFukCmMJHB5i9D28xgcgr1stfNtC9MxNIq7AGZ5KITuaCVlQ6
PHNdNi1D/PZHotobbCAlf+69l0F+0XZA4AEC8HhveIB/lIum6uTFN1XwuSSkk2AD9rx8+oGjuZQn
7cW3leS1f4QVt5W0L4DByKlBvi9CxLIl7OOMDaMPp0cykb9mJbEebRgxbjEH4XXo33lOinUyYrCh
SmTebhtA53hBXgNiutQbOQh9MotNZ34JwTlpBJGCqMPNYYiXbf6ZMOuGSvWFxM3CBN1D5xclZYpE
w222zMh/Ost0yi+ZlQqQsGqP9SkMGm30Vp4BSqp3vNiAxlMU3NmWs5KEhVZhw8cJxQ0hRcJYHUiD
wJ4CLlCHQpJExWjUx4htj3C9fTV1gx3HrkEIyzWJwKSpOcaXjmjJHr5R+kkUUIXRlivbNYvXll/U
mD3eeUed9AwmpUfvxmhpxf2cLb4/TQeeNJ583k+8YE4A8XVfSg5tzExnzFzj7sJNcoCbud+5+IQ/
39bwiM7SqQzf7EVpB3f7Mb4I4YQ9IOwW91/xXmqbbIuSiqR3rmWGvhjnZECrVCZVLz6tDKWXLbhj
reOtn+xgxRZRQLPib4VSuRpdwcLBzxo7zc3slAd3ZDN587AZ2xByju01ufv2tJ4A2HtSfE/ObKRS
i53dj5YPVThy1KydFRJOPbD3hsgXliL4ISxO5h1/eTEXxVm6VX3uDmEIGhYA0RrRW7AEooQxgv6+
rVA2kBcqpa9osOcjevcDcsR14K3UP2y8YyB7yFxAzpQfe5YhRICgI0vEA7PBlK0RbHeX7VmbaD72
WXY+yC8cRFSscJzW/3JhbiX+j+tyIoV9Bq+boSXDW4g9pJBEluJ8hKy7Y+d4X5TVJ6VMqJGra3HY
V+ACLw90ttdEGf9nKuSDn15+aFeU2rqEWnkekAWWigK5qVOXasMC24r2tQV8dZv9uhRVHqV1pI6a
21HhclpUaGyNg0v97PMP4mcDNcCSPS7+hmH20Zcl476hDHsld6n0XmH6goGQ/G5DYdPunDzmdmkJ
xg/VAl4qoOqwFISU53gtH8a8zsLbWBCP/SvDusGe2JVcFF+mvBJ/0pRiwuO+WOSI+s4yAZ8AMZNJ
R34HgMJwxomXMTg9t+hZfuHrV0rtyUpToLLkW9zPYcizokjX8lyg1ZDsGPuMJaoGhnv8Bc3QMwtJ
v7hzwk6fnrzeCK+isxg+BDwsc2p6rGlBw5K+gQMkD6mc0WAUjne4CWl/RPHmUBwYgBT38/mmpy3x
2o6ugTbgxkVZ1DI3xKpoR2ltzlan4OSTtFIwEOo02yWBfShtdU5E1LyDQr8F+a94uInBXABUrwEg
vqZwj3wlbmhJzQgOIKOvP88CIOP1nqcdUunBTnOL1zJvUbSN/1DBR0P3MJqGIV5ZJB8MQDUgtT2K
HVF2QqJEzC1A0wi5PHtUX7PfeFEePmq97PjyUrDND9QsBLSVWUOIjuVFaPm25ZjwNo8hDlt5Y8aB
KC9vKu6VthfsGe/wdmsSxLIWMI9LYRr3W+afmnOEWPAfR1wcbXdvzCRdZRS+HG50/d/d5DZy+nc7
CyiJ9/WrTYENVM5ZgQj1RiALeu7HXbCi4ICsHc60OVPiKFELaImRvBwUoU/hbCob/vIAmgayafrr
5X5uRSr1bbo/B4KG5VFDOrf+BR0U4nijyPUgLtRcu3/gh64Z730CljWp83hwAEd/ZmB9BjtpVaPr
lzMXGtbvGZN2kPqQ6WtkV07LzXt1BgCpw/AZqQkw3q5oN5tdD/kwbq0dcT7q+sM7m2VY8HswVJnM
DpbXiOK/IZutUBsQN5I9eBYss7O5i6uE9f4Ij4LUMp1giuuWDvgc/fGWrjLB+9Azg5VCBSH5STFq
rRrAmARIxVHiXertVv3begxdvTkxASV0qb4DSSKyy4C81YUXE64jV6WivQCdkZDqsbREt+EnRBwK
3WS9D02qxBs4HDnj6Kq2AxAI6QDZe/iI/67eHOG8iEWQGzbPtZ7ms4p3payGjyoNvDm6DRjo3nAI
DO+yRdMFuCxKs+MCMB16t07Y6B44wyxDuOx+ndmc6jW93u79D3FA8M2DvVKvb9SqN5/4Pf37ADrr
+TlM/FEoz6Tj0+euFgRygQ32udcbhjcPPwKsbOPh5T7pZQVLEwF+O03SHFE6hDB6s//ZO9qy9tym
on0ng/KiLZ768v+LyZ/hhs6hmRpTpUK6s0uJ/DF3mnE93+KDKFLgmuN4KeYuoO2d9gLbBoZshG/x
k/4KKVmSUIYvbY78VgY0Tu7Gr4JpEZNlBktNUHINoq+kUxphY4rtG6JoeoeSoiuca1m1u0WB9lj/
UzJNToFjgCM5ULoJrF03RogG/1Oeaj4f3WiXQ7zm1UbqAHmcOczabg6dHbyoEm2Sr0m8OnHo8f1o
iIqdZBKISseyHCT39TIKT2FPubHzSpnBQp7p5kIF8aiJ3p+NQrM9gtTBVPl+Tz7Xl4CUY7riRkOl
fUWvRT7iEZpDruV8cccfMiZNzvRMnZSn/5L0nY6TBLk0gvZbBaCqDQeleJP3zPKxgyZCbzxithad
kQb21LppbY3JYIB3Eh/rHMTB9+iBV369EAyoNq8xH7OfzKYRrGfdsZqJXySxy17Db/s2P9xX/T5v
d3e+ZjhhPG7S0qLJtX5/EcOVXzhnb4NcB3ZdAZCstZnaUROfTqGWRfcpeqEfuEQozZqDd34N5evG
XMVTs3vmS4kV7AFR/51YtV4cTTUgT8RO3uN9/etDqjYUGYyMYT1f6pOJRXw00PJH5rSMlVmQLkSm
w9jEUqkmNxS3WUNiw7401Vzdzi6MmLW0nx1pe9dgnZWLmUVmIuZiZwVP4nqX31qVTRkBN3h7PrSI
1vNs01tmBk6F8YT+Jot43AX8djInEfTbzDexKXgrnWgQtxK27ldauy5/ndf2vDj3c2XHHMQAkATA
TQme3IcF62ePBD13dC1ljac7qq7SR7CMJDv1BTvq7LCbf3uBKFCz1EAsfnwv1MiWCB3r40U4WbsQ
icBcSKSZKhIgPzSPtx73mkNg+TjV/29RdfMG0zCvN16OUN3YyI4p5DokqmDqXExkLf1k3NT/qq4s
j5SCokmFz52Bx3rmdYww7FPotaMZGrQO16DAaq7ejrgd7nIV4+DBXQNLxZgi6I6SCVwj/81INUbP
mmWKc04NcEizfUUivmzjdLQdJXDYm8Mcg7Z7m4GkyDYibjhY4w5AJVboxkUJfyGzWg0FNFBRj994
Vtgch2gXsL79U8v55EX1wWNu2CljUO0qAynbnPikQI/9m/9kQqunksCMWUlFL3NESwg9hvWe+/QL
eDHPBCzNAWdI8ljN7u/DLSB0vRbypH3BAEBEIcrneDOD+g5nQPk4ljmvLipfFVtWdLafBPXSZTlI
T9Nevi9HCf1goZHtjcQcu/ImKrrFYLn0v+dUKX2bZI/97AzT9BERaEDFQbfw8uXbC8xW2xHDTfsq
I9wbL9RYvdtkt1xudSh/SzkazOPd945+qeBM5o8cCypLEZaf0jpGySM2WimFxZ16bES9dlnpppQC
KSyBqa2SEjI5t9jBci++Q3YwU4eh/aAdGzx7Ow5/hSf4eq6yrqvQsyAASx4wfdopLLTqmv/pnQbO
kdCZuQ1SHWMQYTW2hf1SkowlvacBDpsDnFt+vFfHkBuFc5jwdStsGzlKcDbG/2EfsmB/0iWIcEwx
KljEnyoW5gcA4zdCpOb5Pj8VSYoziV4FBLvK3y6K+q9v+LwMKQw7U2ibuRyCbkWbfrL4V2L4Twut
hFL8qQSqOQrPgZKdXh5fFuGPDVKEasL2BIn8quxCq2tsubkhzq1jBD0SZTgR3xKfYZUojJnY4b6R
0ureTfatBAFiysaG2kji6twEV7vAML2lp/HQQ8MdbjTDoXhmFlCDAxz5Ur/78kmZ0v9lJwom4Eyp
70dbUBtDhzigcHzxxM2rEu7pwQbjyLSqMh0trG1ByZOCy7koWMqCNcC805veh8eSthpdEHBLky+p
LgXTws/NhYq1ZzgFnKjCZoSv2CtocIO9vxic2ON6tvbtE6VBbSTqZYijOOjuO1qmj3Ss7f6Vxn9Z
h51FI6jsU0lvBPte1+pyvqTogu9z/3FeXViMsVSzq+38maCXoZ8vBkS9V6WLCwxXsyfh3P7cV4TQ
CP1B3zFmK9aoWxS2qQRhCMUIFNsPcMAwQ/yL9dVG31ElsQFakuVtj9BCBLxoMM9hEltEEeHN8pXu
C8UYGIykNRGUhGc39Jx7fSdWKt2CVD5FitR5xVqVpEwHtz1PGn3t9vqyIn+EQhGq/KpMzBvVJ7pE
i9OC5cgWH/NeWGlH352BYKVCOfep6cZruRUPDVmfr5OQJisf3lsQidNv5p7MUER8/ChWANQA/okg
PHHNtcehFb/IpiqdSAnpSoCCpW2N/Dyh+KakA8kmh1qft6SAMnXrfXflfkMR0ERMxFeab/PXRhd4
uryiMeEE7zFqC5BRQk4NM9j7HxNyTpYB3BBFp45tRr4J1F3lWFFr5DC0gmBOXQQM5ivf600mrrTx
R9DoujbN4gL4Tk8E9PapTzqMZg6kvI5LhguhTiKiriJPaaHyk37OBrumtcMiyGMTON7eqjXzc/pP
Qj96UqjqKWj2agaeLRvd66kMSB3+HpEDq1iKNVLdf6L/ClvrK5R78gYv8H64TRX5Wm4IDCmqBHJQ
aAqrMZwPUyt6m/lPdNEnNVYIWgjb652yo0C/rPVKmPVZ9I0ZZIKWAl3moxDRfNgEhB932AgDw5ng
qdlSqWFPNyl8UjP0WlQ2UlWlHcouk4G1KCUr1WMu949FTSnC+LE76EFBuz8xmUNEsZsslm39PtaP
ojaheed/c3EhB6VOcJ4SSwNJm2XnQ1uBkXxUgOZmBlu7xqXNrSO7QUXI45jrVemlp3AyEMH/U7CN
WItIfNdHtW+9TwuMMRI0nRSdqzbZJaYL8TOIpb4ky66zayf7tKkHyco26/RwrRuYuX2j7LbxekeV
RLpSdYjEuMkvru2b621WUZZJ/j0tDOQWrYMeCeF3/XDygsGzt3GylAq1dfJOHhkvQpE5fRIQNMej
UPToSLDhKraZFOmjz+Qs7Yb33eOOB8rYenV0qdnFEeVKhB+43T2zGbk3ewRbQSX+QJ/IVfMy6AZU
hPP46hRVP/+bRQAeq8xgwndh8L14D0nCmop0LTvu5SENnrqtfGjhlXGI+9LNpQcIU4muuE69pont
fVPWJHypgWff2uGzQm88JJYLboC6v2CmNHFS7RsFmEdAHM793npfs9jJEfUP+7oDqodxq3g0gURw
yiW9do0qoSvESeL3U1jCR6p2Glz0GabODAqJN0MCrjVfJ09yqKkqUrw41OnZwfiEw5q2bypPVaHq
iUeLl3xC1LCfL7iMiHkaTumGyjY6aZ5jB9kKkLTtoU2Jx+PoftlraAWuVgkBaDULBg8VkTgxILqi
orPQgavQMQmowfV0J43rnqMpBOHJbTPnP3CLG/FHOr1Dk2fuHPtaK5sNIiiKivtjfF0RTKaveyIC
rOkpEL80Djt94QLhs8g848R/+eOZuusTywpS4g8zyTqvfV4aXZ+xNDO+hoObFQBvHdtWV9srIgMK
u+q1l4HCOyhx9Q2pmInNObLi2cwQ/xLmZmM4moJmRdSlnf6Fgm0DqXYdwUkZD1zTYpH2+WmhKfg5
dWUvvb8NBakeUaoY4LO//gM/vVD3hCYGVKAi5XRbNjrvn0mVfZ7LCKJlBlyOy7kv/FxdUqzenvTb
9nZ5icGADuKLPbGOSWK43eTZRZ0nWqxgaffkUBxIKDHql+iEcS0R9wp9o/XBIjGGEuCnY+Wqf7eL
9GSLmK5UMalMgGXtW3rzqnZn2laOwYt8+PcvlMK3qIf4C5UhaJGfzK2r9qdWIFiSdwVNaohyiqsI
8GYlyVJDuc9R9hiHrLzfpdvIC05zDoHSEQIRZh0e4IP197wJt/a19+XDQeyCZLT7YgMO0qUStEml
i9e1Pja/FAXwksEUtKJtpdmnqhEc2m2ZODvv9rD0EdC9OIBxRjYa4z/qGf0I8JlGQXsPu+3mzTyb
J0TAzMqpNxDrjrNGxk6AMr8ai5DZt3fYREJcijLK0p6kx482Q9NFgpq0GAuMCnN8dm4PY28NIbJH
ScyTVIfyjMPMC9sYL/nRco00MbsXG3IpFrcP/G3HxIIeKCN7SSLCHYyAnhPVpXm0hQcy+z1qwqxD
Np3S8vsbAL8M5h+L39vq+pemEQrp0anhxn8oJ4s1JwozNkb1+1BZC2hvb8DmSLfbw5Jhf+Laqmqq
UMM3M7ZkREfxOvnjTeaEcennTA9iyj5NHzkIZJYwV+D8UyzVTXHjR/HE2RdM7V+v4xT7Qh15LO93
hc1l3rZgWH85gTQG69DS42w6eQdGRcSBeQONASL3O1aiMbfDrORo5njSbHE6fM+XOsO1NB+nzX/W
SNuwYeEIQJH0AFw16YBAgZM4ScQABNlp5lWWG/trJdNpbTjwpbGTN/CKXs/KftY4vPGKErnULktM
8jwp2JSISnDHSq+S4RxWQvPCeok0r2YV17JmctGQT99EAI6dFCdGtkgKZHK0TwbxE375Tct+93Jb
ZBxCJy1eR7MI3Xe/ucTsrOPcGPf9tZa9gGAJE+WXGpvfa9IeX04vcZdxavj5xx7wTDbZSQPNGIXD
NWNQrbdpLxnEkbopgexxVkEf5hXRpi+RwWzytLv0Tv37r36GAYnYGuh+W2PXX0iDOPpy3BCZtqMl
bCepL88pUoinvFSOUtTqsX4i6ANj4+v+GpLyKnBr0llRCJfSIaV3A201x9+mXuSLzZ7cHhOmtFe8
1Ec7UirbG6EC3+6kE1HAWxxFi8gPr+tBllQirx2FBjtSoBDvgiAIhUOG4XbWTEWwrMLWNLqO+XMA
CO1vyzTZcivQ7n0P2UDKMpy3vlm70AVMitz43304hbFSmyJ31SRN3sUEJ5Fd7KsuksJ0g/qj809y
QrcLNo/VpFTeHTkSlG4yKjDIe91nLyvMleluJulwJBW9mPSy2Tg+hevj1YpbPRWyQXMgKiPYtZbO
ISe8MwWaFf4agfxPuNnblYb67FG+lMWhS2KmJI/QLCqRzPsegAP1vnzMUi081itzZfloNxOqKJ5P
9IOcT7KQIwWTRaLO54txGn9H9okuckr0RUKkUHuA5JyN0UceJT1YFEdlQEPgujSeEQD16pJmsMMi
lPRo27IFTUANigkTM/jim8AgbqfXFavG0qn+JmOsxUdIrD0PWGkm6kqkudvPYPgaP3AdcGtvCyMk
YUcikEVKeNRvlUuzQefLuVvZ5/Whe9W/hNmrdC/B+cZT0LfxFYSyXk0AH1tJINqjVznm91oHO7rf
Lo5Dht/McT3yZX5C+mAbTAGIVGXfZcqKfMMI+KWg8w9FqaidQ3GC18fgvJT3JmazRh/3wfc6KUt5
CVXi1zTl0kxGph2J2YneIir3aOkWR7Ai3+D7uV/LoXXF2fJ8tLzfsihFEANhLuWtJ6OWXQd0ZtTR
P1vEzZ5rY/j+3TsACkDRqcXryDJby1WXd2hBxSZ4GAt+IY980evmtxJXXoGdT0e6stbzFPHMnN5B
41s//vWv1GGAJ/0vp44nivy9JvihyDLz8U7WenIBWp/XejMMVJ74vKsOuVm9DZIdWDpr0gSXqi+L
q0InaA2jW8HnIHbTe8Czit8m3O73gXqdwPFbAsOUCUmI0YqAKCgGJKGxBKZ9g4yq6jxscaCxkg25
AeI5ojs4PrM9zMkV6Zhg6rBcJFZHQnZUssT/1S17CjHnr2RNcutGD4Sq0ccWTvzJHIAtmHnOLDMR
mRLIHgHnoglBxzVmPSq7CLYk6MNhI53huMPIaC+o8WKunHZ84fdWADN06S+o1RiXUwhYzCWPFlaj
CIqvqSL4yKGziSBkSWLUM3ErSjK/vTZLaDfPsm8kw38ssaFEwtTRfent6qXQD3tqgSfsdlOHdjgE
EmUSncG9wD1xgjWi2Kr5jac23fk0yliKaMv7ZUBHWzO1FC4b35/Ol2FviVF6jAt3n+0LWT2PVEUk
hOWdmLzO0Ia3zN3gIDgYBFs31GzhPWZEXO0Wss5NzuTSr59uo9kO1sRzF9ztAVYMbvaLAih4R9nS
cEf7p9HweoKU/om4qRHGkdvGmcuqvmPIwhlF+eaWb6aGV2f8I2zbcrtMvTl7GtxNV0S/7LYepVzD
mTw7Z+W5iVCnPibMPm3xfWdGJSx/YoSN+HnHbTdEX0eqTQtRO3C06TNZl+UReGN7mpaKlHHMjkVL
B6AvmrlRSvEhhvS3Ay8Y/Jzz8SkXEAA4vDp/CGe4Pvc2fDT6WPf5XZHEzvcGSAjTt5AGXY+fhfyt
Eb9YUaJJgzKy1xukfsVM2zXQOEfv07BSdSS5oXz+e5CkWtRpPNEjQMUKTLVZPv7hs4DJBe+Sk/7F
2PfBJWIogsVi0KYajLZxHL8AoQ2clFiUVxGTXHy1OeGba+4yEVHREdsI1OUs9v2L94TMRBwBPVKB
2R1x4boPTXWSD96MTKGWluSNXpXuq1fdfyFJhVZESzFkL1Fa/CN/sxlj3ssJJ5PW1JQCmHb7Ekdl
1Dzet3cw/gih6Q76n5+HFe7w2Y7GTJdspGtZ56xNeaNZMsnwuXBd8bKW3bhAtABlqfQwxZHTJHye
lixcSuBZxz9lWXo3RvISZLUdIM+1uTRtnxiZZlrIX3QZgtcIauQPEmAZKbQ/sh4sbeteF2DlVFO5
cZtxaXlvHDJD57l/pvRPllW5XqfzuWjZ2VSqulgvtRewxXxYPQa5ajBFdsLsDSW7c6yy+i0lb8H9
LtKiyWzS1VPzhNYhNnaI5cU+r7ZCDPq2tCA+vj6kbzE6FBualyZ7uVwioCaw9CdhKDQG5gFuMlHT
j4991cOMBPJrcYTe9DC/nUPn+4TDxJgm3z7ekcYl/wL0z9Ieow/oLsBFlgCTDtATFhOWyyqR983t
4oT0FVpgwsa9ZMKoS1A23JS/ojCZykWvKvIVfNryCxzt1e7BwyXyqByPyEwYJfiaPuhT6Qr5wSEX
sNa/A18/B57uR/7dUAavUA2glVo8WXfIbGVFXA+6tRaWib/4OORn4t8T2EtSX/EOoOmMisq+6CXp
LMluGr4/9cA+30YcsQ+Oo5OdT0SsZ3F0tpDqnVqhaomqOZYMBqvUGUpnws3N083VNlhUcUH05PxJ
6v+yiLD9I7qMPyG4UkNNA8FYlmLvztrdrl698SkqBfsYs287iudJJwQ9CqhV9qutW5Oh8MTpl9fZ
u1zIsZzLT4oje4nh5AaT1Ci3k0Sd0hSN9u4nPIH90fsWTDshBrLokhWJ2Vc4ZYQwf1BxQRvMKvy/
BVB9aGVmx29II+aKEHTRos3zT8uUl0zA4yXM7p5e+CE9ITcWx2ptLJtYDd6VJ0hWMw6/Lfqv3NOu
dKDjeA6/bGvytbmkM66pfXwawcMoOAa32Ya+owFFwav9QIzXkSKwX/dE/gKQDR4w8I+Kyjo0UzgP
YBdAT2Tbq9iyjBDlUxa7lodHnxfTrqXy4ju4gdHvB5XS7O8yz4lfQ+WVikKWQoYZC+3GAoEpfQSg
AUYFPEOS5OwkTkfazvO8Adh+/81r645aJP/+QhbQaW2ZIyRMn/DAVQyFucFrOrFhIc3op3oL2aTQ
8FGKuXSezlhqeLNj8Orj8k+B1yap7XXAQlFzoxmOW7cnUn3T0jovr4+G4o0bGXLRvyv4ZSYoQGqO
p2JE1lFqkTQ4WnBu+Jjx1OTC0WlB9fS9IBDOK4muHgc5Tt6lOFpF4b6PB4sZ3Jo3stn/MUaqg7uc
u8JjSIaZ8n/lMSi7P1BLDxRqpwnguSZX6mW9zCNgyFH8mzI+XLhVLHq/xdIPIi19YjRPpPGbw5AQ
VgqGFCvi0QKELp0cHqvWmuXndCdS+vR/1W/sT6RxRCfwBL6OGPkNdxAUuvF15yulxdC14p++8AIO
WSUMwCq5G2c0Y8Pp8gtzyPGmRYtHJLxLscv8LcNszMKs7gDQ//PQlgbBYQ7ScRplTdZyWEtBrZdJ
HUEvYwQp/KGtX77qd7X8ckRX6+oWo10eJBtd+zSguLru4NvssC2nKPcFV3rBNsjuAZBZXrOhgB0I
tnqNpXNmcwuDimj7rCIVl9X2fVGOfsAXx4W9FxxGQ6oul6vzTrE54JXG7NQn4YYaX97eLcou1pUx
GrORDKDeEF+7w2NmrAIHZiGQF7/rmLEf1QgF9ptsFWO2tOTnEc45kAd163jz9JN9pgtEyQQkI1sg
YdxoZRuhJWfP2BGfNesTTkX8E7URbpI7CmpVh+SKp6zdYGbtuZFT+MeprbxCw1V1fJE7Wodv7pwH
byy8wpo6QguH7y+X9zdj5jN3rhNXODqL6bd7MZHi5iesdplXHoarTIfgsGMeZ9CrdzcwwV6xgsUl
XDxTtitBNtw4TDYoicD6heONFN4j4h7tjn7aGvg4grZOt1Lzl4rUIeUMeMZ+3WdKOEN2fyM0D89U
BpbElp1Dj4Y4VqJ7xX025TgAJQpHRBjxBJpz6RPfLBtTKG2b8pfkFG25mF5alTWqRjbBerQ48jpr
NS9f/Y+drl7QdIiS0n65t03P0f1wLhJtVm2VWhx9JM4rvkE+JrkG97h4/5+1xmqEdjwzL9P8MlEq
ZnIQ5a0ypW4nPehrBAvj1uJIUZpwUZv5BP6rCQXrCBUSWZcRYVDMn9Bhl2Pr6waT796+cefFtDdH
EzlpSGlz9SWWh/E2AikbtkEp3naudqpPFaSJpVaAvWmWgtEouW29mE+DGb+GE0gQzpUN12g2QNQO
puj4gCmuqxaQclTTbEFfa6lxi+pOWQDKkhx5A8S7enL5BgHXx1GhOpGLLXVkBX4GJ9AkEatDVCG5
AbQCCUb6mcMGlbyiOtN0PeEHfHrz1yO4up/D41sEJzfaZnNEa6RrCmnz/+XB2s7clPl3Bl5NjX7D
lv3+q9lZon7C0vBzzVkTd7lLiKeKPHtHarDtqsV6PQYbyrEFIyqQO1LTeoLMsoyx2lO7KgvPrXIe
dTuSf7TWocw+6ph9p9lvPJXvXRnRF1Wml3GnxYd9AN7xe5VXuJ3RzbX3c1+sLWnsBPWWjo3VSRku
xQrxsi1IbmUJcIag9VMdcw1Vh4BV6DpraXi22bJB6197Z9kKGLB6/423Vmh84c1LiTLQHXwIEwvJ
wRoOmZXkxsxna3sNE+swOf3x1S+lb0qRAEa4UpN8Vj37ofTT7fNrlYV8+6yNMGEuRRGgsOle08Tw
5Uy05L3gdjWWikC99bzv4gZrYn/0edATXxVlRcfMQIZB6pn2ZYWiaagKDsqu2USZ5FgQLHKjgTHw
dwz15idHGcFYz4CHwxL521/5AZw8OZyDb+Bq9yCD0ZnHgSHS8byNJqV44iGJV3aiRaQqYSC8VrzE
9XbB1o12DNfJOMX3IaPmzED2EjIL3njrMQ0dHDtAoKMXpgydKOMzHZjVO7Bq7MbCT3Hq6senDQnt
zrN+sWk/NpGlwBL6xczmJY3BvOzqoXfOakzNyFnFaOriN4sE95TPT8njwtDuA0Poi/mlmgB7HMQ8
+FAE8yp7ww9p43dHkLQnV/GGM4Rq/ZZ05oAK3NMiWpC3Vaq+CffWWf+n9z9cZ93vpmk7iZ6JgxHP
rztn2Fb5AvwUPy+Lq9lle0/cvZnHAC9noD8NAVjDxfFQI3UVrI4J3Cv+xGlW1x3d7sNlWKzDcdf6
hxMlzKVY6mrGY4aXH/eK73l+bfMauakgHX0HgTxEzjaxaQVZGFZ+5ouN13W4YCongELavXlVZhG7
C0X0FoMgZM1Wd9DyZMpt/iRfTG4vs/M0oLNX/C7KNEMhLoOILJRZcrs7Aceof1WocMNzHW+l2Xr+
iNaIAk6o2JruC/2eKHctbciq5YX2/E4eja+wOZs8B6zZBCElITf448t+G549kawlf8e1PHmQrQlO
VfxYpiiWZBbKGOeuj/TBeuXatgfLu1Ie0tjnaVKlxqDG4ccUtedJGTLO1I0+RN59NcwMJp9E01SE
x3Fweh938PwZsDAiHiI841FY14cLelSVr9mJefI/QHD9+3dQW3jwLZnH1l61rgbGXQ9GlbBMKHJi
N/4BAvVKYDhWaIwEcC5o+ALvuf4765TCWJF406QEJHQIFsS2ErH3NTXk76qTMJJscZmdPUKfWefR
NPVaTpBgJYliZ4k8IBq1G3HohJ2vqEJQIPC606/dL0oREafc17IH8OxRnds+CFzH1LS6oo2OSvLu
f28fzOBc1yiopTRnhKRsmFO2VPfrgbBGY18mLcNSnSwPcMDh7J12Q7+ajrZFHYzwGSQ+f3kNWmYv
indX+X6pQ08j0D8s1ZP+Mz+Hsr9EIKDi6gSlQmwmef2XBdfzRUfIgs4n5ex/CctTpBeBVAAqZ3Al
qBFAOaDVoA6UQkNdz1oigKOWfepMOEJJqQ0BM/VC7iPWQ2vAE4mpKqkrc10owra8R9UxpOpiMT7z
ohJl6cb+luDuE8b1sbRgRC5hR2GnVvGfUQeE4TPYhkqsnLPe3FmRO9BTibtw1BHkcCbehc6GUZ0G
D6gGmj2gwtwR8C2ptp+uq5D63ByhLKeo67P+0Jl0FL/Vr5Nzw5JuQqcksO3szVqI/aeA3VW/BYhb
92NgvcJWu0j1oj9IGgtQxUACABc4OaumGDxgqNB+qlBViEpnQXF755QNbCLzCBtSYXoWihJWRz+L
G3LLPd5HN8zJrKIME1ErglQ5y3HBsWtGDdNrFI6QK4WYGrJt9VZEF4H4iI+24yruPSJ8Prx3Wjfx
4qwWlOvuiYZfDtGIqP45ilK25IvU6OXknxMnMZ0JWVeVpTnFAfpOp6xFoldEt1kOlrog8nvFXKF1
XX+sIZQ81GRKFzntGl/onOEEmrdQSn7hyJTr3m8dtASNT8Jm6UbyTg749kWXfR7+r3fPd5i+wbBk
vkEoX+6d88Oj/8JCiMvqlilH/TdpI4ODLRqiE8HMUudz5LqJg1/esExqc2BObsJQC7lviM/LzfRa
2Bvo/lBmYNFgU7r33ddJK9iEhJrvczuDQk0f34jyD7I5YXTNSE3cNqGFBWDH8bypHXQ0igXQfqY4
GHZoLdHg1VaHb3FhhIVgqovYz4uKiAAAdTs8GqodEip3ofCglVvmvYi/RoUGd1LzHECx6naftA/1
SgqK8MmXmaaKIhdQ2MFhNuGe6Bq15R0sg6nRI+XyDUfYGKrETsnBKSU1gTY3bjfHOnBoGlXLf95E
ayO72r1Y9H+5moG97naUMQq6iily6LEipeBGWkRLqVHR+oe45L2qq16e5Ha/PKznwicQnFDzK/kt
UEwiWfmOA/KCWv4k31GKE8KK0rdvTZCAAAWcp+SssvhYpY0pwLRWV7B5FuEziJDsabHiPwC3JSOL
MWPPhS8WYqrnFxL7okJQjIcxttutF0Z1dkMsJ5Sq24QH7Ps/SC+rgtDjQaCj7dIAFpw3pFFH3R+y
XBKDEGJzIwuielcKOywVlLLaX2i/NPF2nhgd//THMKEMqYiCmrfCqR6IaFhIfMDivKuAE1YFBG70
+WEOTGa59zaaIRV4H4Hn6UHbehyfOgOjFrORcIdRHUAEZSTjyVAl2Mt/EyaRfLSF7x8OokgZthnL
FCwzgWKQ/JsUXO7UV3rXEqedFySmWICSCVow+zn7ydYLIuqdOoHUlHqC9y3OYLDYrQpTBwfGqfMc
SmcNSyJwbQ77r2Ke9tnUxHPQv48rhRcA9+QiCUZsowTXpK0qTpg37EFNuerDSTyUNXKOngrT94jk
Opwq8NVwbUfXmcKjDO7ljBd+c7aQMvburRGXCNGT7h0R9PPzxB2IpQVpx4cA/aI3QQloRjwpTq2g
sO9dmQ4NCsxt4LcYRxsrXtYuZSZdipgJA04Oan+rTTEWTmHYp7VGzQdFR4Vt/COj0ZyEGKbs7ga4
VOYNpri/2ud7bSRcoM8Zpc6Af2cSPGx2AhS4E85Il9W7CsM9Meb+UmyzYWrMSoUMZQnUrqGt36rl
sDHBhO2xyPT/OXJAoM0mSz1qI54ghF0Cpell2XMMTvvil3D33MAcX2Hb67QXgAVOamiQt1Vil74V
4orkfp0tnsoSSAajc+LUZWvY4TnKsbPsd+faAWFK129I/ew7DQ+edy0gG9cqz0b1JIfmZBYQj495
t8NUL+/EbuA29V9G1uAKHspZ/LjopQXI8vRluqa8Wk37wmTodeLlt38PwOFKUDw0Sb1fAvDqi3Pv
cPJKEsyK07RyOKRjoU274GWPgzyrMRVFDvV5DxeiLs9b9z1fT+JrCVCRF0P5R6ZSKF2q0jlNAUF0
OOJyjbgzfiFeAIRw6Y/07pmY59127KDDpFFBXzMaFkqRYPKb7Yesus5dT5sekFGBcw5EZh5t5hQz
jmqEt5a+uC33U4dl2M6cCLT8KkVWM6ghuVwDHirqXLbi2jZkNoCGEY/Zk8Mp3xKGh0l275PfceqK
Ul0xqDYRV+EYxLQLV5la5TlAeov7E3gGC2XPh3y4S+txV9LyGP5eE45idOE5bG2QFHUxCzfOnzws
eNyqr5IcTGvEY550wzgNCmfSK1TfsDh4ONQQfJmVMDKpPFXPiXMXSGLX2g2XC0nH8hgq+FGyVPz9
siRruLYUA460M69P8GSegMFpVxUNwyK8bSxEpRHykofG8gWGS1EeZCxnpbavh57sa8xOkUiPvT8h
BdpR+mNoMIkyFmTx2BmmOM4c7y0vBljVZMfXD/aOntGJ58ErsSKywzboJFnJOPaV8Af7XyvpH9pA
i0OQ2ACnVgK29Lonv3aAg2HqKbjU9xP0mrVCLRh82yxHb4QhIINT/4mKvQXc9imrPQTKDzmEX/Sz
mAtz4ivEt/wlMbJoZYFOMT+UVHlNbNSM2IkRi6f3N1zFw5zVwCdWvzg0Z6c1k1LRY8NQDwnSHL8k
9bS7YNPNGpeDgMAK001E/nSq5TkJv6ZCVgyqhwp/StIs6TpGXrrLMO+EDwpYAxpgNzJQQQhh6fAj
4u76Egjjh0hi3mCwP7WtvuF9jr7nEnfuoWc6mvEXMRJaDUtebQuXq6eTxJgYixt5eQ7jGWiOGKXj
Q41H1ouvltr05EhVQjffsp1o5gsozYqL5htzpS80pVziyrPoLhe9xQBLG+O4+iwryIlCLE8t2oyL
QQeV9ScP0ENWbnuj/l3AxggPEeq+6KIG1sZzzcLkJ0M3KBuyPHGk0bz2QB6s0ffq9dwvFDMqP2cy
UE22ei4o8kuOQ/I0PoZ660Z46A7w7gL/TrxdPdfEHlP9EbNKYLyfhsT6ogrGAOtm727bd7s+NBxh
qdVdfI9Rq+hMoRHlPVn65+sn4lXv/2ZlvpwSy94ucFTrAFvXxSiBEXoS5LR4Eq15Cy53pk44/Ih5
z2EpfW684K8dxzeJVs5zMwuXZxxXwbPgrG/BqjHilbjBMkMpbZ8UZm88aK9SqV8GiaosfzAZZHrP
wbGmlc/Tod6q58Irfy8/Zk2KMS6nhdeEJCPxIhzFQum/IifEVcgFsD6qSznuvGbQvHFidlAcKYxb
5tLr/hg2NhxaKwqLBQHS0JZ9htPpO/agRt6yK6OZBAV8Kbw4I+O2jmmcFR9vlaQmIH65X8FYNcpb
w+eLJBLANLIGrrKI45gEpaEmDFv3aBHCCpbPVGE/6GpqokLNpqVSCFskNzUOfEJty81bvFi6T3Bz
JTqdl3xCWXVVA/2U0iAd/bSzQoTY8B3hcKdpj1Uep1GrdlRjOYjB+xv0n/u2LCCJjq+9Fye1m9Ul
ISyy5SO78nBrufN4xy3KOkCSarc6QqjWPA04T5xrH+iomgCv9NKfuw+opPiPtdMSEbZ6U4C4u2sn
FufQ4e6xLH6VjDTjvrO8X3RZMV3DbA1+WZ3IxYzi0+pCES8Omwo0fkrHDaBapbPhrOUOpLZ1BCs7
n1A4lMcwv2v8xBCQKqyHaJz3BeW0L6P6BKWuwJXxLtMtr6fHqx47onC/f9ic4RBFdCsmb/7DgC3Z
LNiy3V8Lw/1Fk/JYSadjAKVW/kgMAO2J/lL1HFXilii7bPIls5tuFBCgpmat5wX73n65dtmp/7bn
nbNeragfy7f2JSRCg8ma2/K8HcIRWfrypzQJWWapAqmhpKUD6bNYn1SJGEjVY0UPbkdDRJirdeTX
pBYz8LK4zgOpCQbDwsI1ooQXZfry1bJlNrbBVnG6ABm9SPCrHCEbE3ckxbNYl3y/WnctA3HSG/tX
A0YdDN7Csn4aKHZ+QdEIDi2y0eLIvSyWi1iU8feCvDoczaVFwm7gGNl4afYNKMjlDQ0aezTzChPS
FHCpI2t6BLT4njeZp6Kh4vZXhHsDHq2vXMGR0CnYCpOIEQDAd+KMuAu/gEcNJ78bh2GX3+zOFwzD
qlHWiboGKF+FWCiPevsCNg+uVWAkL/+X1X7UiYL/WER51elbWypppn6lp40UsKOtAanzQod2mN8T
ZASbiRglQVRNf3xdcfgKkhrBO+uZ1Jz9V8t69Iv/l2+5FJSHOVtQ0lU0Te47SvblnlFniEGpB50c
vCmJFz/N5L0we2MaVy3BE214a//TnK8GMLWpDqF9TQ7GBNi4UfktyBIbtOHipRkP2XHidKdNE3gv
/ee6uT0GlJf/vJ6hwOvDEm6Rr0Mmdq2dCPiiJJGpuqy+tWhso4cqElVggvokplFEnBUYllctL4E2
mW9lNetA95zKEmOvgMpszGbJZl5cebzn5EgMtW9tfXFqDY/WeNDHqtoCC8jVvhCFkAwJlMBSvpPC
HPwn4gHyILUa4u0LP9S6jerfMxR9LShXcQ6TcEnbBnXNHYogSq7TyJawlr5ZyqlHxhEa7LOq39A/
/sE4Y5OIzLVUcDQw/2LIYkj8erfnEwRCECLBwUooE8Nf9hqm8TjROIclQfS18JqRnjivSVPzSaUj
4faBLE6gMGE5gp5nBf7sC2H+dL37ih196hrEu8N7rvACKiX3lWXFJIVcyO2FDaSLbABse1jIIwRt
FcOSW8OvuHeKC/JFBoeQLmOf2qbNLUFSlnO0Wp0YDJxaJM7R+z4ocgM9GhBXmG+cCIcfpwqD9T1E
KwQSzu07S11KCy2BKeN9mlg3Kbw2rIj2krRaEksEOIvQsvz0Kuy0TEzz7FEA2xH5vk4CnA4n+VYS
oLW9J286ntxWGCFg3vGvbNK95J83IE1ElawkkCheNknYCU4dk8k5u77ELIH8yD2nK3RQMmpGng0L
6VJcwXtT8LddyM7r2nEQZ49KqfRjSA56XqIUfUq7gSiof2INkaidCyCpowY/vUREvVRWhFzAZqf0
TVQbmKrXsI02hAksdLGIVfMbJrNX5Us82x0qh5zHRrizUJBps8Vpd2P6KQjTvCCwwUeUMAmEacFW
CorFHls+/gckMYAhceoj9SiY9bf2cIoK40oZ7+L9ZbdJjDqDvFDuo8dNWgsQRczL3SN74Sdz3zwe
2rIeOt46dA9e6Qym+qTvwoguSK3tOD6/g7W5zT5BJBuLE9f68v8GFX+mP59h4OL72uhvQ5nMsmYf
DWPHi4rMmDXXLqkEfqxgO15uoa0DksqbQh2UVGd5g0BYHdszxggwW8PpOHX9JSpuxegeuWGDtIa3
sdXbYjwVPrP+KIWRMJsvCkTrbT1iy5FMYcyTBQSBgmhH5b3reqYAWh6OMxnmM8ZhXWFWUi7+pgOh
aKqFAN1sF7uzywIs7IZFCqiF42DHwyWxtQdwNb0ahdzALTplxHyeZpl2oea81pk9y8fbzIOgVwo7
laS0zdphJZ27RmyThluetX+P9F47XU0azMaSnSt1lJ3eOWQuJdqIQCzJwsvxgxRT/3qqM8ka4iZJ
2keSfMgv3aaDEIQsWH94Jz8ndau+NywKkCdVZJamrFugVdOeQS8pTmcWpg2WUBhHs81Wb2/mRBFv
p4+i6D4v52IdEvQVwGHXyIGaw+zjkmWfmtg/kSIIBfVu5ZQrnZAkQOWZJtrJfBCkmHJ+Gl9rfU1v
7DCRVpaoifjdOVy0M3GO9Hw4cs9BPJebgGASwlrxWSfky/iP5QTg6aspRys8n/nEBrtcysJrL4Ys
jnIjRyelbV8RaTSOYmkqiX0ONZ2kJZQyzpYv7grNULHpjxrHPoHXd9mXaGAmEK5Oh7tkDuWnG/NF
gnnFzjmAwa3nu5URkStIlGH5b5CnqsWCcsj5OzD8yrxjP+J8rsFxeaqhxDBRex6NQVPsnLgkfuIn
/mp2T9DfResHQcj4j0lImXvB6YhSAywpUOqVEbIPt8ZCinUBYafgMil581YEcIyb04SoPb4Wg6jS
5NQeY2Lcb5RXEvIHTEg2tfl5JWiWZyf7zKqTlWB+LjRlpyO0Gb/BUjnJq9ZTkaNjGwvnIIYxY9Ec
jEDnrx+2daazZifADLsaDP+/G6GKDbQ24WIrPNFICzaikrgsIAkGyOFcVQUmatp+qTzEB1oWuqZU
mBInsyWA4a+QcY0xxoSwYIu+RkArNgyuX2GpD5K4KNFkS/6vX5yFJLEMD/3EGGYbUPyO/abeEvE/
CCf47qxoAywrECR0iC+Zg85o1v1tegsiuRpzEhcattDPNhFjrogwatfxQpxlpy4esbtFRO4d03xx
R89c46fGV9I8u33O+2znDrMpP8UKEEWosDBeIFVqPg0ZsZvr08hCrHSYdiyFLAb2BalYoIoO0xlE
inzpdb3pPNSvBCgW2meHhUSeTs+R4/LTrq1/qojtFo9nOVZ6yDQm0jRZnxzvSMgVCcBg/uHRcHd8
P8waBIzF1pKr50eSPejsX4Csldi16f5PlFnVxJKEjuJNOHOauywuDZbHbvp6v/+kVPHJUwb1oKgB
sMDITR7vD7EgSGdrMdyYBPbp03/UTQHrOC9oa6OAXtFvhnuPkJ6Rh62uTM6Hj0kx48oM1nNMx7y8
86ic1U5zmqCwkXiCbIkodeho+WSaPzo1Jfly+vzWfTDgc2Ctu4+SAT6R0w3cvDRrg5uUmGxCcLrd
OsLcRLH2L1aWwny0A7cpLmNA4T5/sozO7nAUzRkIj5Eo2vu3GrJZZQDLHmfTos8s7VhxQ7QO8g8V
BQ2MbEDNVrSNV9gGUpVdo9VD4flj6wLDerjB4n4EaKvKaQqk8bQf4eQlSSw686VJJtgWGC8zdk5J
ppfok0WxeA51vWp759gzUa76M9PhTgGc4nHA3DetGIEkG0uu5EubIlbx0J2fARym2sKpn/01BDk7
rnuN+uiHNyopKMorJnT+jQpSQt7wLHvgbVb46sHJA0l+Dp7JF5KRJlVT9lQFb6WjE2L8SQSciNGQ
YISv78I9zDQxaOprwvO+k5ycYMmDQsQuipjRC2vITViL2dELWsbjN/KLwHuvy9L7SiKVrmAXbuAK
9qdtowAhbGqGNzL2c9wWCWDhdft8bTOcm6G3TPGbG64GfDwDmQ7EXJ2zwdKx9P6iEQXzhGVZfHAU
9JD8Ed+AG8WqQEqBodO+1qNw5XwXRGuV9ODthePagvSV/qih/+4cUSOZ+Jw3kXgBtIZSk/+0D+iL
xrxdElIpfK1xQy0faWpKhRW0LWn1v3oQhQYPGEQSgYapZ2gGLKjgdD6ayvouyZ7eWqftHYn39SGU
Gdd+Uu5De/7MlkO+ZI/p/x3A56H4tGtRv+cf7O1Ph82wzMfA7xZWXIeidgfF5C1nYSmhPPfNG2II
3rzm7crm1t1nLy2Wl1C86geNpz7nthnZLU7EUiDwdbsxiD/KPHhbZ++BMSSCJ6+XCFPVcbMtpXah
R94bPhwX6SoLN9kcdILTQQEQHFfMWp9giD48IK5joOmCQVLufOYKbc2iux09r+W/XRWAHY32KJOn
+imHyqXcXCkaxwaG2W6HEiek+FiHBQEw02701bwSY6IG27d7Wx0XiZovVCnu815ZWiUxtpgIcxjd
eFlfTnsgNZssVejNomTZ2/akAyPsYvNJq/lVLNWEyANRjNIRp42FsLH0rmkCgg2q/SHQR0A5rQrp
3dG+GDDhao/p3cbQxHDyeMNJSnahactb8gUvgFZIi3rth15EZ/3klFM0H7nWX/cqeDh4PChWwb8r
1iunY0aYzIiGErC3ICTorYSYQbEfqIGsEVI3xEYPabq8BRuhNkuLvtsdLRjcXmVctZYeDs3eeY40
gOsH7/OAJmkme6wCXAhpRurcNFYt7QTFY14+bl42sGGfA+7zIol5NyztDhsrek1zTKtbsI1WiVJF
m2nok56X/qKY4du5KqboNj8sQ2tS9KdTVJ0BjzhFSs6GZF1uylxXftrlOEpHY3CzYnbcgXZ/0QBq
1ztzE/GrTtCT/32XyQheVJgaOJfkcWWzCW9tvPSd1zoZX3mSkcPiARnfJBEDaDU+12K3dF5JEnbf
c4/sNc4y3g5nnjcvxC2vBOQCcsxGvOR7cRQANP/aO5fUwjesdbaaog/PRsKg/fPBhL0Q/+4HW1NA
omUmZlsPar5gJBXXey1BozAb87b2tBXFgeClg6nYToimKgnJjFZCwV+1JtQroBpEv7HUA81DHXpi
qOT8i3Rr6CkZ4vzp8Q62JhGG1mMFRq6vFbYsK9fyMseE4vAoH855dOpdkstqEHUdafkWeSSq/Efo
IUsc2jBkhvhIhQCHiHM1K6+2obzetdN9p2xR6CNwtYndPGKIhMagsgJsq/Ij2SRrofv26rf6nqnp
g3bKdNdi85MD2k/hcAum9NhG7EDg8pUqqHd4E3AVf3LvDaozC9CC0wh2AFo0SHKF5De2WQKnJyj8
qRaoG3U/i5gb3PuLq0DJ0s+CenvqdsiGFf/WZEdvlhxG3UjAOdb8QWJ77lbYk3DoB98MChDh+eLx
l3Tkq6BI3MxgdweN6X7f6IRmKGeNCL2bRORyOmXsP9yc1e4n8Q3GCs+pn9JcYPmmmpfu+VnA1YVR
3hlerMJBrt7clNhwKiAHilWpE+mkCl8+UQ5q8+IOTfaY56hqW0kCqy8Xrjg4Oi2r7vfii5C070fA
Cj8o9BPg4kj8QqEQQNkwDjapBAeNDpyeOozSRg+pfjNZ4KrnZ8UYzpsFnp2r+0iakTYQMRBqhBxs
YI/TKgzFW1gknfMRoQ1mxGfOqL2m2sK2BdHgbAntVJJs65VlRtgrc6zWKESFqZSA/2U24x3zg+w1
AdOs8vxvYAWTSATeLWNC+ckdYXRJyTPdjTtTmhnq4A42VIPbWv6nDq78VpryDHiVSJDFlO1SfOpK
IIHA1kph1ZDbJmIMiDal2evpMgVpiro0p3ipShi3b4BnB28F8VLFynE86FvdeCwueZJbb6AlTqOK
ZnvH+wjsWbwbTLGvlOCJjtxpQ4hYhY+pYh5NSbKW2S+xNf8+6ik7V25S39AQ5maayjmeTH7yw0SE
czihUUwp96/92pDQsHIQ20k8mt3gDe9gpYymCXXvzeK3zVCDUjHwvZd4ZfbLOAMnIn/+vc+xXqRc
iT8g0DC5F9fM9ezmD6GpOl/j+zEpjQsOPZTcA+4LxeX240LStYd4KqFfTD8T2ooOYCF4yYOLXrSm
Gsm3vFPwguHQCcpMOWcUzQKjwPH8dtrMTaRd7CcdRvslK4rYSOIPDelCm3XVzFdl7uMvSdQfhr8o
Dc6Q4CHlYisIFdRcK66HG+Ngqr77KaEpiwS+sCwPCA8RbCbOHd95Z2RCn4vx+rHBl1/3dBbJSMOt
fgyHd0ukI+JMnuvIwZWdYnvhb260QjwCQ1IX6EfMVYQDRQUnQeNXQ5jpj9T10odGQKv+M4hSeXJh
1R1TgTTA7hgBxyoLxlR4Jc90CfT5rmPVPqcn2RK8rJlAlTOnBufPN3WucNIypFRPkFtIu0CoCToa
9NElIVjm8g1SjWvqxfwLDuj3Wa3XW6w5vPrrxPqNZelMZGsh44vJ50vBB+iDoNI3VH7SzuvUJTJV
BFneUcwAWReVV/U3UPLBnUprtRKEd7MFm1annG23PBioeFRazYZYNvTJJTnc4KbaJdWXZI6/KlPL
jJhNhlq2XPbzG5pt7703pPZKdD99XfLXNvookvIb0u3dFHVfz2O/C8tIR7yncVYcRelPXkIvWnpV
y2OXlyczSAr74k7YXsnpMGaYc+2OF40vqn1kBWj7hMn1Wl9SBIkp01cA3SLBjG7Pkj26t2H3pgTE
Pp71CJXoCmDne29eruu0A6SVJcfe8dFJkYeuiH4HdegiAFVeCi+pnRsa3bCSooW8nzoT0vLKyHTP
OnMidrQPOf5TLC9SJ/zPb3q09EBXXQfLUSJXDvLfjL7lgDUklpFA5nvBK4yfUhUxhvRmHTS82UHE
Xy97aDhgQ0shs5s2qnKX1ODolcqiANl0BFxMyLnUNG8qrP3pQzXAutP+EPpt0xIzbRzltSbD+J/x
yrhJmkyHxshZvj1QeoywoV/1v8guAiT/zs5hdtCJ44BXG44k6ExqcFRt4E8Nz1bF7GdH3bZvS5v1
SP3H1CDpy7OUJBlBr7lOaXhQo7Oux4SP1tNlyDXSxyq6A9T2PYPWgB69y+3WuPcsh1s4z1QN+7qE
pXcuBjYhPxkOhw+vAUi2rC4m02jllEWcGUKlTLc/Tw21f6tuIdK0xPvV0uvfJtUThLa/ti9fMfmk
CU0kc8fi5/A0lsZ7Jcv6rCax5Cfzwr0D1ykBtSBtptBh+SvNm3JGq9iZfu84V0DapiCvlaRY6Pqx
wjW86rG8WsSyY6Fdy6+SjwVExp9BA8PejjPX7K9XLDsKgvPTNzOxbJiL6mnfDv+ewVpxOXANC2Ye
uv88svNjzFqnfxS5v78tjwCfE9O1Ca9u9/w8b4btnpy6yWrooX5fZuVxXf1/pMwx2ItV5ADSowC0
OptyGh1ENwrX1jnDc4sWyEIVd67i6ZOB5O9Gfs9boAQ+stZzIegXkZClC6eCOeb5F0EdChfUjo6b
uJpoT1o008AHYErh1MQHfmdNMsRKUZ+paTEWymMlG19aWR60CQOh8X7rRCNjuMAHdDvWZ1hRY6tU
kqqtCGZEmDTMgf0wJYgGMM7hYCs1TjxCVrvPxpsiR7NJbYcb2bSt5i3syF1ZE8HKdwgjn+j0oLhr
ebsW2aMi9QN7nWBZrC+Ma+xIES/RwwIH8kePZ3H9vH6g0fVZa9rHl+6sKtLh4zspr8bHQD7YB9xu
LJqR2Qj/Gh3ai8d21v8+9yDXujXaBct+KiEe/q8Ts+WOf9Rlrpn1olc89cS1LUtQLXW+ids7CRCq
KD3H8xuQSxUE//TuHS6Hmvcs42xsOvsF+NmWbt35DLiEjQGmaPD4lDT7061c64+kONJty6AA3z32
yaISQpIQ8mHH6eO5AoJYkwSZ14BuIdk0hYgl8PWdwW5VYwecAXl3BeGOFkPFD4+EQAlwwC1n07cB
RKL56dfVROPLI8gEv3UPhvpxhd0HhovCKjUqRdI0BpoVgS+2qoJr5PNFGhhGXR6VdFGz2/Vr9PEK
hyyaT8R9u6vi16fD9y1wLzqSwbuYhvJAKdDIvrSShjzqHAjzvc95SpxOE+LKp1URkC25EIe9yIad
dcfxc5ACxfQ6HDYoV1dr9OJNN7G3EF8n35rYWlorLfGhyz6e6Nr/EBPu1CnJ8IdVZVDwshXsM+bf
ch4mqNHkISUeddtl8NXnFDdJmR9UvseSYBgKsz9dhxfRhFUgoNY0RDgUbqvK7ffHe5a3QR6NGim1
NRvH3w7otOmKIvktYDwpQbecyU6VmAmG1ozRpRWOyKSK3FDToIXnnAEneoH0WtSA1fqfgVgrIYeN
hCVvhmHFB+BB0TvLDRNXvh86bXWMJObxS4cp482aLVnl8Ug4TcSpKF/kSmjSKRZPJfugnJX8fsaY
MMZANMasEoAwUAGt0M+LN8SkienZXOnoNZdbjCWtfhF657ysictnIsmdVvGmSqQtKAqboqy5nckX
AmK23ic8sFOvHbFBKtubkMFkYeCpfAd/Jvne6m/8taTqT9IDRqHE/fgL9KMXefTHYuPBaPUaLSGR
zDzyZl/sWlhTUXMpTiwNDSSIOFEbJaQ4R+NCsBKTTzcfd4iWPFc+aqNVT5VxwkYO3F2Zd8CFk+4Y
HiE5QhTXe4E8S/FQfQc/1Rej1KTwvcZzFaj/v8waUOOObfSUX3kZCjIdW4OJHi+3/0u5ZpfVPH4i
c0vD/cMenO3LRs+Uoo0wwfBulJadTJomxF7H/E93c+iFrk2lJxBNvL8/OktwrsarfQtXhfmioOfe
dEs7ke9V6f7GeaJAM2Tv2xVVLHDjsAeFGNI3N+Dpc1ac6G89mwCEgFtqxJc3pYQbJopOnHskCvf7
nE85kixR8BxGIOZBI0zHWm+pBxCdIgmjJdogGhruy1dKb5SJUrh9v5QZysj5shEHvlO/Ao+4ZYL5
skipj3+ozT7tAz18jQ4ZDoEF9Cy3uvC1qhswET+2q2H9xCq1XVasht/RK0qW0WFtHbGsr17NTV3o
Biz0urR4hlUlsEHcdrKQe85Ug2W0BV/7ClZQdpjrFpXkPnoRgo7No8NkX+kEJSdS0antaoMFiHpP
ylNydCYTvqtQw/X/bUPFtR/3c7QDtIZNB+/uw2oNvdCIDp/Vs86J4LzPFBZs80NSjT4SjvD3m8EZ
Q2PMCjidUWzhXdwaITNLLUKxRrMrENh6oqdwrQuih2iRoSX4Ua4KNdh13JRcMTgScdYu6S0/Vh73
1SWEQIOaG0oNDvdGbVusWL6NLi+X9QetCVRLA1VGq1LBRgOawTMtdClUsS9c2KqXxtCLkOvIEBit
ItrFWDgjK/9dBDAKZVXTZESU0mXvO+Ro6pTWk2kmCvaEKO5e0ATU/h0QR0r64ooqDbTKkUaHSCRe
RG1N+xhxj3LefY5A2/tKbBAM2m9DAMZK6HO14kb4grdfM5ALKVg/9Q+qwurpJe/Lw/xlSNlMk0Tl
Z1U8EqKM06QNv4QviFXcsJkXcCKIDVZw6JBJzFD8UoMrFAhrannnZpglXizxeCvINxNNr39IHQmM
WXfvKaVUyb9V26H9UfzkcmVXraqrPeXoqvKrc7+cx+qAwgEpCObRE8+HG5T5G3LkzIcW7Fln25gW
MD4WOL0heYOnczRf7VPnu5eQVMrC/IqM2oWj9xzJe/yj785PiDdQI/+3tZLlZzwdh/fWwiKe6ng3
XoCg9ys3vdH4b2EoXSL25bn98dePpw39rw5kaG0Q1HVWfHYCfDwo5tMnredqx9D9LTEEDCjn8Mg9
GI9QL0ueYgbMBUyfWm6jgAG5MKg7a6t8+SRC3en3VdURrsER3ve8oGzIUOEz9RWW/emfSrpA6URR
lc7HyZnVAgYEE8+8KvEA3EYp6P46sj+bjOEg0pFDNZN7F46XH1FOFMgpmPX2X5zmpHvYT/zb793r
IcRBaTiGH5/I2nvxmysLHIUWKFKgUSncwYFEjc2Un6vn9wJBMSZZzHWyUzNdb+Y22hwNliCTFYCi
3hkVxxl+3Oml3vK1UB+TAMzX0KBIlAz29bJ36wdoss5XJQcHsnQC8kdRqunuLyle9yx8yLEr8Oth
AHBWybHRgkV9ibmiYk5oxXgaqHyaB/86+jqrrZS0wptY3GkZ6pKsoxb0sIoOf3+L0H5bACkfdQwF
MmAPPuFTpD2OLAtH5ah1XGtD0PetQb4lMBNFQfvbd65xJTFV0sO+SFFc/kzfJs/r4MfC2I7IjTsB
Y5jJEhqwjaKAqa/emYud9ovjIoYJrWnjfZU/2Gnx4tJ3HwjwPzqGFiH+zJsAvS6bd4zWTsBcrWEt
qZM1uWZceGoFNbIj9ELNc3Z7Lz7+42g50nw/hHOFDxQe8iTJVBp57DT8Pjn+ZadgVEaEKhICG+VZ
nNMm09LOSvKn65VCJ5Ug1LYNevl2iGzypk80Ec3bhQdEzAhtlRSfJqIv1skxvVf+3rrcCbRfAYK+
0vNqOZoJh18phsRYULZR03OB/gGVwb+xPEl83QFQJS/wfQuRX7bI6SC0oXNN9WwP3WNugzBgR4Hg
bC9wBbqR8ejVkTzvc43EExwqH0UMylZeThfJd+GU19sstSzttoz5CbNAezYbhwtbBEFhRcCfzZxP
yeazFxM9NUcy8WCH70NjVpTLrEAHtoSgBefKkIZiwH08FZmgvkDLL9ToM9gzEbPe/DEIvGfCPln7
u/7zb8/TYSWpVp+9qE+dtFbSWeipir9NlPD5JXWRyMxzJUYmbVxeI9c3SE2WtlCOGtotZXYjiO6I
mcCDWeTqyZVXoUpzKnDdLVocP64gGPqKUOddLgvacKh/Iy/bK/CNQyoKxEmP1MiFVlePe5Ts4kFQ
6Km/6AVAJDpp3XJwtLVMTp6a5ACtx0Ek57PLlPM0I7+zrzRo7/J7gNt7i21FPQzVBkuK8nlmg9Fv
85K0yl8ntfhSW3ChTkr+JXvZkELoHYkq4lISZfoE/ihUWqkeLMUskpyorAjWlTricJtrGc0GMfWw
8tSfbOXOoraLcG1u5IjocZC3FCz17gRtpEz2FbtAoAa+/SwZBR50iZs589+HaiVIM9jvdlGZl8Jj
WdyCU9wWb2dn+Jm4PekQ+AGXFN3wC7w6aHFTNhaE4hPRUCEW9nJnRnuwB2BOzjBeoWm4Gm9SpP5+
jYmvyfaU4AiHWt65zOHNB1WRF4lDyUjYlYRtVt8fklGqE+woab6bKoh8cFQnMdYzSMBjs5YzvobD
39stTG6gEllE1ykRZHEZnO5V0n4E7h4lLwp7IHujT1noEy+6iTsUazvZHRyRzrmGFI3Gm6XobyRm
cvqDyJNwVzOzqJek5nz77RVUNkKgoP8KhqCGCJtns1/5cqhOlgxYi6r4eSV5nw2PL2/xBjDOAVLx
UNFT8JmDR2kPeBtizrSHZCy71GGNK5Am95Qnl69B6he105hbGtt1GD1gxIpbUHccdZh0wc/Z5mYl
skQlN2jNlkWwL7Qh+Sv4ZIEAmhh4MdMaukJpiu5Fyyw0+MYq6FFvBFd0f3erffLQ8oNc8lfAxdKs
s/zv1jVtNSMPaYG733tKZJMAB28lZRlJAo9e+jfEDoR3D/MP9ha24KxfYTQxYKVEt8iLwpe3jkcF
n+QI5I+aW2xX/3ZO5eXPu+lUvojbv7gM0PfnIn2MtkZIc2fFA7rLPYnKaQUcoB79n1PRBzaMI+Sc
kHq9rTaxdvhIA/BeXzk+FxeZ7jJg1NKzmjGwFzDqq2WHBBT2MNe8PQWbXwrvTNznGwESoTSSAKp/
8EDKlUT083tMz2qar1qMU5DL8UeGVG/ga5mmQbU4u2mMZaZAszy0gRGrXIHnlJ8mpLY4meW7cg1n
OvnyIIQJpFwfDGfO/g7Sh43vRkV3LrM5fhhxaLq6HIto1sbqFsKppeVuFmFwzv/7LaV7qwV03XNj
pUQsvaNZKK/0joz8/aue+zIQXmshTIiB5bjZMVQd56dODNMd1XJlfoef0XfSRxGSyMp0EzViLfhE
13zEo1h+lGn2Uau2ELQSvtsEyX05K6NUoLAr1YcccPQbKsC84hckN9MySUPCyahd3stWa7T6Wrar
XKciGe2thK++ZwhEypw/0YjJcdufjePWt2UT7BHw4DPqYseUAM4vhPSXtTUMwAX/ru8H+WjEWQIj
1AZE95BD/vF2LXKTyiBLUIIhgb63600pRNigrIdjSmGCHnl5TEMgy2wE38hQB8gxQ/1BoDRjYURA
jIL7bMVu5mk+4oWWYnHYsFOQITRFz/bpZ5ZVNHTglmRBegBQ0dHRbYvrIUm4+zf73P9XP7DV6B9p
5sBZc03Icp+EVhjFP7TgWmuOsP3e8mDx+kvzSybQgztrUe5pNxEkczblmT8c+f8s5hwf30kOJ53M
Umjiw6U42kugi/ooWy1/tmOWVkFtGSFrClTMnuqznPLl5rNRSW+ITb4QboCz8oXacahyt2/wdQto
76blTbTwRzbAzA/T9+rYTGE5s67xqy8g5L5nrVPcuIVVKjvLvNzVk9cyvuid/cniQRA+6sqyJfQ7
P01wtBZA+M98rCHtG3PWg6SjIqDF5AAHOEFchVvj2xISGoTuAxmGc0HfP01yNRfSUfyK4JKis1mj
T2BsccjAPO5w1haiPdCbGyTn2tnpVJo/F5mSDpNqIXuK3YRAIJG2J0o+IOqmYqXjvUV6Ib3Dgy6l
sJxRMtNj+5Qwi4Yrn4X0p1V5JoV13dKSHEV3rrnMHilDaPGm1dNkqbAc7aDgDF8eynaHKHA/zh24
vzlfe+kbXd28OS7CKjrr0Ux1bKJHZ01KLhc9P5HgoFyrK4SGPyIgv5WqzVlA0bj1JxZfGEErt6Hh
p8n3OQfmdQj3V8f9G9CbDQk3QcHr8GVn88SWlH1R64eqACLZVWMaRFEj1t2saeurS4H+1lJcyWWX
YxCmJysveewAPCgk88WjlF3rpN0RwWB4PU7FXnx4saCXEMiQIQcrowIkn7B2MMc2ozkiI/v4wYe2
aquaKQ9F/EaL9P2zg8szRVx5p04//HPzStCXBcAtjSYAZ6o8qYkscuqGHohpjoOBBBUVbs4n0lTp
ImzdvXfEdBBEW2UV+gNJDFsy80YC1kG1uRFv9AJuTHeTDB151ZuKnw7FQX9aVeGwQlMLnhxjF15j
j1AVl0cqM0+xZqi3Tdpo/0gbmC4+HIh/EfrYEUs7NsSa2mI4tDtEk+vqbTeh556Gw0i8PxOykk+Z
2sdMmCen5Y4txGRU76MrEC39V7TNFYhazlY6uSBw3ehfnQCVwymd6avzLo1ip0rzHhDrhBf0a0R4
uhxAn4BtSKGW0szI7ySGu9kvfDsjBqEK1+sp6V+rJ5snRqNmOTSwhWzKhgTrakBr0ulC8zgMnpMG
TrKReiKweFDZVNteP/ThE90Q4eEfmKfQYq3Fn3+I98NwJtnbugtC1yywKUi/ymVt1MOJt4wQkvSL
dq2Tv99nJIwruwoZFeSTH6FxAKh7D2CrgsHXLpsaqRFKzASmNrkzw4HgtzxDInulMgPUZ1fCk6yY
PJfAbwNfy2qDA2Tp7wQ0TvmAOVGOcAUNZe3DP7d3Tev41w0Yq24VOh6IgcwW3U5Cslo3fsMrdUKf
ICGmotDecoZ1iTk+KtKlGJ/d1h4YPhDiMTijnlsm2W6gWYLZt7XO3clQiiHt4YF7MVpdl9XiaItC
vc5knvYNgvRSc8SKuECblc0WB8JA527Ep3Lphg9/Do8j0WVo02m/Xg7Zem1qUqbWOrP7E0EO+jmb
tPZANu5wjJ5CPBsJ4qA4RvCm/OtYnPUyCVJvtsIdYXisukXMX+qfiS/NokNsIJqSzcq9hg2r5gFf
G6xusHkDHH00tDaHNEl29p0S72cjHa2XxUmuTetIfF4GZScPOvoNtZcjz85hTYN2I3/R+AbtqZco
PLfQgESvk+ExcJpFJgWJMJpKLrsH5lo4j5b2OAGrxVG1XtVpsBodwMAahUvgO+2NhTSNgORtS/9K
n4s5/ZDHLqpVAAe7Fok3Za1sIQZT597xiU3I/cjx5+6QoNYrmTsdYQzWKOOOwqgXhC6uwocb50UF
nLSw84XYyvCxUm+va/x14LnAf+awXBFiU1uvolFwbYw1P/nQNrZ8rY/WZdJGyNxysh4ohqpYL8v+
sMMi28Pxdl2btzVyPxguKHuHbDpDd0zXcWCIjTz9LJp0O2IT89FtyUN21XYPSxmqq9q9HKOAEXAH
SPWbDr0+o1uJut+x7HmWJAwFAciqur/ikISxjYg3dbXLUd3nxPySlS/6PGjilprMNqbt6fk9FZ5t
gtUqq57EoFkGKcEax+b672AE6R4f76GFELyIzw/P/njob2xlyUhDDtcGb9i+/mZpR2+89SoCi5FF
zVUBTdraB0PYeGr1sYpGDg96Ortu9/Wx+lErjx6vkw0vRGi6zqgToFZVETVyCgYuFL7KskPDt1NY
SXzcOClAxX9nxhCxm1CY/gVvyUuITTFiiL0jD0F8hV8DdgfcedXVuEOxH2VxU6Rcav75Xf2pXPk8
sqJeklgQ/PWcBnyUnDIisINTGJq5KMUrJrOUphkot4+bMqIEaAOddnx0MwgKNprZ2Q0UA+P9daI8
84n0xygdUKZqpJ+9AefgTpOP3gJYV8bMwKycjSk2F4sLyWXFS0db03xskeZZEc5wVpBHCAZ4BjhX
C+xWiucyWddegrHWmMYfFQvr0RPUiVmD+T2krbf42JDOrJkRc36URXsTh309y1S7GlqypH+z5kA8
8GDw6HqxSBwoA6dzxzFOLXvzJJp3BR0uYYES+eL/tFahFHTkYt4RgxB1sJiXlh7zl1mVSuVq8dsA
ra0SMaRzGyTn0Q0ZgPs1PWR4mEhvxeQYQMFsyrEHVOOJ1qCM7oFJS4wE3FJ840mGKdKAo7pcYjwb
UIJPlWktJ9yOiF3LcKOhd2Rcv4g5xoUmLJ36G1R8bZETQfSX761sMesPLWJhI651V2kg0JKWbYEp
VkFfwMIakTbZn9Z9o3N//iM0UJUi4K6QmBVPQDxZ0PlGvyy6lIohvLKMsNlLwAwTFNVaddLcXDmM
97Ozw5/AEVV4pVMGNAtdoOiKQJ8imk8Vl+hG2ip2eJDuJh0duXdf3Fxdmd11uBpw/Qo8UuPxdW6M
OCfGK7fVd8QjeHcbg8rM5K70sfKNhmOBMH5V85Pj7Q4NH5J5B4wUSzJD5K5p5YX72rM9ouvAmCG/
UiDrJcgfkw1QpUqquAQIfE6/89XR8dlTSgfc53mGQ5xrEn/D6d1ODEImMS5IlNahg1dCQ5qPtmwN
qCNipJGavPr3FQMK31RVyOZDnVsdo7DQDOg4Pv6qyJ+P7LiU+dGCgCiThNr0tDr7nG4iNgO0DxgD
QArJxHS/fqHOVnW/osJetdxWPh3nb1kqgHJFwd5GOzPjfTnZ3sY5nwyrL2NfQWCSlf2M5zfoJGmh
qFyoDFwLoJGHwogY8tg/5otaQNXli2cKDxDPk/6hKhYhDSO6mKWCG/W8yCxtVOJ8+7JYtd3rqyFM
IS6ZADYNag6sJ69DrQneQiF7+QQIcrQf/Af0ORu8ZNBFNu5hReUhAbbueHLMOuI4+6AwmXVSGF+B
QEK6PnX3SGH1XAnVb/0wq3pAr33EEsu1b/jhONbIENlGppagUKCI55r4h5haieL7RsgNQLC08P0j
6Tqyh4tIeTeDKAiNb0y/4Rrw35wI7xC8bkkwPKpz8ao/leUqG3ZtZ4cQTZLrvRjCw9Vj/hNyBOqP
KMAea94sQL0XtIE3EioX1/L3d6lEucwFGQ/TDQ4ocZr0vUMBMSqQ/MdxTFUor7Xy+OC0xJA/V5hw
Hje7H3uOOw+4RaCPgP/j4MjRJ8OYydDZBKEzbfY9RdOQsYmjpsvRedyAXL+A5IxkhPXKo10TC3gV
g1xRmqaHxGFU/Ck0a22TzheO4gLEYxg23G18E0vP+4tJLYm41l7NEuLpCOuBZ3d4spwa2vr3+RzK
zeDs/PTUgFR+9flKM0btvmSL9bCDLlpDH5J91Fg6KY6qYCri1pa3wZPgiyksrHhXgC0qUWrc+AjY
YcCiuZ8NRTrEC/V2l8zB7m1PbI5UEuRBaFa8w22bxIOFe3aH7QGKNAauzDq4BzxHxSI1py65eD5A
K/RESD0c+Juwan5ht2FUujzifhzDctAP60BFC8KwFjR3C8TWOS5RHDjCYU1/x81M4Xqinr0U+aZx
TPnmkzOI3rLgHzTcgQj5VIs3wjuktBoyNg64dPNUC3i1e6WKLsNT7vCUdWtJZ6FitH+Lz4zLaoep
vyt3kM5z8T6IXaN4HPDRbO7rtEPFDKl35guzl71BA0fD+GzgQcQ5KFicYzUQzUTz6PLgkfsFXCcd
AZPe7eKVGeiD5zD4Kn0L3jtMACOfieCPBZQVukiXmFBLVPRDckt03feNM3d7KfQWQ3wkhmopwPVF
PvCu8LHXKDXlBJQr3UrxQsIHbxKVnu4RlLOpSFM/g/9O1WOYmPoHIR2meT2ywronR7wUAQF1ERyf
mgCBkf0FWx1y91viOvokEHfLfQKR7AHsBv27cJw5koqnjEAHzIJRwCdGxbp2xEvU3eOJrhcb6np/
Hdyj1V5cSWzEfp8fidk0O5M26dZ3pBkT+gKocqbf8MhG4nuFZqu9lzCPg1+k8qG2ZtTbq1Y/jj50
pY1vk/An+u3B9UHcgC9vJcvre8rpnHEPj4ul0IU6cNOYbVsbqCRRMGUjkzvEJXnlYN71IRJHHhOI
wezV5Vj46s1/oXc86uN3Hi4r+ozmBAeIoTxrDPy5Ouh1QWSsolLMIDWxGbgr3EDBQX8RrZSCPyKb
zcHWMpp+iv/fxhXkoalfwSpLQcHZZE91cgn3+XQMp6CJkpo8X0pUfd1tTagNaZKNB+z5gZjq+iwi
QcWU4xbC+8KWr3g/tvOrkVFnwmhV/VS9lUOGyVUFB8jYCdgn5zR4RenyoFK2cOFzxYOVvA15RLAd
UkJjjAdUIfo9Or/111LAZE70RSsWE5uUqLb3guICKtIFvyIIiehi4QlWT7rBAMeqOQy9LNmZqlaD
kBT3wOI9UqbcGN05EuwvJXjefMEjFKrjuuZIxAGiqljh7BHvLS4r4okYFVcDWHjfOIcrDeXXtUfi
9E/lmjIZEZFQ8uclxhxVngThpQRKjhC3oAWcr/L5MXtNCT6Ql3CAjVCLIFXK/mohwy91jMAWqDBA
uY/CIeRfWqK9pMr20oq2zsnypvTtkt8sOb7bsoy0Ggq9I5t67kq+s6GkB+IlEEhw5A3QGD7QwhGQ
PcR9QiGwwqNhWiloCYNM9Tr3pccXcAsaw2o8nXQtBu0jws1ArIEvoCcv2j+JeIDNX5WVgZzzliHk
pcMLzDoJAhmhb/1cA9Ub2C1QaywV1h0C1DYKYETpC9WAwJMqh5Egdu70bi1GNJU/5AwQtNi368KW
u+j5mR8R00Ca0BtrvRx0btVb9rgclOc7d293VwcEMESs+Mwm8i4XfMgI2mNCHua5YkxtRAT1cpBz
SxoLqqBmbbzw2JxbT4jUTDVudpE8zVxDXjJN9iY42wr9dPsAxHwEwoURK+wyE9rzEiFFpLIovFKO
9kcaBNQC5F4bUpE4L1ySVpqTqAROenyt8rAejfVc/2Lc0jD5c2QFEPkAdfcWPPmj5pxtidcAE0j6
j/vitZaOFcYo69WpuNCPCwD++EhH/hJZeZhcVyOryxX6BerhJrpHuma5nxDvGsBxQf+WdW5nPndQ
XoHLgj/HUzFEgNDprdDHk8A3Xzmxiug5ZJzZg5SStSTsOAZ/8Nq6Ne8MIZeobAfQqbxcB0PD9ANc
Bm6GrAk8I4ywCLzJdYNOlzxaEslASuhGzo9mmaDVJe/faZbthasbO8madbfG1VKWhCMpmT3fB6no
mg8uGw94H/Id3jxa6SJXOEzB/9b1NLnYYdYHuwB4rTYmG5CccAs66CmczvLYlyMbrWDgW/o55LYa
/JfPaOjQmccldGs3a9zybn9ryvUbLTGqb29sHawA+HfHQwAn887U/becWzHjHPMdp64DgjqgrciP
K4dbEGgCShQl6PxocHjak26QnZ0yyOVmnl3xmxSIBKGyf94BBuJ1VoxZmkKiux+C4gdfPOcTvYMH
fFc74526+A0J/bxod9ZH71JFeXc/Xr5An4WFJdKTxu3NAG8DAWImHNyKWQdIOq43363rUA09sXqa
8ZESJhNeujen3SVfCIXW0OXlXbbngVSxJ6/Npx0h34ezElXaMUFogrOYpDCW97SUdVCk4Dr2nRXt
CBdx3QAwF4Q+xENGTY1OFxs6X6DkYA+SS75SIdEL4TvsJxiX4qndThsgSrzCZ5Dhxp8nZXq7HcMM
GK6nRetTS+NF7udRo+/MtUB7Nq6nzOWLb4+YlYw/RuZiW7osHU5GVrRiVEkUuV2xGpTmJgsdd+U4
fwtfMlob98tJfd18Fo7qgN3TPWeZolpb9JsIROdFTduTffKCGGfU5qgcB8foGG/Q63m5ylkdJ0ZK
HGKUBX0Dz1Ib0Mp884lXEXp2uHrlFkiOvaR3RrKNbFSa+WU3eI0F+IYguewhebn3b4E+HBzAzKLv
5dkj11KuYDOoDc5Kz7RAxG6m9gGyfyh6n8YseDu21XAx/wHQP19ixx2rgjUZ33eyRnZqNFA+SubZ
Y1NO/ouRVc8dLgbAnZSUgoY5j/u2KJKyV/MU3A1cmEjAeikICqpVDJ1dPqsJufOvNAGQtCkNEjga
NiJOLZzQs984t3RoqyMcJQ624qq2fAS308wP+SQadG946RnIfPrNE7AQMsO+ghZZnICHy4MJOYlH
EsUhjamCziuS8XKF6eMeKHaD6mniD/FPK2ekVn1ncB3BxB6VtfEEGWMT/MDvEnGwgDdgLqmFQf2u
i6zmFgmPral9zMxcqr813nCwmL7F2cC6lIP3+HzhbyVQvVv07QUm1apQS60Mlf0FEgTT+2uXUttK
c36XxjhE8GnTnT7mAURfBipcGXn60i2Di02whdyyPhjAEAQ5+ktswSMalNZg/BtnV0PNLXnSu6sk
fTZZfIVI+lTQZ7Si9bG/ika24VqQgiG2ptUqU5ccZu9vf/6tj7OGWd7MNF39cQ1zY5tU9VVzzYnA
77/qKjYRucrpHEGHUmHb/Z/7NMS8vbhr2hIDDxEiCLY/3yhmBgMz5L1MlN/VkpXhkjYrW3lVGPax
YOEpt0v1xj1K0eNcxwN/kkqJ33brnVp86G6TGctanNNCGaU7V5zprHxkB/COCoSu5XdF9Ebbt4Pm
JtF+tY2dl8Qiv9HJqazUMz/jeII1fVD8awasTXEExeKR2oC4Bdqj0ohsdBou44e7CeRBG6Vn/iai
WG33xWQ4E/sHoqjPL4w7EVqNuh5YNGffbxektqKxogfATK26lfrfZ174S05B3PbQ9XXZ+em3Ad4M
0vkRQaDk0yIvpvFKYKt4BQpBekd3ouWc8aQEgjfOc3Uh344isfPnpguHJ0syJAybayICXE2Vwwh/
ZgKqY6NHSqws0HhRJIJjtT1pxZZvU3Tvzqq7QC9Qeyc1hp3shmOMOvx14DIBe8X/UCnSn6bePaci
0/dQgV3chDEOjxmyHTA/GxK7M/5MLmgL2d6a9bOwJDIrnBG4aHIbDQuOl4uwJmAP5fxR7xEtUj8j
gqiUvGo4Oelw3l6bRh7pVRHOq9WJAVSEZpqO8k4zAnlECKcfqvmkYQwpa3q/52pRBuS8PAUU/39T
OGce7RVxPPYLrBHQeFZ/sFK0WqEetf4dU09OD+oGOYu7bccDoo1InDFF3l575KlfTlIp2EEMZqq/
lnLnqJdxZQl4sve744HTpHfT7KSDxz9+q/yIzs1tKWs6GJClymqZAPBRY7C3J3YZoRS+ri5+/0I3
RIG5GHS5/dwqINyjvXXUl2Z+yK3uErsv4IfB901ozS9jCIRSFgCtY+/9vVd/DEdete0PIujNM1Xm
SUwmbO/a82wyfN64/4uMd2D1CaKBsF9m3MXOH8S6Ji6YhlFb2c8V1FmY2pSbQYb/sQ82ygw1ciM3
cyD9ErjgiPmGfBf/7p1KAUHb4GQzmaLjfVOeiiu68akKst1GgR+TPpZOyZFFx0wASg7tKBFoW2gX
z0Cp8sQW1Yj6ueEPEku7g7eU7VI0/HzEOpGWbg9wEkSO1bGd9lljzFBjnAXMn4M5USPk1z7i7qJ1
jeSPvgioGfD2ZgzTFUVkVG8wpWFg3m1cQe5UiULedxkVMbwXWfZnTVXbIiLnY3PS8gADKq3LKbyZ
ZT5700ZcMexUXwi9ILPMSTiyI9XsXB3t1Fh9jEuTYwHunvGfqW1h9B9fxDutLx+msl5Q4NgzgAre
48tYMvsFwr7HGRIjUpQ0ZvQuu83zX3gh0xzsM2X9y+ks8GnXNgWQ94Lxwze4KK7t6zt0tyGQPU13
DOIZMmMRBQJKf9/MiWJ/jxF1027D6vT4TjU/N7wZJbhDSGrUReUGPVkKLor10L9l6uNJBhI/NYsB
lUDrGUL4SckWEeqkPo4AFLyMc1wuZj1Vu7GCfOow2OweUrZ01U/oM6CS1MRac4b88MyePnKFOBgX
AbPdA4Lt2IU66wV5dlbcvvzR/g4ewNWp3PKeJIz68ElxgLjRvlJoK+ULuK5WqlDK9OU5qEx3igYt
vK9g2W8zu3Hd5KfTuclmHeeCCaRFSKLi/EC/Ps0cE2PBQyB95Qvvo6C2jQuZQikrobthKiy1rDI1
VwyVRd8qbloTws3mVfXjHLtR+EfnDQP89UWgb15zUnEnrVItlvffkA5UQWprFglkddry1t4Kmo7r
wCx1sCZw7pSfIWl3Tpqyx2SwFte9UtXqDp5Y8N0RrrHq/hAeE0ZEyqMW04hgv8UsGOPUcb51wx+e
zdXAP3rag0QOJ772yWTNoUmhBPny1jbp+eG1DWFmGICxAbgYpYSFoMpILKnLYoUVBAdjxRBJWy/E
zXy/fc5J3eOBvV5LC4K7bpwB7WR0Tb6W2297q1xQfhBifUyp45H5THVvnfP4SRJKsfQj5QaoXwiu
P3H9GQMMX/n0RrAPkgqtX1o5wU4m7blC349VpC/odXRFwYMpZgk0DJDnozBaOYhi45eNJRmAOOjw
CQUgkwK+HSkj2ZCLPZBdkaDvGCYiKZDVqZM0g7H31Vnu2yd0IjTYGUu5GNtJD+16lkalfge1Yf7I
syJ02eoYtU+/M/2ZPSeE4JBhwjBAMQBhHaj6PxWDluDu30f1A/3wYcAq39NioffcvOvyoqzddOvw
/+snbVCiQBdR+ZedKVAZnVXZryZyfCxE+6+KxcZNx+apxzpbQIKY8vQLojlR+uM4wPEHqcpOA/ni
of9drZNESOYuHqfmozL54rjQy0DckRe6+Hcv29lzNqe5KugxFHhm49k50VCbZntT7S2OWoX4vfGg
jtfGSslj6lrChzhSbp0hDOWW+af4+UfPsP5FBgtgLZV8tgfQEYxJe+gXMtjc16cHmKsTYsI03Cd6
U+Ms24Au6FQPevNAiszl8gApl5Y5hiiEruhpZRnfYzSrE18rS2Fc0KIp3HbHgZFtTe+D8ruLid6o
879kku9FmNnEG+PSq6sCMktVXoyZJgwheIpfKqoZiJgE9r1fGbdwkD9YgvVtVZdlkm/ocjtad5cC
chMuVEs/Gi1BUCYcQ7k+JtKykzT+/f4CunI0Z0KSfb68pbPkQlaszg956qfDLF+UX4MJ3S6yRgAK
ih0Tk35j7r1yF8WVWnPMmzaxH8nKgQg+BhSsRYjPohDjdCtmBuiNhAKXmRn3TeFXsbEjM+z/9/zs
udV0YbaZxovtQUgmXnTzVh5VTcSj5n6wzANAuRHs9snO2tSFKrKdUuxOD042TeaT67zsEstkna2J
GNO5AEJd5hjPhFczeHK6BEtLFpTYU1+77sbPAtp0JRu9XvMM05WobXS6X/ax5BG9BDANg769Ny9q
bUkskw1E2tzKNJC1pLEPWWaG01tlES3h2P39LoPTBDbJaDwmPjMDDqQt7gxt7Z8CxYiovOC7TClu
+WubsMi9o9Va5NPcVDM3QzDL0ybBSXB5dEZo88i8Bg1WrYdJ+PIzgFmobbmtsFiop6KYkJBPrFeP
9DJmxoVsfykzuf310Nz0OHqTlouMGkRY6Cr7NSi9d9qRo4ons2Cwj23A3JBifEyThqCuhUG9yLug
t2exg4BznMZ0n7RVgQSIBGaY6xiiinOSOOTw+Tv0DK1pOGOwKhcOm7QpvYIAyGE6GHHlNeyKZMYM
jZ2EWJMLVqNXyh++uWMlV83iBIp8PQoMxxj9ySst5AgRyUcioY7AbNmyORqd6L5e5LYodz83YfFI
Erv9dO22V89eBrg4tVY6BzdB85dE/IChLdAkrUAZ8E5pKg0ZNPFAY+o4HVGTD5JUT4cfsOdmlrxF
qz9VtiBdDTmIebbHqxxLWHdphEXsHu6CnVKp0+HHrEa0FJoc6MyB8yKo6Txy2pbCEEVgudPePZyL
bT4bVaE0nkcHyAOkCVDE3PvmeB8rYg6EULLU5Z0+Vt/2szwIzwOXlV2zzfxgMewjqXEKvitbBJ8c
181MwXvpVVEwDF0u10Pd6c9bkSX0dbBqywVRu7Kg0PD/QizJGjExxF/bfgvzxoEktY4pRQJDbyDf
TGX1S76M61/Hwi+YD1cv2zvcv6d4BXfUfi7F9iw48dVWw/y2TxFSJWmWyu/twmo8Kifrwwql32G4
BssvQ12+RynnIRHD5kzZ5BMmanbujw//iAVe+HiqA87fVschqPGCR+DEX5RSaivIOhJBvwQ6UpoI
t5Tddr0ep3RZaFBOTAhphPfIJNQUGGU2PAv2ZrPPQ5kTRymcfV1zQIEl1ZxCyy8uN7ntSwKOZR+a
s8XNlq3uL++E/LVOtSfJrN16ZZKOsgSyBOZkOwgk7Ga/evKwmbAVF3DxoRSubJ3Bxh0ja2SyfCU8
ln8y+Mm6mlXMkXC6icljznJyUCWSrRb8aoJX89iB+wbj1clYVpWT039tajNmqRolBAx/9UiQwlKY
v8fhzgMuADW6o1/HiMJ+dqLC37HgrbjVugMFEHqJAzBMzeKAKtMfVZd7Nq33noroTxFjoYO1P1v+
TpZRVbqLDaWsIsggiqj/6LQEEL7b+bsG0d9UhZW2B2wPd4HMe4k3a0F1N0D+qWcWgfg1+RfqW8yT
NnZu6yFVg5om0hP5NHqtC1EGNOIW3+C6glzDoD8M2D9JMqCVOkHqIACupHU8wVyvRb/YCtLVuhUC
BsRvYIf9ZG1jjGtbwkHCzkdb8cM+JpAtX1q4kHo9jvA5PppOP9uEUQkaLm6iC5nY86KG2bKbK30e
DUB6R65B7SBX5mb3Fl0TBGBEb2RJiLRbf1iVyA5LWrnLL3Vgk8OvZcx5EEvYUYfvwp8G4aYbfaCf
gijDLef/UMYNDGSMRl+BxH2/O2D733NM231vZoa6XaWvB5ukUuMDuh/7mCxsbNZs8s/CQbiiG/tr
bw7YP7IUtun39ZWeeHLACgm5/j23WU5FkCSa1BNqp16esxBsZaqhUm4+LJeQNOTlOLS65DOLaJTq
kQEqbpHabZabrHraL0taeLaVLs7tFE3qh52udST49o52vINrO6G7OsbdSHnHfQkkl/sL/NgjLroi
kt0lSNRcdLX8jar1vZkw9blBZ8a2den7MxbDyEJNkLHws0Q1F/OQJJpSa9nYIX9XiOXdrbHPOfSs
mlnXt8+H4FCkiG5Ubd/91Gzfqq8ClFW4Qe0R6W5rN/b1tIbJHtwTdG3WtIlrzkJXEMl2DqAlDgms
Zddq1tcvrv5zWzYKXRssmrlIR/0zGSybDWl3jSmoPURbrAJ7xFemo6MOdtYulvexqS3ScTr55uhb
VCLWSGJ54fQUz931XvljOebAGNxFNESS3U5IMCP1RtWgyAzkNAGcTk3xZ7XGc/I1iyIbktw9mo58
A3JPiPh/UGVK2h4HpHpOy0zHXIJrPEJ9et0moImDFc0ngCGNvGz1oFGzWFpuIfZXEXjodA2OrwhD
3gGoNfB5LhAL6rExo5Bk+Cp0BfUnGyftOrK2CN8pZZjshsb5LCxR+J4vIzFmIUIVb86TS0Y7fR/o
Zygv0/8HXwhtf8QQTAyRbVY0wU8b3u2mBHG1cIbg/usGuzuyBxjR50H/2m1BAIiHP5Glqg/RCBgy
zithIanDNT26crIxIWcAn1wz2Hx3g8L94r6cZsSJi/OnG+XGt9A8Iq+zXC52m4QAWX4Cc4NYWQar
Dh3ttaVWvqah/EqE6pW7mpUb6aPBEQ9Mu2x1H0Ci++KMtAEOuegKtE5m1wR8KrsgsDru9WrMgl5W
RNT3UxS4Fksn6AD7E29oLX9xw6C/KE6bQlmT1ZxaTKGJkrARr7SejrpxtvBDIoZg545KLsWm5IQv
fu7RR+ozZMKPfwsAN3i5PsKwfvwqFSszUJ5by3LYRu7oowmatxyf0+JomsGguAl69PfCFOWEAMuP
U2ie/LLg6oQXA4zc1jWxONoPfIg7/8ZlHgeZ5S+8tF3+ci8uGE5LidhJTnJ7B/CijKF3D5e95TM9
MpKU8lux/PUnidi4mnY5xFr+pjfKs8FyMTGmh74DmZFytbjkCejjZditT+5Rl6QK+L+/JcwfZBzs
OQDHL/BWhJSqgISwGU6Sb6V6jvBXxCk0Ji15fzVd3e8bSrbBHRI4PMYsaunYpQOmnnaOFNt4ErjI
cRMFynbBJlBNqwiyPM1I19PWydhQ+nLmVo+RjJQSeejDIaM2o3d0oX19a/Iro2600St8TzdAxFHd
qGwK8A/UT3oN6WIxyAlL0cmg7lVSKzxV4PM9t3r1B7+aiOUPFWFSw2bMLC9Q57C/fhi9Vv6+c3qG
cEBFYYztoLjDYGyU0pO72ZqSH59qSgUNmjNtGHVDA2GgRux6xVcp3p7kDtq1WVRgXdPGeKIrrJHm
Q2IXYpKxxs6H47ibIFnZfEz0GE8+vdmWpK7U5dmnsmq34I/b+is6iq8dULFlOslnlEh4hSNPuGOf
aFGaVYhnGITuP+BaOU2YnvHXE3SKIDFS2IXuGd5iXxCqMN6MS0aeEb+KMzJrkwOsEXw0uXCAPbWp
7dh/YdLKoKuc9IaG9IGdcQOQsS/XdYg4QBXuoFUK8wYt5LwisRU/j7yDqtCJCOiVAdRrddfvsH6r
rM9qX7ZXhXLb/65K+4H8fMEoO1cVnq2BxsUiviKH4p0a+XOPdqsr5rTemm+1LurMBl0qc5DOABi1
vxeozQisj7BaogGncIV0pJReWqwJuX0OxwGxYW74g4Zoqj2p7bv8aDOc0OmgrFWrCaudq1Xp6C/F
fwqACTmXjsfvkx7ew90TRoIVOrRdiVUR+LUWnZXzbOvfvQU1x+RG8MZpsClyJss5JiJsmaosfo1w
JTa+eXI/2q/4yzgA9t+A3aegjEfCCGTs19frc7A1YfDlugktWmAukvHQFyFZ4xf0ZjIkFbx1qkmf
gj1wWFyc1rZlAp41b0G+Fu0/NnVv2TSBtHgqQJao5X4qaNKvcl/czA23/LlsWKKPwJLeqjI3cD3G
QX44z8qrOMy6cvSsoqxgWW+id/zAb3gy+nUQj/zKiliX8BVtN6Ua7un2PedDwf1IhnKZaPvYsDxY
ekOm7Ivd/5A6FMYcUdYCEmuYrzy9/8agoQzdqZUyB2T9v3BPGeFFedFTBRcddJ7GyaRT+uLScRoN
KCEPSL9hcCkg/25RxZWJFjbhww75AyoQmS44K8N0q8e71+g/Aq+rksSN/Ml2dajXFPuubNEfu56K
D93H+MnmRLoi/Rh/AqE50ub/EEZz4ZHX9JvY1ZC9WuBGZPU7dCHdVQ3Tf0Bx7INPJRI3Mbj7Ttej
hoSu308tt3esaMJJe92fiYg1tJwmUDjuhoO3j2VuS3kZXBO/SGmIe6I4EG0q8yPOQ+3ezdtOAd8A
Y1g1OFX95GIv1Kl+iHWqFTJNpP+igR88ny/CNedxO+0AubH/PgK0hM5Rizg02mat7EAorbSa1LhN
Z6Gyp8+7G/hlwYKWYCHflX3bgzlpf4aQ0/K+GVhwLmjnrpuNaJgQZs90ghPeMIQip+2RGqnzHLHW
NoYT0WamXyTrCXGn4aFEQlzCIlOvILaT3XnlJBHX4Wm+jfTsee0k/PNXZ/2ntog+kAcyCaJTizxQ
PLMA1IkKWLb7oKMCVpkOyU77fsw4s7jmReimTauuSNKXs4StPmRlsKVSI39IABE2TLTQ5RjY/VuA
PU025HCYqThM1pkWCpuP3ujwE0pn+DyJ5F6zGcmYM37DQygAup2bWZW0gCpO9XD4MmrZ73hSBsH8
gjA/FHwWpA5txYdQPEd6KlAB0/Nbzj/1yyEKbGpNSdQZzuRYV9V0f4xH1me7aHpLEGV1DFmlTDBc
d1k/bYgn8sQ3bTZ/Gngq1k7ILD2tC77aPP2zIOv1NNk4m6kV8NVSR1e6w7JY61UNVaY/b56QWOkG
r37XEP8vCpF5jH3na2vmyOh9NEI8FPrfXDeS/8eYP8LHc4pR7eTdehyuu/QHh0CVmmf/3fR6uZ+F
kni0JhcqA8aKEBTB6FqmHU9k0MKG7xMO3SOKix0BzmURi/CDyK7POO4rKEH//CpiDt3g4YolPdfX
38O9fj5+A/SciYVHAgZbu2FF2OLckuZ4o3Oo0CuliIaT+3h5Wi/zUt0SoFpZl7QgEp+lKM9bZ+G/
5hypW0faFc9W3JJNfHPjw2zuo+EhpRZjNvlji2Zvmat5jLzsbh4tyrxN0O8NaYSKzr4Fy944i0KD
kLQi5t61ZpcHOBgaTIKVc1i3Sz0/CvEyglpk2oguBB+OiGJ7F056B7S6fpi7lO+YskIHkVa4+U52
qHKvAYDidIDNEEgzN5P/m2cLz3Lu/ckGWczYFHjokNlmtRFF3rkW4nd8X0pLl1UTHm52sJlsunZD
RsohBFIYeELM8XQvS6R31b9lGlADZvcj+NmeA/YbsW3+hAkNpIWnYmFlHhjYHqmqZMHgSgOCx8p2
BORCBVf8oUMjpXd6TjmHnTnqFSDDVAvxCC/M80V+lQj6/vanzI84anP9YzCLm6a+OTObpQq3Y+Jt
9O0r9N/JjbVONhnIq7Lnx7eVpc4z2n0O17YT0X7mbwWc5LxYmh4v7k9s9Hq5iGHZlcGOWEhKZYoF
ftIh27xXSoYMTJ9gTSHC4sh9hwOnNr0VYf8gZwfXigmJ8husZ9qHmo5I8os98V3Bk5BPZEOPYYB4
SIrI7kEFoGx2svh4U39l953rVEhHpQa/ds0uaL8sTHlCJG4s//q842n66AOlri/U7lRz94UDsv8f
Knkj1sAbdw15nVM6ftUARywxRr5yp6s64F8CxbJrXIsSCiIDMCVN7RRRwH+rd4YfZroCD4lASPmI
jRbN8a4FzekYIiNngYMYzsKzjTyHn0gvB4iI2FXqYN4xdQ//PEKZOsGJ3Z85er5f8mLbAyJPQXyR
7I09YP/gUdrxEMEAu+me4SpQuJqkJ2qevCLx9x7ACIatxV8q3Eh7j8GieZWwXj3FR0ndfT2etGDc
/1+0EFWJj3jLPi2eJ9guE64+rodgeyzSmzQeC8YouJUlFl93KLBNe5CgKDKm6nJ45GQD+/DZRmKX
VB8NArRSaDvkzBrFnPubHHuoatjQPJi0CrGsuQA+rD+matCDZVAJWECnoj2QAX2rZ+sN9FSytFzn
QApu5CkXbTL1oA7wI1Yr8FtkhTLQ7GRVwSg7j7Yr0O9uYj1ekkF5NK9kPqhWRqKhHY4qb32/hSKx
uIfqAGuPq3hGVUg+CtoeunjPQdfbFn/cXdCUD/mNkPK5DVcitkUtvtmSB5Qf/xeFF4uiHwgk0LKR
oJEORme6Z4b5nfsRq3BT+KpAUmA6QdsZZhZYEwTCNNZy88EYJv1Z4XNE4nCYIZE53U0ZC/83fAXR
jskSo9n7huhWLwfqUJomFYahPXBgUMDicvoTBuRmBcbuiX5CW6EaNhvpAcsmJfxwJqobi3V31vNd
qdatFS8topHPGBS4DP0Ms7mBlnXONe3cd+GJxUdjT1dYXWrEDaYoZMfHPrvKbAM7hHEXNuDvdrXd
1IIhffu9ZhKBxWFTb7sSHmelt11OixUuR16c/cwzPBxauAvO06NDFq7EurfMK9JeJ6S7FRJ/VPzc
N0q2x8D9xhJ07IKM0f4k+qLzFGyjBe8/eBkDyVwWgUkaw8DZ44M6+IzeFhLAe1srptYRTcx/2Zf9
KEzJdOnPpEB+4eigk/ZVfOxIOgld8EE5CilUltsh1UqAXNToFma3RxdnP2gqh8BNgsw+JapQskVT
aJ+yvYd9eFSPSCeGDoF8+XGNl56vZ0MmGRZAo7wbFjkij93QCys9JkWOpDL9sMd014on4Y+tZPGW
xNh9JNtWJxxOFKGy9GqOnpDSvsjoAvteVaB4J3ZhqGsrxbUF3MKc5VNe8Ox1Mx6O7S3lfYkXFITJ
KPEVv7tQkf+JlYhJYmDGgm59OrbyH3xODkNcW2FbqLzfE9TElo/PDQznmP2ZMj+2IuqzR/KstZZs
GMwJO3NejkNENqlFQcdALorwadtmZcrErg85yS9axMkxRFriKh94SpMsz8pqZ68m+4LxCYd7bmyB
uRvTTDeB/XlvRt6IER9nVy8iRkYrJdV6q+GXeoxm5bPDfsY7Wg40cAvDcTYqfX1ex9ngGXeYWaCy
6azKTFGicggvVvxvFOSYwQ2+VXhlpmaDNxo605RUjgOJ9/2MVcSmvJqD8yuGUzJ5JHwwmol49Y1j
S/9AaY51cWajqlT/RbB7c0xEPxf06YuiVDQ+WcOMCLRC5S8Zbz1qc2sMGtWApmOyO3f+ulN2OSWL
eVu7cI1Oaim+b2fb4H8Cwa8ugEtAimVTCRPDzpjloXX/MehV0NNAT/SGA1VdpN36xvkw+y1fc/Zo
OoZbUDOxNd9ljcaeC9sUHy2XfFVkmC3+Fszu8PLU7a6UrgfENr5M4syqdIOYccYh+ONCcubFwwBM
E4F8kLcjAp4IGXhhCIdes1QjP6qM+Q/t9NsfHBelaMGm95+ul31EA3HE9ibyOvmg37+y6DgKLDU6
TEZyU8WhWFtvHnMyWsEGocIQbkFFlofXgVw20n5r4Re79Z2gYgnVJCapjWTp/Z1wIthtpshcK44M
ypx/FICvqIO9mvkD1u8ifXASReBeaLz91BV6JWgeSKdpmWaP1Rjquj1SFgLFEF4/2mgKB93obVH5
YD1NpcfgYyuDqhWt8pzbBbwi7fG/Pf470x7hMo5X6XomQmiMbT3KvtmZ94HPDUNemZjP3cYajXXS
uHVZ2X0dK9JlxIU2Ee3LH0eqKb+QS+aOSTIYSuUm3g7VZ06x2UHeB8n32jD8McsHdS8ag9U4fWyR
ik0sgt6+xwn0flfU45HKw4D07t7S8EGXf6F7sVQXTyQAFOoaiawYUnH+e09eIojN8gOdtMyQG1ma
hYzoO1CbWs1b9qQ63k1qv/cZKENhKdkxngjXV0AIy94LyQp4ZwwoHwcTzrxitVqc7yyZ0Rqr0R0b
BWboksYPD5xwYrfITfzSeB0bSBnQMGWNW6tBh544iH1lfc4v33DODJJB08XTpconMCBU4yFGJvLB
xe5sEwTW1vnkVphkySwShOfqnHFv5yPt0M8kcaOp8Gzr5YyKVwaFJYbVc2DnOzDNux6B61RCkAj7
JgamSXMkW19VKrYcaGymf6PrPn/52crrd0RgpF5uBoDt9+naPnqGHQ8td+V8YOQ6s/5MLiCm4rpY
B6BlJeKT9flwAHx06X5SoMkyU6VsQtK+TlLdnSsK07+gIENUQi1HDGa17uD0TZRjc0nUMGm+Hqea
uuSSXrc9tNYqEioy8vR0EAVk58/sqpE9w3VLkCF5EeDvYt7j+xZ4ieevKAOF1Y+TA6Ibf7vgtOoK
nKOEsfoKjaNO1A5zc/cVA88gFJAavShxN7491ke5Dqv72S7Ud6Qt9URFMRkOKzO7fTZl2RMj/2is
aVQBGsbV6cWA3bSa3Ha/tBTG9oacOMSeoVtvFUHHXXpO1RtOtQLJJYPGlO6ePJ+AAtKRjFFYIkfs
Z9QPOMj2edNrmxglVOE/CDmM6yBn1NblIInFn38fJeiW8lawwkSAJ1+/wO0sAqlgDTwmiXhieEKS
KsFXxSxOG4Eaz+5O7bBfxyFguqg616s+TCpYpvSLeG73S7RVTiqUmbHTE6PEUZWvQyuhoemYMXlN
R61ZCWqY1ncQounXKOKgsTPrmPWHvymCgey9YkqMMtIZgkiyGuFT+y0+Mtx8SxmBqhllaa57K9hL
4/ByoM7osNAjYknsDSYT1KpMINb7SStRZweIZshZ5QgEURB26x7BndJsXakPfDjgEWh2tmDKybn6
Jw/7Isr/MuVx8ZVmeGE62U0WWzxeOsgsOI3PQymC5UAsHEBlFwNzgrcqD2dF0owsAM3WTqpWO9iU
9v7qGy9+PamKppwfq95P2xoNuKTKhpD2A18wJC3uT63tjcfr2bs5+kT8loZn0Dti83L2pVHLKnLB
xPUSTtQufxIDpLid4OLO1UmdA6FUltTvDHTNYBHmUT68ZvNjXQwO0mRnyTjquJ2uiMjcvZBta2Aj
OOZn9BEvvg5IP8BBqRnRfABKDqp+vnQGB5p5D1SYrjSqe3VAtavGI7KHPkNGvQ8t0TMMyNMvr5H/
xiy3K/9xhf5Rnth4B9boH6UMtxrmnOQ5iy0KczXVbFlonQinnenljBMQy7TR5eVeEUbD3zn3Sh8+
IF6Ab6jxoU4jMBQJdQaAa0rhIzuX11sG2TA2YeYWanzyYk5j+5O3JbooQ7kSjfM8oIfULlj+Lh1+
jCqPKLDUlnWz+ACbUIas33Iavvpm+FcKKkB+OuyeNcZWC2N1YxasIkN9zerVUA2XoPmKlCaJkt7E
Ph0zuvqO/+M8GrOxaG+FELHsRWupvNYEJS5v7qy1n07EbsJvtCzuhDBz2Prdvwh1HVb7HhljHyLN
R7sPCSQ4K0kSeg6Vc3WJym9U0vFxX9FfhP592Cu7l0AXUXgXh+7JXeb0j/iXMw3R5a2oT/mrMMTV
zUrBKVNHQBtnaK0SjOZBa+29f8xzvHERfFajGVf4sqeOvKc1ITh+Si5V2Cyz2q1ipwbR4js2C30O
6SWpoBQLMxFQDGi5qRJ6xBrEE67fgeuA44zij5LDV4OmXDb4eHsu4q/zISG03R3BWyWRhK7vbfKZ
mZVZl/UINwIV4k+aghis2sC7FV3RIIxorBdUXqLiuCxW6Ky4KRQcN3VRbnJKDFbTC8v2k5OBj75S
bjqxbTjtD2oD6PvUFKDLH41P6fGXLPlDGTbmsZ07AfM3rmpzk1d4N5J3Ctl5uOjBqHTP1jYhjvTC
XVuZwIgMiMgXob/nxOa/yaYyQXgxoYHjphQSJGkZIdjfA1ypZ7H2+ztx0KwxVMr53GVw1A5xJanq
RNA1ZUmv93Sa/GcwMOmh1v94ioO8ulBtkNnkHrn7gN4x2bz0HsIXfIa2ZzmWjVcT1IZnWbaByccs
u41sucZSm5rWPAhTpgh6FLrMEHBXUuuDRjASffgykolv13mqkTj14a5oEVPgiu3uFonVcBHi18Yn
/uXi08X/4LvymkfhFJq5JtOw7aey6aVKZAUaxJRVvVnzr7ou7u1y9CRem4MAErYKedJ3g+R2jhTy
hpD4JxVnHotJ/Qzfq/JH+JJKjyfmmt75VVEdwByzFGGs6jq8BXWy1YbINsFwIed0Um0LeV3eAQ7R
Pd5v9r9riuctpJzyQRW1GxOVX5ld3wBN7Lili01ADumU+yauojeHDlJKsqsnQepiiKC3Y2ap9zSL
4g4vgrw/UUgNC+EPtkSXQtm1BcHAc3fy3vShQCpodJK1TYlWK43Sg/qq/eVZr6SVZgYKb6wmAW++
J5RBabvAnRqvF0DzhWyG5xBleFqMQgx5wQwXLZFXLW7w121G5QkQHGeEfRARZlesfvW/ZMNN2C2r
Fkz743rjTJWgjgDK74Nhk7/Sb2/AR/0mHy9KzKqyzcwFiwDf7HzzJCAznKARf5fLK9q5FTUH/ovG
RpPoFPA6ygcdPvozRLnPUDLrQdAPP32aS3eiczKQrmadA5iJEPHuLMW2EC8z23ZFAx9Rh8slkKuY
3Y4X/RFSaVOrKlHrXlQtOLg5/WvPMZtgGAf7ur6GF1eN6Nn38/AWDyw1epLWWN1U6e/BhygAYPUS
gsARS7K72L5iYYs5KhXEdgJ1vHuhmSXUPu9ofx91j3JEyhmUNlfOCNt6fqoX4G+6sU4hX3JdZGBQ
s/9VhUeRS7o9GJK61KCCkz/hl8MQCSxlbjYgwW6pIc7NA5zxLhgEDpTXJKVk8Zqm5I3zN3JB94kL
AmQNXUKJQD0iwiHvCmQmEhV53nEDGQcdDMDlMNJD03PsHEP6OR0kecVuZDIlgYK55kmFgzRkobSr
4PsNn/mUCGH17lvmwdAwuzHzCSz0pwSVqzGk8q6E0q53SIJCG1EVvIRCdKoYbt056ocQgMezLKmv
RAWH2oTz8+VXCYChdSHPf7HjpC9hdiGHNdrFKicRHBAm1g3X46dQxdhvbKr6rniNenuyPmqtBkzk
DBKa1ZH8YkgASlcX641L/JM/NGdagO0tSG0T+Io9Cm1G0CSC9kOD/NeUiOnsaMBFoawMWxgUezkw
kAgJhbR2AidrBqPujroFckQJ+6SbQGrtNe/fdBIhqsQhBBlgk1NpUr38rPbsWLD65B7B7QkwO2cM
XtnBu5qDpAtqr6ckC7cU+ndIOqirfKrOpLhXtlUFw5F6U3WVgbOnHRXo3BtE2QbJEfAmKJVdxslv
VeyHKHf11b8xVKh1offwCK9yfvaiXohRYyDZWsQQ2sN4uvzMD0pu0JtBjQXtjFrlF3iELksLELzf
17ujfk0JPvEyYlj2UXcY28L43QEDIBxqIJBASQcJNNCYOpEMTa1+PuWq5UEEGpdK9iAstaP0qT8X
nyoYrl0h/Fz2B9MncHVRYiptNRA/ihqe+2g3ziomhihLph/y8dwP4u5y++VVCjIG7JhQgW4mlR+4
pDVI7k0J4B3enmUzPO6tVU6gxxt02Yo2qOv5kjAn6Dd9cDtL7eNrF0ljcjLVb3XCWD75GPvZsERs
zZM2pfzu6Ya5VAhLEDIDfVXJ4xV6GamOAzh7osAD3wKKUBpevp1GgSObqkYtRdIkdg95fKRP+l5U
KEDBqmj7GBQd9k953T46LQB2yJk+X5549zGJT2vgkNbsW0KK9AnH6x+++xOCeBGQOOSW1bbnKFbb
uYIMZZtQfZgMqSINpJoP5GewNB914U2t8KFAtSWVc7XmLmkxJ0gIgazgCsWxruCnOsnvfcBxjvDM
wO2EpZgkxlhFUxd3QsGudXNUZPx+l9QCMaC3jCRxiH63Zr1pEpldbaXyxmRlTmtLwb8rAKmhcKI7
NHeyIxxgnA2obNk4yqGqx/gKwhlKpBeCWAzRmn9zpSwx1pkTBU2pIHq6qSVK3fuViZ9bAr5di4Va
5UykNlLFS8tiTmCz7wsB/14J3osbLiSOXrUnsaeaWJNGOqN8q3JHHEkuLeP+1IohEutj+9I9UBRu
JhSfB0eXHzuptqE1FzpK4kTP4yGJBXlAy2WR8LHfycBUEAgd37TIxyzOcmKa8+ILMOd1GzBC8LFy
x9WG/X4xINB+QbLBXkprZlauJzknVCIpVQqBuO+e5Uyw/ek4M+y5oCyo6j4fRCs4tC0vMPWKenl1
odhO2FYcuH21RIJ29GRr5TNDnqUFg2EebRNUbc9+NzsZuwx/b5hL1qPEI3yR8Uf0P0xJDGMlMHRS
F3Z4F5GPpbEZwr2gWnjT07gKV8esIhr04AfFgbIVYoWK3k9maEZFWrkx65yC0kFhaSJ42VQqmoPq
P06x80RXkmkgFoejIwu5Er4zoD83aOulklWTNuy1xpu9zurTZpVhCxl3GHbwNC+mOFMLLW3pwFjR
jnffrc8s6Q9U7TTVE5CBjDcN4fc4giFrGjvsJsDVIqe2bvMRjVoSieIjtdVJLX2QqDafiwQRaKyF
/bRppCi8euN0rnwfTwfKdn+v9uoU03gBev0idNOf4Wqj6QFhx/FtpJmP1piswUBAt67pZbwXhMhk
gRoNoO2GVIf3GE23Q06IrtYiNZDkAdJYJdUih1A0CQ0NMyMpMcb5gpRWUmPX54qVDXvEqyigFqb2
R7V1YDNpbTlEsY22pp26i5rIlIxPO+Ii7eIx9VhjzNYIzHgmJS8eChqpfU9tdGZNPdV208INvXQI
JBnx8hJxN3zFqGb+SQrPK2fvMUtoc8sc7wiFxZGsUtHNvw6ArQ2Z3s2IppMLfFHiQXMYMgB92cCj
65o+oV/BkiLz97Ohx/qHrwWu7vrPntFUnZtpaRdbPnSmjwmke8KrsShAzoGbL22TjTfvFdQvmfZv
4BDPS4d2SyVtkg8AaisGmP7AwU3N1FAYWJunpZfGsFLJQsDrpOfUfUS/Bqza4/u0Btu/9duy/Gky
TzUkFJRXz2gHafe+jvgaJahtwV7N7AKUoZvUt5yBh/D6iT6U4w7CprIu9WOhGHKdhh/jLf4plw8+
yWg6lk2eBD7c14dyRk0Vc3ahg3cUPmHB2PP7u796VaKS5NhlStM+ec/kVHb0QaVJWS61s0h+YaLv
773HTxpk58U9GQFPL7rxJ5pzMgUB2jZ2IkIZlt/BzKAsKVmvG0+ave6Tqh9LZkxt14AZ+Lpgx1ef
Q+ZDTffyoqxB+84P4dtM7yM+wz0/5mrea1DPjLPKFwOPHITQI4JVcaiq2Za0WxVCnEzYhFr5LHSZ
N7V2YKInzWd6W/FS+eYfKGImG99qt0GTV/eXuHWJABISiKSUy/9j4YiVBSWWkXBGOr+NGekGRzdR
yKONTz012gT7uiSZKFyJjpTmK3S1MnP8/vZCNMAtdyhpgNSJwp6gf0TZ1OydBUqQEYdi0ULrU2Ld
0pq/uYlSow2d02XZNfYAyqZ8NiRmwvOOG1vn6pP/qTVcSzHYhTz+iHAxQnxQJsipxh/MBkwRuzwB
GpkGEKLvaZzP9fcnTKHEO6MoIVl5VeR8532lGjnEpLCxLL2mEQ2Uo0EF/ZdoTLhSr3gRtK3zRVQd
+uux/pP7PeYHyVd2dHWo3yavMcQGYjCY5uz8gFmFnH3IJzxrrlzUeZzf9jRPIK0sFMLFEJKwpwpG
KFOmWvqTmF0223rj40Eey9KbHfKE0Tt31hk6sCSumjmllG0717ZBD1Dtc0YbF3vXOckQ2ZXktD/D
GztIn8rLrpQlmlVeXhMRmW4Qrf5iNsLShxZbmEEW7svf8iHtFbp3Amvap0fV/s3+m8w9AgA/NJFL
G9A6FzM4jiHiIw2I4CnMyeP5dR4+cKVC08czvZe6PHv8WBlUeQ6O/ig9ub6/XqRs71ahfQd/umAa
Scw6l2TNK/Wj0BKt3BijMz8iL7cKoj6fP7LhToId1KmJV34d6Hd3EghpwgNdfGGPJ5g2V2GzNHNz
B9Y2OdKoBYMMOGjbwRBwdVXV2qOBbythggMDQiD87u8IZSfmDUN6NOW993KtEUjURLd7CUg39v0E
xJcOhC8o2HJx9gQMjKKN/W8Qr1v3lgXMSL4knBMcThsLI2ygxr+flrzB5QnmEVo1MK9HP2g6EhWQ
jllaCjz3Q8NXNUy0QBMsP2Z/+yR4pAdmR5GV1XZMo5E2jR6fytoQzzXPMlB7bfEe/ktcWHX+EUBP
TVytWNg6mpkzBitslQem4ipQCafeN8pJ5cCHsPxhDUxxe5ofVwlZ5EdGppOAXVpQE6b6caXm6pgQ
YsrU3Ehfcf10++6KWBTGDmgr1+pVoGQEP+KcgcAxFEUqSePl6Fp+czh36b7HKkEYOebIFhThpblS
vsiYamSJVw48r1XVMyCktLF35oRvWuazLnQUWgWvUzKJLIqlObU31RRuvQTSxbPP+NVm8gFqMKVK
GyDHAHoL4f+FcdvaSTufrknRItOFgc6eY4ioJVf6R7Mu4Ypu3metmBdphsa6dd3OepRGko30uTuV
M3hCMFK6yR2Gn+geNaIU71i2qvht9kq2C8EAy+yZTQmM1d4yFLNhGdc/FjQG/+wSVYAbtdoAGCDW
HXdppNHh9Ay9VJ4hm5eIN+s4nb/bzOJ7LTIZIrRuM9lRQ3mv6BsoO4rOfjCxLAPDUqmRcYfheXkq
P+Re/IMC/UHFy5oP1kHs3de6SG+n4HSzQe6swidYLDMrad1uBtyNlyMjrWGlzS0TzNSc4hVDgzaW
JfkIpGIZvQfmoIhdV3BtQeuZTx9/8Ymautx8FCXC6ZHk3myevwuI134uJke437xxLGFfcJ2+poFZ
BI/MUfuozmhzPwh3xslZCCbnh6tkzyR9wl+HGQXcj5fyQJEsBRO5qBx6+L0cTNjnjrK+LFfhG8dT
fXP2rOnnErI+YqWB0v4GjL57rjpwgsc9iLQ90mENlmk+Bs1t2Nc364XRN0qcGR0Cbd6rB6OHvzY1
pH72QlM/UEGFwVfahN5ocOFoprvxNaTKxOrcetP2938JNhK7S4PE0TEbh/e7mEpgNxCoEtjSGrWu
qDnuw8+ytA+gdsg02cJD7MkEV8KCkO/uJV9unpHthgOFz3e3+BPqe/JamMCNvr8GvMvEEfxbM59d
BAf01vlNKh2/wQX8qExgMCUATlsQWTWFoxYf5xBiBCJLVmvNO0RrkCOnPkrfp+KNf/byb2wINZCv
1Hfl5Gvpeh5kifyAifOdFXFxrc8dFXe8cTySvsRqPIoMKuayUl+TdfJvKtxlTusAPs6O5YwYWug/
TpeDe0IVYHdXj7s8mhFbIGlXHgLK2NGmeW7e+hQxHuGCnwjLmJ2Beaw18O86tnHbm8b2ZGgVNdcU
eWuowuI7umljMB8iT9K0jn+a2sHlQTaq6IYV1+jQ6kydFLBMhkSKBCV/ASmIu6CMCPevVCZGuod4
dJ49EGRWVGPtt7CwTbfNng/OPhCOXb28zL/1nFdBWsCbnD0MatT5FgVNEBQyc0GTKAnqVgOJV8Yh
I9BJ9AgdpWk5ncFdx3xGx/yWp0Kqi6ljJvw/HApZvO7ceB/IF175rsx95IuiyZrYSniig1/7CZsc
/nqda+y6cfmkCsbDz4m7Q5sLyTBnHwnildepvNv4qFQArSt69lB5dmItWMJXRwmjdPZy5mkjY19g
7/5hyX7LPeoPKtAlQowsQOc0Z6F2h+JtoXomaMmZMSNfdv1ijKOn6ev3FcJXFfrc8Vi6xxnErgEE
27ZbfPh2eUjRIzRpGUKLNf5vGPSHp0FXExEhA9qFRiRmPxCfQuHJ/kQbLmSzlbq7YnnTcLar75hB
WtDofdSkmulJWOyfFzp0u+TdmQnq6uBimlwBOkheoykR3rWKScsDolV2eW3ZuZGQzsxlb3CqAVqv
fBoc0yybYntSlP6AQjrnFTcnOSX+UEyLPlN1jXaaaDviHZJCl1J6u523kzCeZkuw2XDztX5j5Mp9
3ZzSF6eoa+PNc0CXTAd6MPMBmQuOEmg835PYMKLsLn7HciUbzLQSo7BW9JwnAVU8l9CSTs+bgWeQ
dkTvbQMIVugrYjeLt+uSIQsvKlovBfnT0DPXqMqwwN0CsNtU1I/FTW9rv7Xm1A+r78n6roR8q7gf
1+9FTzAUsA21r7Uo67hsKqtSlp0keU0TjVp6H7kFJ0D3Ef6pyZZB0bZEfVMbytkcZaKJUJ+KFh/9
n6SX/jHP5Gm8SgoFblnO6oKxXlPoGMViJB+jdoJWB2CshD3C0VoFrq3hPbnsl3UMFssvO/DewBIW
N5hSC9VZAhFPbIjPYF5tayEIH3dXg6rQCxvuXfT9Y1/4glUt4Ndju9/OzUoUboJwXQgoGzmsBN6v
Tx0p7fKkqrtz81XTPMixig3HOInrmh08yKf0Tq5N2h3dQfxWoaOcRMybI6PHOsxfUkHRbrR7IYqC
N0Oxy3NU6C6/MyPtZxWTSoRqxiFCpuffppynMUPp60OLB33zjX7Gs5z+m615+kjGfrGIxXAQ7Pfz
1RHTKnftvIVWUi7tVfo5cul3sr+9UIrZ8Vh7A3shJlIsLTBuy+p8JGpjR2pLVN16+KFp2il7joxH
BU2mK1MXk410yvt72Na9j8e0R46kfgm+I76S0j9qUsh+zAri7F4XhQnx43HqOAhmv3MehVldDF/6
JoQ5w9mnQGONMJ5l0GclEJ/GkhLNc8wdR9OjWfT2+j97bohtTwzaFCEK8kneVowXWks7uqYxCb3s
B2yHSExBwMaPRex57mXqsn6P0hj+nIJ1bvv7gHta+jkdanZZyc85Xf9KnBzLUMoNrxdc/liF431W
DDTnb1Zc2LVdGV6RkT33Uo9JzxhbuaaZjA/4Lr/DdqcNSw2dVmnczGQ6xSHsWKN3yfAfGPPB9JGp
Vo361f1Rpj02IScyawzqFUru0q2zVnOr+Er1uKu/bSwKcCbE9ZCgG31YYlsdyGofiaVwExjc6jMV
8HBHclVXYkG6Q5D3a9KJ2MHwp97TyE/Ei/sNF2qq79Xl2kivS/GxOQ2wPSkf6tCLuxLCgCvisFp2
KbxAaMxW7eRCpeC+ih4eXfUduCvf9EtrTatwo5xjwI6l/vbnjKjtCePpYds/5So/HsilufkWTGHI
Uyf28jbQxoWOCegOdMGiT3FofFS9w0AtPBIo3Wu/znJwqwDLq33uJlnKOSc9a/D7KgwRJ5tuorYD
vpM42ujsUrfA6Oehr+t5jjnFC9HojU0KM5TH6KQk5NE/cMmLUhBL07KyfSb26l5FT2BoybzyCMP9
K4gzf6oXFY5iNPq69VyoztSepR8UzH/Us2jwqqySDEsu+rid+dDKX1xCxKNzYe+Gs0gB+mGUUcl7
ZkK44yssoUxSlUx5m/cTLIJVT+kzvLIc+EMZv5F9Tpu8bKOXXsZsKtLOvZBESJULv/KvLG7ShACr
ElBS0mXFt75IupGaAB1L/pCbbEfb+jb4pFW7R72zCdsIaP4VjdtpDRnFVj3wzNXLVPrQNYbirF4n
15lpFJQ8mgg34GLX6uIrscpMwlcg2Dxrlw3BNo6CLP0f6kmRp+YaHDaMcgswz9OprMcvs+l+iYKi
2fhZzAJtKLbUJ/d7LFpc7sjx/P0iJ2dbj0vHfnLAzqURGVcDXEczK6IiK9qSI9ciCZoXIgo9sLUN
cB3Ce0Z+3urt86KRzl7/V9ob0De2uECYfJNElCnpDazK1YNZlVDciUAwooba8LAUijpE4Nz+4VtM
1LHtOd2RCgMEBVXZhZ6o/Yt3anDJtf65a46Z0FzO8ituzKXxGzmys57PAEDfb8/Fo979JVS4Ikzd
tzsdC7MyeQ3fRyulg1jBdKmzEEjOcNnyNkQs/lzXbmHszGDNbSCpFCHrQKjoripY+FoudaJjhXAb
HDSnqX/+QUXh4NJWUnLjvNL7e/KTRvrJss6RM9cHq8ALhCcSN8dD9eUQZh+v7sHuEuincoBua3Ah
4XpVOYHivD0yb/krImemI02I24TlBAq1gAcYwuu8qCTYphP/HRL1uu6uld0PWkcY7fp0PC9FBgDD
0YAjvw9XDFUGHTIsbNpZi2LWl7ZGbNzgGzxvC6US4Fdoj7GqABkUj7Byx3jEtVUUrGNqqDFNuV+G
M9TVeHzWSCgdqGGaAHoqvfWMH3PTRo+ERmUH69GM9vFG6ME9jyN6he/fPeHxzMCTCuhLq4inNdap
4DTraUay6RG27fSelcp1jedi3J6BBdNcn20c3ofjdJi1BYzS4bNkaylTesE9fTg2u3+ew4/smXFi
kQM8rofle77VZ8MvtDkjulm8GBV3gcSnXWppdKnRkGza5s8y+zss3FK/2ZKIMqV+GFi5jZRZ+vEq
o25Tx9EmIzCvnRkQeQftAYOcje581bHfqIUdnWuFPh79OxzYHjofp/461HfgDy/RZhOY7HxgmxUK
N77v8w6VZST1e2t7wz+V8IDSBRQJBg6T0I1op6Tk7Fj6fKjdXcWIKlaArp/dMj4+/GimHJysyZUd
V4TjsnBwxUV9zh3LwRl2MlYE19tMD7kpVqgCukCXxFxLG7rRLFp5E7ZMagyICkdX50bL2iRP1dqf
7pPSgL8W5hZx4D4suP/G/qUliF+EXsT1xmv3PcPOUX7kq/1YFKefMn8j2wPdXpnmZDoPdieOIwMn
c7mjziiRDUVS6CtYm5WaYxKgdc2mwWzSCawDSVNBe5miTwEEaW7yRroZ99VE3sIzJQZ+ZZY8AnZn
bH5B9Lx607ZNgpIvi5Cb94oJU8SxtEFrqsQbac3nN3nlAc/juVSBL+suzuvNS7rqETC2Yp4X5DVA
SdTyefeuXxboyEaUMjSPcpGtzgOqjNQUhUuT692+QWZNuPjDuKYKyDN0tX5kiDtt4MZQZjUGe27u
x9ISth/SE6QNo8BAYGg++mp6mE/CSGk/xuV9r8REWkMjUdXsv+8x0aoH8ODSF/S/fTO7JyF3C/q1
9aq6PA/Sv22FiKkbYeIfIMENj31jBXsUOLCOCjdacSI9Ya3ZnW/DYfUqgARgSgFfcRt8/uboGEx4
wOMz/xyy1hvsn5eb9rusHZSpp2tcMs2GwDFI6oHtmZGG2FFxPrhA+GzHVWX15vFLFYAQ/WPm1u20
Dh2Q7c8iUeIy64pid3oUUSFxMFKeEiGGDHuD1H84lL93EGi06JpA2opMjCThhNP8JA/yIFZZ86A/
KcqyVKUUDS9MPD0D+k5gM81bQhggOVhG5FqOQEYePqEZj16xkZu9dUVmtqoS+21JYE4BGiIpS2cK
v8yqC8/c2rX85IkKulGYkkQ8LFu6ujT52wqUHLWWAgRbD5F5534eIqr7UyHnULZmpBbMw6ZtJaU1
zns8YDH3EC8IshKvwl94ZstUmGr+nzpFhdQfJ/guurrTVrneHOUiDjX1evKRvAIrCRBtTmBCowzd
v74yK/mdw2Xi2D7CraV/1IKu0i6kKq9bV/JMHLV5PGUuUNPFhDpieIYa7KLURtBKekbZlp1D4m+T
OTThAFp8QzmuZCNvghwvAmc7dzzkzq/SL/oT7M2AZG21f+PViPJd5uL9iKfIOivAtvbpOH0yjcRv
Qwjs6u5+zRShZkC58lvvrXyp4dPXdAYvdXBDivPw5EZq3aiSkEwCwqdY7ea8CF0uImH8rvCzb3hB
GwJBzPIZMyw4YulTELJ1HEM3Il+cFga7hP9XA66Ck0rNaNHq2xSguwMfKFNWO9NifqkkTdB47QP9
xdq/puh8TFTUw4irrQZ9uAAaoLdNzP7CcemLN/NjA5jWWTwy1lvttZjtPDu67zz8GkWD3CzjwNOL
YOrIXOsJHcRLq/zockfuar4M+Ys+98RJQ8lfhlWBzsXwcHkftUabDHN2u6CyHCEgGQNazzV207HP
4Y2vj8QQabXz+iuWY7OP2s91w9bggmm6iB2DBMxxxnofgBooTjDTXLq4MebJqJmVP1yo79rH4PYb
4B/n2Y8bjSx7h3gB2y/bVeJRW+xQ3yK2dFBRwS6+KSpmmCxX7yoX8aHKDa2gpz0LHwfTP7PhJW9X
/gzLe0OFgHomn0gRVofojUG1CWOaGJuf7w9t9RFP/1t6/jRqWLxroDKxjZUL3kdom1dVhEVHr5TE
E1awtGuhEZuxltyIlnClW2gaO2LlvKNrW+feyyLFiKQ0RxKFdzM7M07b3ChkZLLbiP11gUY0vfP5
RTxuM+QhajT7Q2Gch7/T1l3s3FYjnxXQ/LqTUaKpWtMVTxOPjEtU40zJ5/Cmo6IhbwzGHJWN1cqM
G3F3UY7dyftG5MPcSVRRWd724ONHUQtdIRXWbhi8x45LjaWboQ9VArhYYUR8xfqV8fgJkcy1z1yd
1s0WHnCZLQg+DdB/3XbThLTUQMyFgbH8lS8di0H4pXM+S0InXQtkNO2aJypumWhtEP0fSVUrXyTN
PhQXx5cDaKcG2gVDkpD7bNzw/GIRe4iiywnQgY2Gk7ldiZoPzIbG+yppzi//9jGWFFJ4/lLTpyxU
nYZirIyurtQWXlI44gEdg0eTf9/7rrjRaqcy6G+NEft6KIpzruWDR83twKriHUdk7+dUlnRIB4Ai
q6va349pihyNT+aaDb5BKrzYvE0RQN04bSHQAa/ppt62/yFjoARFACk2cWBGp55dzs9WjbzmgATG
TOywVraLjegiIGq70BY3GWI+dM7KUt6OLxlfc6sMuifQv4KERpx4/wAbB3ZobJGWSkOPIJKGrRnf
riE8tkgxahUvaVSQRoc7ceZTX9KFCaqEq187kWRPSsNr6Jn05XjB4XEyKR1nTmPK0n/IBL95/53K
X8wbPStKeZSw/xCps4OVAPsblKiH0eo4y/iXBG9MlGSYot14tY3vkNPrOmHsrUKR4OurSWGcFOtR
DEZ7WZpcDCvSRHStvrkFUg0Jz+eCGd9xxc7sMkLPsoKB4PChR9mRXriwflFiKZ4d+ar6G9bcUcy3
XHjGJJedIqDbPrtdCEGsC6n8aLkhubJCedugW4KnOEyA8AwTckPlMOseOMHBWzsdwZ2qgaK/YYkl
hDYdELQfNcUTaxEa78+qh5yuiowYSBuYpDWGvCrOFGboJnq6rj8O3JnAzabLFJbghcEDyS0bzyaX
kJOTKG9Y5w6IyfQfJkpuKCZt/sZ1INovh4Swwr2LTkgzOqBjRA39xmXuB0hNzibAxclFHHZ0RHw6
rdeL5XQrruxGqhcXAufsocCUtX6imZydzDNDdBTNSN7hWUBDEAvZ5YL+v80JLZLd0aL8bESfHzXO
5R/HMGqRZ+pPm4m5VmwcQGgc72Hj6Nu4txj8vKUJegoO8M4+71DC54MpYA+MYenBIZ+UntFpMpWt
POmuIIKht3Etf8bByEcnKHbSc5hIgLCFlK/QUuzIY2RekH3u7/desUkvNEh8iOtU72DYBSy4WlUQ
WPya7Mj/r9JCRwHM1hI8Rz9EJ9ZJVtqDq+eXsjdAD/FOs/6hDCJUghzTEwo2o8DWlIG3vRFP7oyO
m5b6LM2WAqM9q562d0uFg1b3QxdjLq4yzkm1tlbb9zckN8Yt+NfXQrcNOkWNFrGq56Mv59v80TjG
K3l8KJIMQPppysqSOpVx+IP9vFEZHBOFqWNRyCUk/8H2KRrmUQc2R2k1i6QY3gOnJeTR1CxZiKjj
Z6vq3uihmrzqNtiqplWtuSRsbnYcW9/LJCChE/PV8NMfo2LepacghRtBNIxMxZ0z3my8ZYrL7cfL
S0OWmPW6/KondBYANU4NtMsd6BxiHXE5FrBerdQxRaYYKOKrdoHWek0KWzzKT3qKuF0gA03y6Nyy
YPcc1g8CSef/eYbqSMElljUVvvb963V0wbosuTSbKaI71dvdB1tsbsUZbBi6G1lRXKIXWrkssuB2
ybyubCCvV8/16KmK4RlnJMXykCjn3O/2ehWN6a13+b2kVl5ktukMkp2pwv4bLl6y4aze1uou0EcJ
IhdJSR6Yz10Z3mJW6+p6Aj+ccWUQlCYsbfhlrbion0d81en5tHjfygEeTA/k3zHUZ8gKrIHdY/mS
TbuHUDKjGfD+WHY7eLV3YPU9+0pZE1qEF/LX0/gjOgQyo7mjEJYush/3i/5lIrvIStYda1gHhsZ6
vs9aVJVTMjhg/FV2QoHIydibqN2m/w2XyvbGYSuKQOzQS3bvsVXGxkzZtzJTYfnJZauRW0ohDt7U
scqE7F8BOozspV3RibL9RGzdyNMTuz6J5//nV9+HgEK1FV9PkmG+5f50ZAgsEvGFm4KUHE0bKOMH
seFSINrkhYD1xssNHLYMAbBuz2377gbOW1xoS1DqpOC7Eh7gD8vDat2WSHtxTcsJP26Qcqs1b2g7
uD8nvFuj3zF941xe3Zdtw35olIlNAmXatfUnfgbQCBm0QvgyaS27B1oafgtmnu9UBdYpbRwKwQMA
gW2n89GtneBGHJuH2eFOvVqHD29/KAyzckrKVEElXgKcG11aOkUuHWESQoBd1KArChqIgOmr6/tW
wAwagGkbw+vFbC5L65d3naKui0zGZWDHHhXTJe7imYM+lbpCZ9yZCN9Wp9pzb9xewLQvFzdEExwJ
6dPWVgsDMdNt7qhw7SXKBWuqcgr5bBJaeFLTEgWfBM3T3dwSxre9esb36/0MFkGgutu5G6L6ib9q
kJQtmF1iOvOXbChFT93LDqUogoibbk9B5Zrwpipt7S0HmQeHINB9NGlF+MnwICRJZsl4YmDnrMBG
UTDw1jTjrdUanlNEkRrXBcSB0s1uAY10WhPGEjALjr9deP79nXMhfSeEhQzdcf7lykNN3QdDVvsm
O+Yxe0HSb5C5452mbTjDikSkca52wbxoVIEcyqF9Goel/VU+7aQlpJi4xc4sn02+BGDy5eoN5DD2
IS2vdGpFuzzJnhAfXDNq9h/sm2QDWMaG4tBS0nHPpWgqK4TkYFm3p+/FUpwDbwI+h3RzxCQ5hDcB
/hc5U4dsgZO0r0rU/+T2oRCBfhg3L5aKCxiSV9tnGeECOiBQcV9cwn8dzdpW88Z59OHRunu+M8xr
pCNrXOEdUnuxJFqonqIwR/zZiFXmVyanoLu9bheF6C+3n5/pPhiDlmUD+B3tVDtSbgDKKoJNI4bb
Pw4tjRV2AafOcQNx9jWTeBQt5/Pn4iuxHMfiR/jmblHI/2Dk1xs3Wm6arUSF4SLTkjAjL+rolI9l
WIQ65omvdl5hss/famft1CdylkSaTLfmelP2mWQEtbtbtcYCSskuIhpix2IZaCra3PifT1dw+AAN
oKPETnfQ6kWE46pSjvOLVGlzipaHcWTbnDTRJMfpDHyhq9hAvGNNmetQTdOcAm7gkDzqHqCibwKD
ls6jBexDBVwn5Up8nIWmdPFAJcSoGRxBVpUgf/VKrucYQkDrj/IC/KFI3Tvc3xCAt2/poPYiz7go
0O3M3qdgSK5AaZThuWxbzQEQtg+ezQ1z+YW2mQpxT+qGiN76xsmP6APWysxHS001rSEtpaPdyIQd
hrbPM8kB8qtVDVnQ8Mn6V7snA7P+7JjwQbRqpzUftZR8G8Ez73nsydUiOS5dQ5KuozXZRHfwnC74
XLX8mpOj4VsO1jRQoEsxW9/S8B085YGku4srS+qYbbJcx9U/XAbnrRZP2lU5g+SK9aUvt91S5xn1
3UIa04urB9F0C+eWMPQCQbzhymDAvUIoGAB+K3P+mV8uGCy6+9RyzFZ4yuqE/a/cwnEsfJqOrDSH
gt/GAduKE9TMyIRG8kwJoUMyJ++GV5LkGbVFX0hwnowMbWO02gjb5shcSIBGN9YZTTIBmyEICq4M
M0fCocpE6dhFRZ4Ib8gURzum4/kE4VueeioC3ebNysyzzgztecuurkQLX3qZ79YEOI2139ZEkHTN
oQxDN0P3HeVA1NXhjOCArXoM3PZn8/lLpDgHjL3Z9CvCH3C6czKK//H5CNPVAiEOWo6LeCPKnGfQ
8i+CV9G0kXQ9FlOvofItPJfcqipCuA9VAjXP88f6VJK/b+7od+MDDqDV74mu/92tJKHYZTLtO6M5
jgtpa+dD+X+L99VW1pc6VeVkMiyCLO197SuOp2UvUiV7A5NS3333cxnO6PtjSVhxtO9TKphbrHsz
jRZmhsXmQVgALH/JH1OtJd6QrPQcv+kPZ3v2ntmDZMfHCkUZURpdTo4NM+yfZwBqQJ+Y5DuW3jvf
1XyWBwSpu6DWbRlUajF6tvpvRXtBVUByuq98G9BxFSBx5WugLXnME5lJ4bw8M2/mEEJ38W48SNPc
7ZpGJql5RfssRrYoltxzjf8nJB9oc+pzJ4WLuzpa+NEMzgrkDbx7sJ327jOFU8f7DXfRs9nHFQOn
WZrVWOZCoeUjrNs97nWaip4bJ+rLqYsxNDssVsYkK72JPDcO3uaSav7H8YIa6d+3+jd3YkZ9c+fn
wnR3qIdS6uCaaMWBzr2e8dSnQrm47IOwTVOtSTo9GyZVlz1yAnlRI4Hsp9rswBwxOCNWRIAYbPgl
uc2zUw2EephIKAL+EZPjd++xQ8YaXlPulqy3WjYzbwJh8tw4CUkw9JyEUkbfNBG83Jatovt/Hp/7
G9eB4uhyTPNvh1KTC17FPlZ5hDFcpBj9ufY5sn6dJgo3+qQsULPORZLnmJE9IQohBA0UJP/a4skX
m8H7FXdLB/gYN4MubPnqDM5EJWcKkaGDX8b1JYKYVG5LyyrCAwOeR7xaAW1yNihQzybcBeY7NVa1
e9ALG0+CxrXEtUR0kt5qnsVK8JwJQ/xJUBELjaw4ON4DpYEoYRtnUMach5n8e+Uu/q40OgpLZ54S
0vGR7yWtjKMz0lrq4OESqIFfYxAGtM0Kc/ctgeN1YVqfX0S7dY62A6+GNtNsSOj3Xk3VgxQ6b2uS
CnL7YTzBMw1Fs1GdX/5gjPgKDWfsM62Bhl8G6sZ85+6wJm0MR2squvkMB7DnhaMnpe0YUEfTKor7
Eummi9CgU1WS8T3ewviQHM+ciu1wJCxjN8jL+zBw1h7fNRMtneHxtNFWhyhRfvKS2gjKQ3RTc6a8
+0joiNePo826i92SvdqC4iXa8JNc8+REt02hqqFU0ytK5BiTRvDcG4xq+l6V6eSrDox0el4GehND
w3Hzo0fJZo/8x1mNWanQhtvhW1RVYV3GL+1srSIFojzW5wYspeEnLNNH/MQOD43SDM5j9ngAgGXw
c+RCCn9i+TByy2V7lA0ojNX9SzkRIm5OUZ85oLD2pPYpl745GnON3Y1aVHi0bi5a8scDoRIH8cKH
6lswR9E2gFEXqIPhHYbv07NCCYhPi9iG/NascajSskEBumEgGq9cxT8e6tLVxg5Hm4QqMvQTqaMI
P7pILsdGBejciAIsvKBVkjmT5DY0NpF38bj5OsZO86DNV4/YxUbMiSXKbZU2COX9Tg7jD+UnTYtk
6T8rsOyuHUHZCzUCV0UeiK6MJXH9Db8eaNOZeYvhb4Tb3OGFE3i9xG3EGGVX7NbMlJrmfBOPzzqo
BsYDq8NsreupyhjKLmYQxus4eSQFWF7JtfCPCC8SFVJkKFevb3mQ5ZpPj9kxJX2SkVZ2E+1L3biQ
b5W2tdySQvH+nPBxtGFY09stKBrO91NJOuugSW0kYYEkcvjMr+W2i7PTVxNn9UFgra47Vn5oj4wa
GBEU+hsWlp1CSHSMUtXLzfFUY3iGHZgMprcUuGWJOSYN4w0vfSJu55cL27qf+FoEi/fMVZGtyQ/M
7oz9VJiyKeSQwUEhNWB3+v26jsmPdPJ/ZsmXJx7hMOkUiN8KaWK4ohWGFjKm9QrKDi/pxy7AgpaB
bPSHEqlCdsWKdipEmh9U8ixhiTDMIgsGCIOZOSOklGQNXpmgSxjI8dk+vDp/E25mAGgMLGToapDQ
FGPv3OtsUjE9I8tfkSCP7WENSqHY9DDIFdm0l3US+BapRPWVe4Zp+uuPKVSUAdKmPAWsezWe4gjG
r+jXPr4spQqH7GXMV8JHYRh4vGRNwaDaLo4SyepgkIzanxn5/3RLuTaCMjA5aL8sup+LL1GHqB/2
vZcy2uSpPVaThgetlnO462wV2tI0q6Fy1ld+U8dTBfDp72AuKuTuTxNc4xgLYYS1EvskPWpfg/WC
Fwpu3Mh42VU1s3swf4mCkXefGX6qdpNNH9jtQnC44vhKzO7xqdw1oc0mjTA+5Xu60hO4WWBygFJS
g6m9k9wUbnmdFdpOleb6qhk5fJt5/3FlLVy8VglUe6kaMVBOAsusFT6titJs5EjOBiImehwr8xmz
JWNMBHHw6m5uAT8H+xPGzVkhdOM4Bw00yEtWAofUbQTlLw5gjCzL+PFpp8xE+o3G812qC4uTWSRX
YxWu6lC3GqJige+bGSFcYeLM6OZ7rQUJyt0l/LdZLNllIj7bJmsWsgcM5BdISx3HWGa9dUGSgXQj
I6im4GY6jamvNel7BfDYD/QWTEFq+5fB7+q7Dg1DEzyyd2rc+43xKZJOfQEwO3j5QEMOnz9INSn3
v8FcwypeSquozZNQpxaoKvKr7KJKjwWVquDBhHH0dZIwKiQWf2nKU3hBe6pcIQIvxs6vVFLV1KSm
v+LUDwfFXpYH6Rh46BO8msj4rAPy0zgUjM/YAOTkk7uL18mVrDNht3h4P9lPA3lHuiaj/tWXGphm
vSW8u4JbZxUSt3SD40R7sl40FvXcG9BN1DO1UIdd+P+ERId/v34a6c/Q7bi0fFJUbicVhja5/DWV
Qkvyv1wnek7Qjmm7AGn4Icov0r7X4uno/wdN3NiIwGWAEYE59pWIREhau44qmrtm4G1TY7GfI2GC
u4m0Y9OrBipU+YT1MaO42k31cYwR0+08ICQXrNNDJj2V1d1I/K+MXC8oLDu2ooUvTrmANSuwU5vC
xyVq3WiQRKKymil2w58cuT/PjNRlsFbgL1cDuUw3yoiyGnD1jJ8x0wS/AY3KqyYVHk231B6JCdY4
jCVJCWm4PVuu5DQckqn5g0iQHpE+lsZza5OwuJD+9z3xQEUFW8fU8rdMfMpQusZwzTRJsVlA75sw
/b9HG/R7foKkfaCKdTNQhDmC5tr+o6nsmKd1I2jdODBYrfpsgyWF7dOoUwUv1pvo1wW4Ibgw/+/C
Crd9nTkWmn4Q3iY4iQoj+aiG2dZk4y4LM1ECmexfbzs8nc0KterGpGhMKTMxocm3QdTl47LpxxhW
Z/aZ6TT5OWh/bPMKUhNEo/8aKLAEpR9DAfv7yKo3FYIHsWjUXxOeTBQ2SIqBiLhoesClyklvYbUZ
8OmpAZWV5XOvqSysPNCITNH/qp+/kqoP4BGEV4ttwVyKqHMixvUWw78isRracfDzN9SRgAVoP30u
51c/QOPkWXlDHnbCMp7TNHQVjBMyQVlfxtJhDKk0WyJ8QXfEr9oQrHqoPCs5w3e41FjxU+dNS4ew
/OvzupGn4fGDmaNGvTcRUnEPqx1V79YvOCwVwFd94e8dibZgoMMreVsSXvhlwqiX4JAJW1mXtJ6o
tAbigVrJEIhVHpiykwh33OJW08rPletR8HVhqSb/ymi5Ka0eG9HFp/Jvx9xdvV5szFFv7cMu3QaT
jE+PqL5zovT7abOOICXmZSymvUhlHq2iLB0MrXUVIMMX1b/PRn/KnUNypMADiypJKwnhSXyGREDU
1eTNJYAzLIAKnqqz1wInvbfNjJnSN+IfygiZCGOuaWLnBFDZo7IU/WRKM7hO6dfL2k1pHhBRnpuQ
aSxRgRyHuLmIz0+Kvba72aBmy7f2uR8xL9K65QOU2wyozneJmYFaceiLgWkXD8m0USHABXQMoYJi
z0+SH0CD2oQG9rLQfkCjMoWf85Kx1dC68cUwKAZ6vgxOXNo9bBbwG3zottx6sOtId3BeIWoyISz7
B4MFyzeMOs2FlCT8DYX+7BE+GdvkKXEXxhJbhxRlmD1CRKqRlWOs6YeoxIfm+2fUoRfCr1HpnSGr
F+zTCiKHT99cjr8ybDmieEu6azEnll4eZhA0exTYddZGCFXNifICP4lg7qRdgs20WPdV15XH2jFi
ZbNquFT2xKn1t2QJw3WCgPSWojV5ycu0EXoARSA/+nfpkeRaCgB8MAAJ8FugQ1B7E9BrIMgIl7DJ
D+2x4sRMKnjZKxPpoDKAHXZtgoGqcyECyNzqjJ0hKoExhnP5JtY3Jq4JziMyaKVJQ8cVyqcPX8jw
UZr6i2pn0zEpJhvFdtCYbYgw5sdiJXyvne063nBvhbF8/5MgVvni2oDzWHnTvlnVd5hYJcD/CSNI
snVFw2DF7Kbvg/idQ/vARXtSp+w2qJH4wdvx58p8GtGSFNe53wHn0PiBB5L1I0LdGCfjIDMUnz2g
+bzWr5VkXGDbfGblmGdKa56lAdPkLCDW0NpPcNzgQ5oLs+inmhHOpR18giVxLAieCrRTi2yQb26D
l9y3y3/l1w4fSb9UgZfy3t4jl5UOKe51vRZc3tdS+k21fudoJ2jc/vx5p2N5KR+HlPZvaWtZk01f
LmX9IrwdaWqMMaLEEfeS8oUAAvsqJM5irRaIw8iIJ2iJZ01QwrNKZ3+eA9KTZ22R/0RfOvp8zA/3
bg4fI3n5Vx62QSCWuATkspZ/x7s8910m52CT7S8NCloFbaHnHF+VYVtHZCAvcCFc243YukuFy4Pg
3udkp50dwrjQ4Jafy/q+RCknV2fHQAHiH6gkbZJj36kv/8NB4ard7WGMBaIru6N22nhL1TIy7xuw
6BSYRFF0TPoXZT8AGjz0L/8Epn5ksWWL/PWBO7o9GI3Dm96MPYXWEVpQDR9IjDHszcu94vznMKGa
5n+m6vUb8DEqCf3JudHrKz7tYb/NnzDLsUVkeXoopfizjpbO8UsCFYJVDKBIWNjQpzhPNepdxKcX
rLAhRYr2CvUHlVI50mbB4wXqRJS+23igOS7oOAmWQZJMJzNHpyjSAt2m1Rb+GHVu1jHTdmzQftbz
wpw4YijAjcMKsEwyc3CuJXJxNLIa7E98VT9mW/AYMDjgEAogCnxewoc5FauaFIp/csAZXJZaiqxr
A7Bd6RDP2qQC8FLb14W35onOjI6nLZQ0Biw2AzNcYFtdp/sZ+vTSg9xYHFGtOE9GQUyLqXvp9iYK
WyESAg4RausC2xloLyoN2oVAb3TQcBdyqBCzLrbKOPOehqcF3ktXt2YG2tpuBtIL2EOdy0P5qtxc
LjyxIiOB9rRwrZKkK561cj392mt7pl2ryWJToCVAljlpHB51I0+OdOqwKbsPVMGMxHbn+kNS58pY
TBQVXJV+wgblnRlBY+cwrK88o523+rkgzLFFMABc2Eyrfu0PePYgO3WqsN8IPTNSyHSPnrcjrbvt
bCqI07TYt24TyEAaVfmmVmgylYIggqWMDBpckWF7NrgD7PJDabATPD0RpV1rqQgXsWA/P862JaaK
XcsBejCdC8yYTmojB0D6CeZqGrktK/LkEE3lsf+DEVzfVoH2hN8ns2abcf1ubz+JWtCtU2PyCxjU
Ust2I7iIfshHE48bvZrUfiORoXb/25BgSDR+hFxBunArO7TOo0NLlrBUDfSgszWRACjDPjZj4b+o
B3rBgrxsIQMF41sf1iDUAx7q9VlCwoN1qrmIXam9MTxpUjxmKu2YB+cKsWxFwpK0SuRktQdfemG2
MxUyiTOR2kWjkSFl5XnSfsiI3NgQvw0tPEBPx4LKWV1GbpZNOQrruvbEEd5Y12Q7LNX13nG1+5DY
Uzw+fsh//CQ+ZeHNK4b8dtQeHThoZn8/MDRISBH/W7UvYK5/oLQtyYMSfwjwQaAM7Flt7D5TQnha
uNv4bDC55QDkfuJjAXcKwZki5DLibjLn3TxsgrVNa7/x+AGYt1SKgToW47zbfSX1hPdfAxNILvDZ
jB+oVX1sV6L8D0FHAZWq7C15GrQpZFgHHbZd7HlqqP3OwurVzFZAp5f1FpmqTWtN+InbzPnwJ5tG
ZVYh5eUIESttUC++6Yf9wbrX2ppKvcjzpaPXwSBMaIGJ4Eh5NwqDmtallhtq7hAz3nT+QPDH0WTk
Gh64KNWFZ1biqjNgnBl8J+ChqxOTtbubtsA18p6Cqn+9mKqLuqXy/oqA3Jz0X+OXSxWmALcv54ZE
1ahDqnGBNZLuS6btzrC0GMAVQNYMOmTAg1qZ5taqES2R8Tv7ObFpdZ1w4YyoqkQVj0uXweae27zX
mVo/zRiTSMRYyXEr8Wg5McEmcT+CFNRDcO7f2/DB63RvnACNb51K9KE0aK4omVRi7uC9bXNXlR+c
WWsF+Lqn+sYXWSJmU5i4RUWPsvkRSSaukeyQcLCVkPnIu7dHFygECCrUR5EeHPMJP0VsTYeMwWl5
tQeH45Yf103TWc+Ymi0Mr6LbBLkmYJHNwpHSbZhReT5sMOfu4L9d+P3K48QrduQPMZAXClgzqdTi
3ov0YyLufbplWZ8DeqYiPzYQuhaP39AJKoKT24M9+MZ3yE0hkvh9fuJgIxfiKDK2L2c2BpgT19Nh
7rZpLxTejYODqmsc3X5H5OEl7Zk5MnUTP8IpCQVZSHQhPiIfdEKqzBHlmRrFKuQSS0Qqfvd/4tjG
t/U9VyBnPPvImWdu/xCJZVmB/CYoqpCPyjJzwnx/mpiG5le25oqL8wBLPByD3hontGdP6SKQYJZz
+N2y/wONiwnU3LCSAFsxE24r4NUn/Ww92MrruAJWRQBGwzNE6210aIrnefSs9MPwxfUcIOOW8btv
EeAS67x8NPkU23ncq4Np5+vsaCLmrJ/x38pSBi/lkjkarrWpFkJQnDvvIPeSDwbOUclUvLNUgMm3
4l8fk4rJGdLYsRiM2kJWainukNUGqHDAsFwDfTKgFuro+VnwowBBrWK8i6djLR2puqd7Z/A4PxAz
n/09cmC0tH1ss0HQWiodWNrOrv7FDynz/moJqPKqDdOV28R6IHN900OBe1fGYxil3xYlVX8rw+2t
V/Bgsm/IhQKNtbFycFS4UUniCB7d+RL1K8ZB7Ks4Sw8GTDlFn3ZTaEOyd+duwm5/69bxGnersnHy
NDC9/sL/UQsw3Bg4Ml5T07VBZWHTJEc5jtymAkSk0oRs3ljxq5Uh3ZqS2247NwSERUrKKYvVktXI
xtj1j72J7Ii74SeY7QlXib+/0QXH2nkl0VZTMsvHxti9cDypsXUySF4g2EJO+sslpZj4ilI4cdKb
50RHC3lPc9XC4rgxH3wYBjNPZpdwvM0fMUQm/r1kPXtrAEI3e4z/5OxDZpwF0QMWaca4Vlbtw9v9
ikjvbdWFaZd0T5PUJ8A2ggvwxgIP0VsUD5yBteM3x4uTbpbAJX8jQcb7ZJVigAUSFMflK1Ki4Z+F
sZzgvoH0bg4FtF2yqjcHs6vugfnknjEp7ZNh3jdyjolBeOj1VYwINWPC1K52gU7IyEuh9v7IXOKG
F5qUW8+XwuTTCf6BDA/v/o4yFLfwfG2xtYGXpxDTlbAMI+8iHNKTfYlt0XdqQds58Iv+qV1vDfr2
MapyiRKsNtkgcHQOEOoc6Kt0rvq/yteWy0XhMKliAP5fGTE3cFtQmHS6iWWi8vzRrw/lfe+lXhPO
E6bbsvKLpVTaLTjjd/D6sBjJWpEdLxAW9zv+u7YF0QfRKsRNIH4go+bly+fqCJ15YV6ZO3syUZ6z
WaNwDVFhnNj52LOS/SGUO/WaNHKIRrrQwd4s6uixrXPkwKQzd5CJuht0/QSjvZK6F/TeDS5jVhlE
5kKhURANOUeO1O/48jJmKlIYESDkKIT+fwdE+5Jt2CImNUaJjkgz2lc+GKz2YP8oXalKNE7Guoj5
z8m4fq/LzIJKKUKLPLruyBlk70SE9SbSMKCJZ5JX5xur5Fz3V15zQKC+SajRTQTskbBiuTU3qNF1
JBOW1CiWidOI5qts/VQ8y+dpfJ+b0EKqpx7G3RyEKzreZg9q5qB2b+zHRkq11q2pv2wf0qgJALPA
InK8PiYIlyALdoaSgCabPtw2FnNsJqGc/SkWjUzXY0puJDBOr0kfW7GvtcbeKWJEPT/l4X1Hh5iA
ZN3rPTeoUcmbp30YJHbd33v71Dnd9vCE5GYOTqcTbKy3/LyXD8Ea+rsklsLSEZbGZiT9EZzeDsRv
8gY15Scm0nV432wl5shKv4nSshO8LRBqZf3FTcoJxn9VkoNDSgZhvnp0mwTAede9t+ohu6fRCoWZ
FQajsxc9qvtBagkF66ndwuqCwlnuoXMuDryww/OshB5AIN7UA/YEfiEhr7QwkvXTIHsE/ZS5G05y
Gm4EpNM9phIcEQ1yD9f+H+T6DZtO1szFHuUFUbTFdXUck+zk2LzBPrkAv8moaG7Lft+afu748Lku
C/G3d1NZamGlQHI2wrkc0fjfNlwaR6IPCOh1SJpTtg5fHrSuz1wdb5oa4rMsH9w5jdkxX2z+N5xP
1fO3bNefyA0l8ser534xKq87svYjXjAmh2Rpqif2//kZaACCe/Q7YmYygRj46+zrbzYXMfpDoUm3
8xarfJIgoFcxfLJ7UQwpJ2XtVDiis+T23jNHSV99xucY1EfLp0E5e4kQCanY6VJQV+xLz44ePqaP
UeQZ8iL9jUqcnI2s+CRYG+5S6eNt003L/sxJNEhm03yuD8wGndWdLnl1phnceYZpZ+dLDkKhDUwO
Sd3XDIiQe203rUex0bx2jg//ONHB+fYyWNDCEvpyREJdThA3KqfHh4X7hjPUiVu8UisqTGAkmwKO
+F4+ft8Tjlcb0cTWEzX9KGhHCJMYLfIKzo72lFE3r7ud8POYbYLjGkn/kSMvX+Zj6flUGuOZvvIM
seXR79Rq3FfX38aZ69PiXE55GD6DnekMJbCJ5jQccdru1naxzy1wZySLoCl9lTf4LoXnBM0XjnXV
GRpkSADnZHNqXhsTW+nEiqhQsm9KJ/bh42eBKW5Kn8XO6MKDETFg52E+WcwhmhT4vzREj65xL54r
nv+jOxw8dsAxdVXbUcxki2W2c6QiJff+vrNSHTbhDxK70noYhW9WuQPO0BGZoUG0YNTVAU1xbFAw
Rf6tynI9YFhwKCLNWc537qUVXB5/xkRAGuRDEb7H8g+0DRNmF2OFS6DJIX9Q0zZ4MKHeQu0iYNf0
+2EDn6VKZvBfKEsDcAgfdpwp46lDXwefE5l6EXlA/KejdenY3uDbr/BofeSpWHbg0w23KR9rvDPf
X/TQKlnrK8ap94LK1CnpZDxXC96sVOKY1+yuVIKYSCuQi76VaJiwiE5AcBR55aHvIiuHl1FKwUOU
Yw6XrZ1Wcwxtxn8NIecxAexeAZDT0xXoU4Gk7EZLlw23XL00AKZK/P0CmisA5cIBwuqxf3Gz6AV8
6JjklZwg++u/2G8exAfBgFk04xv/fmhwH6D19vPTD0MOpOsfWSpry/MG056q3r1kNmmrbSAk0GsU
xzt3bduydETmjy6tNgdKGxO4F6+qJUnE92DBQHnGUm1an+gxzcxOuRmVTvFSVcgudHO7Wglsf1aN
wUadtcELQ12YwRk3197eEWwj8TRmcoVM164+jx8VMCbtMt/IzsEZ+3XN4WnXfj7oGvAyc3ckatfQ
YUIw8G4AU66FaFizq3/nzrT2rDyBjzIsTFvwlpXt7qrJb88Zv41THaxxtM3Redf/4pxhfJr0lfWz
UbrE/qLu2DdH0qS02KgnFf9TKFyk9xXLxp2YE+buKur6Q930SDQcrLqui+aTyuxf/qyUkU0WNHnI
7fJKrSiOA9keqwnG3ke6ne793pSF3bJK7u9qOBuVBafaZQFIieasyGz9fcX5y9IN0SKHP9GnfOx/
Z1/0vZ5RpRKWypndzB8yuAC/Nbde2MO6jpuP9SdG/A1bd7PjyLFertRxezeGFAWAU7mn0pL7vrQ2
gWzKKf9dhxDJPeJDq0tiG5dnaL3PopA/9zcxlmz+Kqyd4jfgyDqvuVXPnN3qyObNGxzIjpyvYpco
amC61/DbGtAjza/4Whz8K8UOdHSsPiS9i0D5CAWeI+n+/zxLNuwkBd13qR21tFa2Z+tiBJJ6TODs
/72yah4vuYXLxKIa8PFqOX87RcTPaAfic224eHLF/3ntKjHTeh+b5QmBCz2MfKbTpRRUdSqXONsj
4eVzud9QgFftuXpQPd74AXdz7va87D5pV0e/r4vzO6BM0aHwgc3iSMzjYWcSnnaDfDzHqBny5GSd
WUztnKol5D6fyK2khtf5PWhhgOURQQIa2yZNAVTFeTzjaSdxSfnTf0rgBJw6nNr+b1KXLxZ3ZL3U
GkZfMA3KHW7FvV1g56FKMHNTHts6yTZWOB69i+Eu0co5NEQc1TayWi4fq+MVLk0oCAuZ49/hJx1G
bpBRFrGfKTq4usxI5sSzhblhu59PUWlJhKrHFMJS7w6SamzTS1jrV/pgAAWqFgLh4RmkB2+z4sTG
l8VJueVrLs6vEMjiON5/TVylk8E9kLDCcHxkOwluP1CVF7OmmSS0e0fY1DjXeeqJ4yPY7FdE1A7p
UoK0pbuakrPZmZrXyTnYI1jlrT9aO4tm9LmVot7U60N7sqXmLyFkAwcTkWqYYzMQCJVyHzh+swKg
cEkZiMwiUfUddutAamBRvA287X8rVjQOBODV2xt244doouUyT4KhorX+j+2LeBlhKrPRu68ViYzT
eEL+OLjmv4H5SSY+0kruEpWvmJTKt4R7/HYj1P04CzHOhAJ10qHKC2Zi1jyHBxxccjm4naH4OpFv
fzKth3fj8KlHZv7pSb8ONcQx2t9g4w7Qk/9bvZWwq4JBV3cBRI2JI/A+qiyaHmEgrC2Qckidod0M
5gl4YfAmwgl00CVI6aXwoguotYxE4s1EdjiyU+uuxtRsNOjj4nsWuQC++ItP/lSCmc6Om/i3M596
THlIBT5Q2Oz9cImw2YsxIxTLFPMTMRuTdMuWBJBzXmRgSa+uQZlbBvIxGroyOEaR1zbNCUDFIvw4
AmHHqUqMDqRfP/NQ8nx8wqMbkwDN3yvG64ZZS7OfQOtAGORgJvOwNm2ZUXJC4zrVCLwblA/5bQFX
a8+PsAHqod1ySLtOo6GiG+Gx7bPfWI11i31YdFNeGS2sXHeWu6eVsIWntElTLR529OOGTgES3SmC
Pbe9jYEEm1Z5BPUHUMJ78VgMHhOEtZSjW74URl4Lel3hx+QZlgLt80oaJmpPZsJnzCgTh+aZEtTI
+Z8cGBGw3OHxzXEgC80SZ/Qw7AStpJ/G1t9k4y98WKwCClBJwMo4w1BM1lf54lkrnxAj0KTvXqtz
4ErwqGYDWqVzWXJAs/833xNEZ9I5S7MGPRdFSjStpVNrR0Bt8Z9Cp/s+bMy7mt1zIiY2qNAEYuWI
qMExJFY7rN37f9s/jg2VPnHjXqtCGR23zXok2EZDyPy4VptDsT204YfRI21Ai2xaNPThu2X4pftk
HtkVm9EW/OrzzMGrc6bv4lRuiblZtYDrcBmRn6aLUYEo+Hq5VFptiDwidaGcl7hUsojxUO+vhWb2
5nvZ/4oXsvmUWiA5bhlBJvA65Z3G6DiuOY+tceqCImW3hG4hXAE5CihMrbDXsKZ7L5QBmoU6l7Zm
4szlKI31ewdWZz/rlM0WXQ+hyNBD767rJeMQ5nOOsB1k6z5oZV3cZPmkW4ipEn1moZHrUVwnL6DE
AQPFtoIbWkfp1gY1Xt9ZF6XPTlo6vOrhhfa5kc6eZJUL7rsA2IIzfD9pE+j0Bwlqvbq8dAOeJ0rh
6X5hjNwD6umG+NVNasjDv7Yo/ZXkjgMBYuNkZnKVE9oKaY9WmA+iVA2A4qLiAYUenw18eTsaferc
LyL3IFB2c1Nu3T+Y08SaNefTVzOy9o3U7D+/Ulo/JbIlsOs5In2McCYRjxz9N/HGhFL7mBu9Qat/
T7OSiCBRuBq8kVpF7lsG70KDxcamqtOzH7quSz95xOiEWEw7J5l0QU5IVzNP1QzYusGhaY+otIIG
HFp/+ZzvSA4zhZ5OoPeLvz81AoiGaGUCEA69zSYUmGHNKAqiTnHVzWZD533MiBhulfNz7pPUuEk+
hPESyMsTwhDjjOVp3elPXST7G5C/mKMxKVj7dBAHJq86d6WAcXqBycqTXaMm4kvhOOgg+fwPu7iY
KoE/pZq7ONz/5rwx0WU8cSydXC6lRIq84PfiA4vRsnegWvoVfjC5HuX2pLoXiU7sp9vWeAgqdZ6p
85hgMqEXg62FEOXBPUKPBuo2vVnntKuHWxLBFlp9mwLtvHRRfGfjZzDw/DABhCxnvtfPPGOtwfUf
PiYkupzbKlIfTMu8JflwaBPPEPaM+XIRz+oNdRv8L2jvtkDNRRI/aVrhcCwFyS13Wvyj9HmLEY7M
4G/mOZzQAhUG4CBmdZO0k8Abz+oB+vQeAM7e2ECe+AlBsNfW2NkiK3Mlv+uzMqgcpL2owB8zbNdT
qt6CMLRY7iWfrshXrEJYGTWOaK+EfazAKSXkTFB4+TC+BWHqmAqtunvAIyPrH4RUyqHwWrMTz6Pd
wnneR6j2gSUdNlilExoV8ivHsSbuaj/ZAfXiVYGdP6fLCFBYuKZef06yDjwo/rOopVfiMfGAWAxr
WwNgLlt464Fsm5giCSEd+Nz/moFado76VYfyNv53KXTkZBnZQziKN6l4dpLCk2lhi8rdjL3W9GyV
2Iq4WvabLa2IpcOZiVJK2AzHJ4M5Ub3SCtHtZcn2L1fFk6B62OiUqVRbOxTkvIJufreXdHxgg2M7
058aoyCWOhHykWqcXzWsW5QTqSU2og231eJFnZQFW8ELMgoI5jSKRY83/ZVC+CCgqywdA3JoV8NJ
3DUc52PG1lloUot+zPEzSW9e5XCcVh+X2flYp7uRMeBQ1RYOtdaG8vq4IXpHDfdioVjrrjNnV5wQ
qXx2mC0iE6ZzF6iL2jrx5SBQzuhXmVFZQQ3zndHA/UPeMv8LhONQlTA/Isnf5PWibiu5e1Cqqs4H
OJ+HASpZodzf8C0qo0WwB243mxu4aXk7u//u6RXy0nBR0U41ebrsE1wjJyIbAVkYjkS+ROp1DdMj
HX4O0nygtFz3pc+mLqWQZWRThfCjgHS+zHQJImk/wh3dTYQTGANh0Kidun4GpGL43pQPpxA0IKbG
wzKTEu2ACi/M31UmngcjkiT9OEZGczCvU5YWvYymYdAT5qUGUqNhakWpdvtYHOMBrFzEFqBf3atS
XaOGxiF+qrLN80GHOv8IXBJ3wMflLasZuBHj71wWICKotX/9EA+4nCznGqz+XoYyWDJcEel6r/tC
Njjm7S9nQim2GSebeo8thgYUwFNq9RZBaKeqdJ24ab2+sWR3wWU6uyxv2d8vlRZROUAJPai8sESL
djpmijm0aZSzfNHEECKvsbfkBNbXGuNrUzWkWUv/Zer4yZJK/gmKwVcjgEpJx7+X2G5ArlNMDI2Z
UQQwwjrXBOJO7kNeuX4GJw3BshkJ0Kx9ZNYhaUtzNkdampbmZoBuXsEIhMiX9bdN9b1ejrfkftcY
0ljJ2gGK7kwKc2c6dcdge2Fs3INbVhedsoVZCgoBXKSwUBFp3JUE7mABYAyXM3lQCEjJwmTUgI6V
zm2HG7qQoRl/8yI9NAkeo4hk0fDUd3wf5MS+xKHJS23S1L9v8XamInMsLE4BcZo4srGC47PS4+I9
smb3ULzI9FhTgnvJeA+nKdLpFuw9tBP/vmJHEL+l50xJUv2AOz2xiFKJ4gErR1KeIFaUQInpoa5R
PQyRhf880rMd3vAUOLCFNTHdwXLxv8dGFWBFDIth5utAOeAfCVr+1a08km4Iz+i5+8Id+6vQO8OY
6mq9YuFnzEzKeRtXMITNS1plK7I7uj/RE4Re/lxZUXelChJNAE8OX+kYlvXE9rgxz0SC7DdhlY/3
xqOoYDx8UK8kNg1zl5t51T0L1h3rdFb6YmY0c1Yod7XSLeO1lhxV7IcCFuMZMZ72uG4YQrYBAW4G
ToBqjDZkRjvsQZUy69Tw8y1GwEUi2CVA06+djBrjkRxUIDeS0j1d+lg177Z2UG/reTo1nVVbwajq
OweWxtZu2tdxmxUgjSHpNAh4Lys0VuCzeofoEd70ZxWJdS80Gr2MIMme0jA9icOloeAKjo+m5Bi6
SrGpxaSucUjBhKMRlCdIGSBckNZ+/RzHZAv+7XSALQceLqqH26IXFL+K5CU97rZNCAKrtgyLvAD0
QoE7iZnUutMdL+de4VDdWmK4GLmQ4hgfJgTh+yjH/ulxTsxyfqLTrtFGFbZnuhRLXnxJf2RaVSDP
UJDaz66mSD8Dv3zh2Q5jbD+gPME0WEeIRBixff7PZqMD1kCdHFAXoVFRCcoaCCr5KaMjpKgjOQtP
VHS7z8iFZdsOMiKpX0/DisEkjPm1DIT9KOOG5QDzB8a0IZabpJoOW6TFVfKCAl7g/3LtCXqdS7KP
ez5tnUXbnSddD65bF5Lp8Pj5w+UvXmrTTpfzAo3PPD22O0OQ2J6bwtB8Sllx/3j+sm2B6TvgPrS2
zfCNTvOHJwQ0mugh/dpLit3L3wTyPT5z3F2I80vUbk7K6LvvSdrs1zAN5j2oX45D/ZQNvXSyqQyd
rDjYc8+Rx1hdmloYvIKrqSPYL7wJJiD0b1y5iEwmLi2Bb+FePFDJNsH3jst2qz7UOyXoQIY10Q7X
F2nAaxsokXMShwFwTMhjksagkYN00ZsJ2K2qEKJK1IMK12ZFuhaGqc2oN270U8KRodtfz7XrSqeU
BgU/6TWyMFkfHpjWVzWU3c1B3h2X/klFf0fP4uCBL5V2k0QHvNrUsi01R1tcaz7L9G93WeTFSCRF
lZ13x9JMjQ9xVPHOM8JUXGJSNgHF2OhmonQIpfw1jkHMn+aCL/LGgDkWCDztpB/ibayCgr6xA8xc
oYXq/NtBuTnsx6+x15t8vWetM+tQYVg16oUU+3AUqiUfsvHu2yL01oT0nsnFbeLAo+yn7MuENuY7
IiWCLpxe85XSoi7XIygCajurbpphUOUOpn0BmTB7tqa69P/QWu3XxtGqvssi/5VUSI0wlRnRlr7d
aViPfW57KUFKIwucHjfX3pK7wDg+bfYGoWmBnffEnqXnPZuLvX5c1jTWD/GsA16aKpTBvWiJai8e
i5ARy6kfaR/fNK6iahvIUKGVGZB+EXR/XVhfvO8T0zOgKt2nLslZBYca/u795RIXaO9jAWHPXPpt
HQ+L86CnO51VvmBr8E8cyzDGvHhNLHjvP9ZXtkIY9n8YKArS70kIcFmpqSuaI43/LYWUggZNXBzE
zIxwfghkYrbCkHLQqg63WytdL0Ngkucz+nA6SYhMmA/vRG8OO1kfkQ3U3+o0m1lOY0vm+s1yAR2v
7mU7ilB+xqM/75dgvm4EZXUf2Oj7jFZ+vnzLZK9FbpbXBStTMKdrr4GYRv6gf/mcyAZVfQUb4q4r
NxjPvhLZzJ+P9QLYgjXccJxg7h2IUM9nUT6BhRKUS2MUcBb//Vc4fKan054P3QoDOJRy/M88T9ux
9gPsbtlPL/r6wvgmXr2kuq8aKNZOlVuyKEABi8Y0ock7wAuTCZcoL860ohBCUTJU/DvMMFqxW0rd
MifOVvyCsdU3Iy4W33ds1DbPvM8B3Wh3Eoi0XBP42AvdxV/96n2Da0m135Spk9xc9u/AFmfaNOAx
lvyuLFUccWJeBeX68+FM0w1Xo9HzA6pENxe8qOsvEuOehg3Y31vjvx6R0OSTyCifbo7UWbNl1sK4
25arWmwQx5PaYdfZhucwv59n5ITWaHZ7NXSaivDtlhctMpyBw+MgYHZgUx2lqnjR1M/YULYHvIu/
V2rnpX76W5tpt5jg+jUJo9Q53TEDXOoF42ECp30rMdz85RC/srwBsF2Xp0vHZlOg7EzzGgrAoyvI
sYfpLx1fqIBl6n3PN6vFuE84wPkwnDtkELJ9kGvyUZ/oUrgxfqA4KTWnNsJIkyIhnTQzVzMZyiY4
abBVay1cGPKfOfn+C8tUAy4x+PnMYNqK2IBcOn/q131Ui4+yH8J/WGvHTuN7KBOtEYvv/z4T9cnY
av2qIhLi60Cww2pdEYtpPXpaerDs2nTWyriNjTi8apnQvn4DNrgHoeu7XlhYLgaNBXnFuBA8ZEvR
7CLn7Q3aCtVKogmS31imcvX6Fe+gB1l8faDh4CnZ8mw80TgE74ZYq/TycYkot64iXtzIv/4jQ8gG
pD01lfB75BFjCHCJZqlAzoLaCyph+Tc/yhBOdyHRUHHluUFbtSgw/bN3YnEeVvWWIVUTlomYCYyk
0ZEU3lKRKtPUzGolL3plsaZF0pZQjC5o17lPZ1UU17f8IfsvXRHEa1oGKVwBJnAwAc4vy8PvpOiF
qcItkusThNVwjOPhiEGmI/lAa+LPEggpstoC8KA9adl5lHqbZkiknHtRu3UV1SjFgst97aF35p2H
uqpdeAsRhhGXgbPwyiEFH7tVRODthdDDcLeuzgJV/qWFMlaC3TxDQ4G5MxqJo/AM7hM1D8hI9MvB
KT4NcBOKpT/GMH3Blw2TosALy6x0r3TpxfMypuVtzzG/FtOWMbzkavvV2h7XWUOdY5We+25bj8QM
hnscwS4OBcVOzZ7+VkIWUYfcaLIbiHCSWpeuxpBVzlSY4E5mYNVqz9zlfFBuBUsUxqywTdu0YiXc
H2+59XtpSiI4DjoFGxeQ/BpbvgXDP4FRuOm/vsk+VXGr5q+WFIUG8ZnfrvNdjbchcuoGxZr9grSh
GCOuWCK+ZCLzjvlq3Lvpe7qQ61t5ZiNDJ+7NLjeUqZyMuyKADzFvsxQf2x1CVhjmDyWl6eqMCgHb
Zf6kIW9lWngbEGwPm20fFLQeaxydZz9s76m2kqsTs7Y/Tvg5QtWp1yOiDi1njQMpylAsHwQr6V4z
pEN/wMIq0h+NGyRTQZXdcO30oDichWf//vCWL2OihToZyLs+ElBZF/uKb7SrnCfGLcm4lL5C3kCp
ARxO2AHU+3Qgfh/SShq0p8pcp+suLnwhNzTiQmdcSAsX8azIWCYpLZZ/+aZM+tSP7rLp0qlRmKOt
LPbWP3FbW3vXenTu9DhhjIre0yKwJJtXJKMf3wfawHtWaG0bxlTqNYeNXKzCli2/eOYR+SednSFE
tCdi+T3cMexTe8ffiNgPE43aFxcTDrbQfe/Ao8ftVX5XKvmXI+LGX/DSikYkRfYlD95dxol0duoP
biHiPIvZV1l5DPRA6eYHD8InRLOnnWPjuM/8tU3J9aTZUgnVYEWz68BAy/tuNJopCXmLJgEZNO/I
lDAu6WJ1j3luePrYSYBFkdgewwyzfeDVmbYz7jVs3t1HcjC45Gf3lJ0nekA9ytZFyBO7Ayvjk4Co
ggQWJ+TZ8AuicherMHASLQf5UCjJKE899ra174VhPikA3hPD1pbwan44hueThmsyFIk4I0nyOPUZ
F4JA85E+wmN/u96yOIJXKJO6h5Jd8UT8k5b9nM6lYpw23U46UNSYmVtPPlcht61Ga/Pb5s9Qz4iK
B+WrIRC+wHww4ooC4iY2ipIqLs+kI1cZ3YoZGJS0tZNtVOM0IhB8Mp0b3Wb/tHlPFQ3R8e3Mc861
3+kywvlTDwK/ehXWhIRIobfxDOAEPtG/nwKQkBYoyqJgkYayiokNrJkxtdUmOra+i80JorV07r9H
eZc4g+/2UTyEjsMBZDZVR9E6dv3I8VH/Yz6mHUbPhfpuyAKm94Py/dmKhqhPQ+f+daLLLErUYaxv
1k3TZIgYfdZ0eEL90XkXWy25HvaEGLYXNsqNRmJuYVnMqhQkpDbj5TrHQNjqd1f7YzGz6aJsiykM
z7vpau6zCtVNrgUqOjqBHaXIjRn6PobJ8KS6G51d1O9sgdfF9KaWUQhiS5K3B5aWaAgp3jVqA8tN
0qRzWPgFcQZ+BNqcgxLDaZxfPHI4fAF95ui1tRGFDoWafQ2upkbsXQmTD78dopJexfnPKPvbe6y7
josbrAEZUTmOPgcHfcRksNEiDz19ZzHj0ERnrNUuowJgOaR1+a0Gy66RfGjXC+9h+35V/quHhovE
caJXCsD5O++Y1yCEnIHJo84d0VsV8R367sMRIq5gi8gbh4PDqnPTSKo99PiwnntExyTccDyiet45
zf+zbI6RdSZ+h50TZQdTFR/HEp/7V5qLQfI57HL1SCR++cT5+nLGcnVz+XrSRNc5KkkhJKoybIxO
69mCVcHYUuEMsV4oI9EkFIyMIlCr09c2cHlDyXipMdKxjx5JRcA5dSWIwuBi1HB7ni9oGvyKDPQE
sGXHV/5juZkBEOu007t26vh/GzHy+QZZGB6eSQcdNbZXz+00v9ZEZFRwwwNOvyvHmRjgoxb2LRPy
vaIky3FlWoECarZiRwkT+cqnO3IAmDUKbIbbDQlhodNeRBNgpgmKjZMDWroCuFao0as+Nz/WhJo/
+UGSf+IjZ6ZH4MHFl9I6vd5NjUOqStihY8vyKMmRrrViwiCq99irgcYZEL6JsonbqPgDepNRhTat
n14MqAQxx3JF6Zdazopq8ACtsslHlz+PFzEitjrOtGuo+INBIgFTw4pPrShb+r7h/C2zRGAaP72a
gwdghCU8icZLFujc3rHeKJ+Zf/Ep1xMTMUlGavAQ0ysgwpiDyZXJ2/cQtju3pLjJBK/x7HQEp4J5
l8O6dpGWKqTiAI/b+AFqV/9ocTwSKc/EWjNLv/Dd6WzLLDIG9ncPa2jWLadXpkkVWRZVQQkyRHxz
n1qAMs8qxzVWxBlWLdjVfxMgIruYEtltALxAZp/ioVwiruf3EajGKNGOqGndsXXEw5TeTP2yhFxF
gDsgdQCCWE4POGv6r4E9TcvNxvTUkR+Lsigoc0Jhi34m0csdqqK1+LbrVLN4tAw5dKc3+zIGLlZx
UdBQ8KzMG5rOvVSob6BtQUX7DlIY7mnTVG6NlFyOGXx37JWOWxEFr0uATZ0bb3W9Xu+5q+VMA81i
lLpac0ErrjPea+DvdX+ladoQeLUDVL+uoMMA6D45jFOM1TSXm5acsEsGqtHH/cM9aG3b1TPW7X/y
2WlaSf3JqiZ0aNI81PZjuaZwzKjvDu02tDqgzOizc00dpmf1Kq8sbgwe8XyRKOgqfp4AwKygi5QG
iiU5CKoTXzAgtCizsmywhg4RY7fbYtjwJ94wZLKsiJE4kHXFiJfd/+83W/K7r7CPgNvd4UhHXKPA
CRN/j1kVUCI6auCLAt7w2TYXVkh3VVoIuWv70eoI7G8ONdBZhewhljbBNkPniLTfNgOegHRtabe8
V8QnrSAaRViBa1EgErKYrYPD075+XRC2n7+x/OTpMbMYZpMNfjwOKpofVz+uIU6TaoG87bhhveZG
YaBo4DgeZ/QQSQQlpDjJM1xJSc6teWqvVHpnzoX/OaVEvpUfpH5Y2Jvi8+p4Fv65RzFrDxJ7h85L
NwmaFr7FU+35CGSqqTR3B7SJ42VRaMq10vf/x/K/t9vaFDvojHGogw+uEU6QFunUOqGGgjYx4gMz
3xRh54yYUqk7MbhJF2verA3eMJnCxf9k56bOwmJH/hupb5VKMmDw5AODGfUeTVb7FM2opUZ1TFnm
VL5ae9+Csg/3aKV0LapvLyBpDPxQ9tKvcbxsYJIHew/cNV3Vlbawg+ZnqmG5xnw4hQiLSaVmQzp+
ErryUhGXwiHIIADGeRnnEdyu6NE4sd9q9wUMDaHTvz51vJH1wxLM0XBFo+gK5GenHK+KTQf47IbW
BTTdo+ImbPGoTmxm/+JRbgkH9df6ddr845HgpHaWIertBv9OcMos4HUxtwz9PrrBIn5GB/SHPGKj
ozk9w3oYkGGVo7kMHkKxaqqh2pltvsm9dNo60sX0m+Mrbd43BQx2fuh4/ocdY6yXBsyeEQlwOxHc
/y5MjPz1y0Y4/3ZTmcQOJ/HK81ZlBjCUTvLfoq2olq7GxOaxHCtZfxl+LWcIVLmVZ8lkKS533sqM
ebi5ogRaGopZBr5ZsTzViHmROCtPRG6ruoMSwuCrpW0UHANMKhcnt+83kjU2ukLi+pxhzJq3OQMh
TO7D7vNUkXvs9ySN8NMwpJvzWW+CzePPm9d1VohTjjBm78c30MZJwwvREXZ6QgSC4leULlqy7len
rpVjw5VIJMBd+bPhrrrPAj4inLEoJQWNbQQkMHrPSaIKtIBZeQfEelf1bY94u8+rXrzOApReTpHJ
n+Jsi0sMei3KWmGrJChMD3vUZ69ytHGbAKveZfReELInuUeGbaVYAUFCBgkCT3s8X0XKtkjyUsdL
zKQOH4VKqwlmgCXgpS8DpKHgzC8YCrncop/QIsuOSniNvRX2OXfJVofqYBP/p85g8IWBZ+nBFI62
RDlwhZkFhJRcqHNhs48t4T5iVikFtWbAN2MDbPFaFlSbHghEg1YYDifx56nNnnaBeFhWKsY1zX1w
ROnzTjzKxTXFaiuIJvcFDWi+1LHlXAtaepsxB34vXpmf5r4126ApXxLSwnfzXk4z/epGCtVz9/K4
uJsxVkmE0dAowMHu4q/pFbZcWxpj0wDgkh5HuwRWN+TVfnc6Xl0p4B0pwkRiVl81bdeBfUrVRl0t
+X+pqIEq6QV0OBJU8KsN9NS5er9O0sw1h0S8IN8rjfM7gmN0812dlbIDvssX6PnSlA2NOorgcApW
jgJXzquLwwJdneQdtE3qnwwVEt6V/o+hGBSDCB3I6AKZeCTW76sfFJpjXjoztYhDszWPYFfJIKxg
nkQ7maaW04ykDFsZmYNamJK0m79PlWdTFq1tH8MaXc4g7bcmaIWO9u22e3dJHspUxwdRA6c5oMJA
p9/RVxEvd+Cyd0OxIcdu53ztD5BAbx8bNZPEoXiDqrSlGX1wJzjw7D0uo6RKfCNcsmUsZEeHV6ZA
s9bfTtEnrEsx/sTIXlRaFa0L38xGZOjo5kph7hm8P+GvHzLtRaSkls7Tw/PcSum18ATE+yibar3E
9BEOaZNU3mw1/rO15rYJ3VwOaY4KPfbOro1CkhX4AM0KUkRjW5f5Jp+uEJNpDHDcVMBOFDDk8jza
aZlQNJrUTv25sdPXLB4uKSeJZrekGg8j72SzFDD5t457gaTtZb4aldjjVTML/L4HRpELIwQ8KPV8
cVT3SFbleNV5XdaBTeDSByHAN5BKKs7PWOzl8TiN3BeA4q9ag6Bk7YVcubmqaWVMyH6W2kDP5DIT
ppCpXBainNTrdynMb4ajKkVzozaaJKCDBoCmpA9jaHBpwYckA+erQFuSrfc2ZDyetLzkHuhQFAwN
jM2ChI/8klOR7uSII1RwH2xAfYOQt/2yuo48or7crT0zDO49SxoW7YZXXQ39lUAZ6Ea0ytX3qqD0
O4hmDCNPWrOTyWe9+j6RGJ1/EnuN2kV076U++nWsohA1kFw7dYiCGS7Mvq+wHekM80M092CgsXDI
EvlV/6HKdTTUYbba9/2dn0PjWZFv6zPGF2PptzrfHYKMZ70N5nA2QdRmAKh0EucoRBgqv1tZUQUr
V3VlSr014pywGUE98rqVYo0pqMg4sqwM6QBCetBitO+lZsstews3hyUMp1ahNxhHvpgTw46WWOCB
EvIdauu0Nlo3UIHiR7cdLYO2qPDLihRtq3VMlooPAxb8XoejiRrfo+O3e0mnMPRJlqSuPsJnDg7j
B6SyvJANVdUUiD9mJrSivhe2VN0BRJQPAwV8EnVd+2h2JkidmkTms/wDlaroX2jLwOBXp24pYj9y
ejIFlssoNEQJZFT4MpNmWni0RkNv6bDEYlz2xtNqlkvkt30igxTWQZaMImHb+2p0zUvRehGOgWZT
hVWn9hZS5PM8crrxtAquRbVRNOfv3y5QcWoXecC6H/SaseeIu7lfGs+VndCaAv0WRK4nBYhCcg/b
io68sONEl7cs3iq5S2dZFlaqoodOYi6PozrCJSg/8vjcP88DlsZ74JubcMyGYCaWkk5LNe8qWNOH
VlbM8c9dzwlEK2sQNpFM22S9BKmw44j6t/vi+h6gsWBuhTShTs8DPBt5L6JEzxkiWcqBE/rEDIkV
Ct7ihj+lkX2zZaD5YUmJpDBZpw37jQvBQaXVP9RhoSrO3YFAHOD28O+UWWjKwD0keyASHpNDBRkw
JtQD7/sY2Z/bdp8RudZtNqaND507CgGiq2ucdUciHaz/cB2Lu56BPJXCuzeLTn/fU8Mz9/tV0u9h
4qEy6Ye7C/xwdoiq9f4D5PJ73wX0RP+VfJQXlUgfcfpig6dpGpJZBVVGFhXDVSkZG7diHWGGdB61
CSCZRpr4FXo3zXSA+Ri7pe0/0rJL+3FnbskqaihsybFAGn2YXsxX5m4lpQZ0wz0YeVW6iOgkgXeS
YK5QKvREEHG/TvVLOScmHbQWDS+0ZOwzZyQKsDtqJGZ/i3itaZ6L1a2BYd9GqEXeB3yoNyRITdQw
ZIuENFif7TnZwEazcdfYVRQwylGi73Dr+e/5jDOzA2sFubJJdy26uabVhb8ZxYfo4s2IQcXGjuZE
t54NLMbhqTukZYQD5nFEsrfaJ1xZL7LD/JQIXJ4Uhl7Q1aciNJSdC8XOac7piS4l3nhQhReaNhuq
9tOD7agfT3b2toDW9nqUQjdSdcdUc8qGyetg65ifKAnomD0i0YAF4fY9I+LH7tiJbDBimZtQlnyL
nzq8IopX2JjAWlUpgM+DnIByUz9jgr5jW6SrYeaKmo1IzGH/m+OE7NGq4IqidKuSrh6xvbj+Au4C
YUjW/fM85dgtmsusTXOXC/gihCUr7Jl0VvMtPtEfiLBIBZ27nuZR6qFkN7zAClFABb1HR16c4KLt
OQsJfFOXoHlp2pnQqLd20aSdLSgYQl2j1SWyGqnvSCHCmA6xOr04ViQK4P14n39+zZzQhbUHMIPy
ul7DvisGlvHkmXgliYQD3+isMVJCi0WWdufXH6R4IoqdVUdKHlmlkt+C6E8PauCIVWPM+/loYgKL
rGjGC9mYHwrr9+TSdWPEPsN5J1Tarh9DUWEz6Rh+QFZ2hVld/jIrGp///3K5vG0pwH7hldjOOq4E
P/MZgesqi9Ndf4okz41xfw4yfHs7Byrca8M2jb/TjWrMZFRr/pRMz3lgjx+Zjz+2SVNaXhgtofMt
9CvrSGVviqbIsEFZ1gpvrWOBGi40E36cuBkrClpglqBV3VjizXgBIg7Hg0V/H6KA7L74g5Pe7T8f
30t1dH6WXKjU3FQO6XcAyAYzsX8xnCA2INmUxPIaDTl7kczeCuWY08+jfeGfJeCIbiQ3p5wTGcjS
lzeQSJvvBh9KPWR3u4bKkRFTcYzrbSOK4kC83Lk2V3LivwhKaZlVaL8kDogldSpIMePh6nxAKYZV
X4FwGsiWyFVlza86d/xpHdsZSREV2hd5ilW9CcYi4mJQ7AgvOpsPTyp0mdJTqq3AyN4A9i9jR2JX
0hwsuto+RJZBv0F5pHwstwqLrQrlaeQycd9TJdEh0jLo2klqjToGqzNCkA+B2oSCUEnUWulcmgbb
UF+QoyrB31oiImpVdXgw4oUqrWaeiv/Mzvmyz6KKapdbi5FK2raXmGHp54mPmPt646sLIocARFtz
qpLeNhfm3Pq3RF2Qg6Jgfw445Wtg3yrlK1bKb9/SqUN/Rgj7tmKq0jWEaPTcYvu+JTEdNjJngN1d
OdgFe/Kd9a1eDPaEV90uO572JG/UMw96wWllNIWvQdnVRDkVt/Nb51xQle7wtIFxK78rMzYccRtU
2iDfOIb3P9RgemL89eb4UCEdcScrFg4QYJ+KbPFA3RgUtAL+U7gtn/1Kdp3tP32SHl/VlnUD0PeG
4yvaEclKGzuEjZ2Gj4uPc6XUELWbiNA12HRnEav3dAMQMKalutKQtblezWOZmRm44tX3U0lU3yNf
5VG0y97OuqyE2z0VS4Dr/sw3MoMsW64tjWUuInGiQI6MF5RmmBd4ELKQHIiwrED2N3qjutmwK8yF
sixdXflScPU6x0IGNVaNhT5bG1OOyjj56X29J/sIWQd1cMUAOBb3VHY1XusLfxZitMZnvuSTVz0z
637PjnDOB8w/PqEopfbbJIIU/eX2tUZYabRi2oDmW4yoIMJHzPJwCsFGJUxJm5fTPU1VB+4BEu24
YcZtaOMdYa05cexHeMKmUFncxVu3/2MVVxMOScI9EyJfnfUMHw/SRryTpCroD5/f335/WL3R3IgE
O06b1u2u6KdDrI90sDmpaa+UISBvW4hF+w3O9/EtxSa8Fic7TkIxIa2TfRJFyqwQOq/Ng4MvY/By
j9i2LfAQo9Y3EgUc6RZttMmOLn1SERhlVszW6nM3NoC4tSRP9IpMcs6TAcESnCmN8FfZNTTLi6d3
Z75PrcZjkAIwzTPCetc7Am3/bRUkKbS5WKYMo0dBSU/4AZJAK8NOBFniRIBT5Y3Q03LtFQH8K3aA
sE+GGN4g1DEsfv5IyTc6RzVYIkBWMeoAK6LWxecRVVAxDFShYMoLK5zCMwTghoD6c0NkPWukbx2M
/Afl8jaRWKGclARxXy5gIJuPcx13NYlp1zuW3RHOVsXg+fgy3GNihCZWQPoiprNpXmAI9hJ4hGQ1
HbHP40cdD/0GOIyyCdZMu+Lc7QOesSotHWmVMIDzJDo/f/uaHF74vAUtku13x9b5zKcKAAt8a/3j
nL3rerkLDjPJCFrJ1UXmtVCExLLG6SqZbCTNxIu1YayEaqZ6S56/W8Ds9o6WfJyAvdEcsC/C/NAg
RVUKlGo28RJW+7oyeHKOrJ7cYGLo80i447De86iG8ZBcv+oi9mLQpMvkX7HZQRCpEztE+aVXCew6
0ZPe5Nd8dsKHn92FMWv31k3s1lWySNaAaK4Qmf2Z86Sbfyf28zLIvstks+XR/P7lmEOLojL/50vA
8XQLzlGLZTgWH5TS5tSChfU3aKUwvj0U4+ZJSVHN4tbRCYqIjeZoG0I1sTVHoUgQuQp9lHcR1qhM
puC0uAqtQFnPPkmp8kNsWKcsKnuI2XvOu1lKZ0r5+7PZqPwv8E0OBEEUNfas+B3vgXZTT/0NCka0
oUm0zvm4X4DUUr9+4OYAJQcQ/CMi98ec+ZhMURgvlFfFtB+0CjzyqZ1SmMvK9mkB8lrshkGHG8t3
DF8H3lK+2Ji6GY4oTE9eB3BV3Hlzoflea3avl+3+TbbgaU+P5qoR8UYCYsx6LjdJo8OnFKc7nDeK
KpO7vCl4GS2j93x5vr5e11qgU6g7lekXIg14lD40pL2N6FkxBgJUu9QyWhF+MgjYNBqiRlFkOqhY
ypTg9pOwLDCODfW5JghQsnmDHpVeEqni6AIU9OdyZJk09oSBs5Pc7vkypYadiXZTS+1Yr9uUxnJG
9zdS7tOfnZ6GKcCMON+8OIYhX6lp7M4yu+0Hyuiz4/ULqi+foiLHI1pcniGi+9CYnFlPbPljC1T5
OgUw+UqxT43COAGMR/Jd5Emzxk0n45PxKYyTHqKFUI7f/tNTZu6Qq4111SlpBFfRZ8j/Ay3A9Bfr
kKromJGQF4xcMMjpcxABQiboRBvnhcJrsa/4tvkJW6Dd91iz3xhhFwU1WXRSgZG/JF7OjuHYm5tN
q3FHO///Cl7qhBcMJGvVcJRITmogLAkr4h0Rjll5bDJGFZ/Wi/ho9d38tvI6id5+zOOYcoQyCrh5
ZqZYixI8JYCIRVu0tj/B05+YCKBtOGMhTj1AxFrVuEFGM0jvcAk7PqSoYHGlkGrxqrH7v4JF1O3h
FGJ8VQQ4stNZQbc6h94wQjQc3tNM4NZ5Z9ba8O3B9mMkqdmAXQ1Xipub5PMPtR7QA8gwidu0ktFF
t/IfJWPw/t+RiFhLwQSda+hixvJMbgY3wnKYhOsn8ZQUejwerjOnQ4kQ6rMd2fszknDjw0dU5zMi
yc4Ssiw1RYkZn1Zgpll0koS+PJ4Z5+efnlZd86uhdSTznMkEWU4uUVNK9EexMVrDJb+H7Q2L3f6a
8J0znCZvvoWXzTILqVRgvYSN6midhMwYReigOQlIOcQ8N9wfcv4D6WJSPO35LnqGvoHYYTqJc13l
DCWKX7kVCqZ0f+LvwCnkfTy0qSeXMlwW5+xK7LwKXEcFMMYH/6BJo/Ly1+UJZv7ttyx2eZKVlbpA
/6f1jYVfJ1P7DReArXvNg+js5YfTPVLo2xBZEAvFkWB84MSaGRyFpbIzctcPZ4uxOgOKI0Awoq4H
joXw98ogFKz6rasmyOYT5sy4TeRfajZb7BKxjBbbi6X3/UawsC/cnYlXvK6LLdEElGuZzCpRP05h
DEgxbsNqUyP9m6zGCgNe2Q3UgiCCGEDV1I2OJIQk05ysaX5hCNQOWsftETUKuIX9huLXtHHBZgtN
yW9ogcxo6tPD5WD618nJGT4Ve+jGb02TGVldXYIzRNGCpX2sv0jrINTdF+w82BA35+80jCOeuPV+
SpNp1ug6BwqAjuaDzKmSqYREHloIMfJVSx4sBqJ/AzAsIcvdfDZNSksR+M4sITnQjMyGoAA52Gtq
VecYg6Ntg1p/vsauL7NPOVCMzjdJR3iWP7xCLrj28ntZXxUGRnbEpHuv1un10gnpoOErYkgcdUnv
n8aPkf5ZoSwR3sPH9O3OUBgXA84+Rk4G3squQlj+ugNqP93sQSmqXacMvAma4cgQ10a7tyzVQGDs
Gc7THEZfiN2EXFcp2KojA8pK0AfMsQnK2EZJXnRAbHGdo9Pcf/h9EZNq0K3IQ95NzeT2YQgZeQ8Q
IQWwqYK/NvRaMqMhgvR9gqBAKJQfhGcHbDL9SWzWIYrEn4wjTomkAmoifyU6F554QdOV5Molccxl
6GzD1hNjdvrd0hdBsuwIb97RUFY0D8YXimDMMf3tSPqmizCKOSNXqFw0MUJzTzCbP7J+RZKdKv92
jOBsiUqTILEIJ/GhJR84l77JDei7C7D19U9McQP1IvDSw9jJOWB7UyrtywpDT3PQq1p0Tdf4y/3J
mNbTFRD6mGivmmxiXyh+ld3yMalLzLo1ynBaygJabKaMqnDRzNgU5J/l9UYjjmiGhHmvHFzB4Q6K
+u38Ch4ECf1VbEJwrMgqQgBKFUFMEoJIIYQKePJt5pavaWyQ2Grl7zad5vzhXW55k4IefNOk7CPW
ozQ1va17vibfL9V4i8Ley19aekuZFKeXqwBX+cIlNxR7StPsuSg4xJSOsu1DqLiKVf56MIS2156+
lRBTBac86Dl1IpQQM3s9scAEVcv1Q0Y1OQken473NPsz8K2AJih6XHHggJE7Ii5PwaR3VFb1YaeP
IlnVGY4sFaVG7NGGCMG2LFVZD7pCSMBNDKXRGBYE0PJQ5IV4bzFOWwd/DkuZ/aEDX47c1hbhosmG
d3XyF7UqE/VIsXXVAjFbgQCzV+uIISdPtFNsCKM46BgKWATWnakXCVzn49f5I9u+7R8RhqTIzECC
5FCNYjiG5zSm/owct1E4JCsyfa2ACVdO1GW/oJgdY8HKNu90uwQCIxGzNun5FnPCAGAsCOEnESlb
TJ1YT/QR1KcV+obzv5ahKVHPl01iFeN2qScC+P5hQ3yqrigSDvbdHZvpE4h1NY3kbqXcR7F2zxWI
zZ74k2Bgf7tWBzYhPElxQWGA86Ueg93oJXIou9FSvHuX3+EVd7ZPbtkpLv0qeazN+kz7yEuJG2su
min97Sk5s5Fc1YEjcaCAyXcbiVLoaXWi0F2mzkhKJO2TUSukdUEj+SssTFSZH+C4AU5aplqyNdzN
ACI9ZMsiveolVZ03NyE5AEKEK/7BkqTrhDpiu8QTlSIlyz0xJcbK4/WnIpwvGVVf1OTSsyD/d56o
3u4jpKE2ZtDdNCjewjKNnBPLawMh32SHvuyrz+jXtAPJ9cQcGh++R+wtNcfQJ4IP/PAnAYgIM9h6
d8Dr9lTadKHvKy7YxevxGwiqJSczZLxC/3jbPDVojeVq8HVC5mKXCSm3RVGi9ZYrvUAvGtSvt+5x
Trt2KPIbuKV42E3ToHUz5W3KH3/0o9PaC6gWpVbjRtZaDxAYAxzp7dwzf+YrRX4GoiR8EMACgu3v
zWXhEn0khRJlcaE9uUvrj9+V/UX0K3GFxBqE7gI4/l7LzOLLroaNy9WNP6EptXzhydMXbPQHpDcB
6PptNo+xdyFnw6oov2+xNMCmoIACMCr+/1lcG8jnfuX8g+BwH/WnPgW40RrBvtZxlKEb0YW/z2db
PU5Jufwfd/+kdLPq6AZM7sFLxxKurlsqSBZY/r9hZS3iDb/eJIxFtfUo9AI+hztdEvHk78rw9vO1
Rz3TvcJCyUL+k0NLPfXGODKMtdllNQ3X+4sHwHxxMHPm8kztAx6PLVjPV1C4ikfrOsTYjZYU+5+f
J1zFxHO2VE0YxubPYshaZ0IEkoTzVBgNAxUDX3DUNbbeFyFN/GjpuFcYv4aKJtoEr8UHYtr633V2
mlyDxWHS2qq25Rjg22pKt96AKGpzkqBr+H4dxVW68fekLFKVt+K+PlDOyC7B1/I6j/zsv20WbKhB
g4czIq2Khbn6VVa2bKojhmnA6UB9CQBN+d+L9HQnzvNVEXIpPSRMXHcfnCldRC4L8ephtXZ40/hq
K6a7Khy5YLSMCeypkoprO1nHW+08bMd57ZF2p9gi3QWa5Ukqz2oOa8msBvGIq0ldI0HTKxb0R8x+
bpcOz81dNJRKHaLGEOuUG+zT4QGuNKBZOiFCMcX5LXgyrEGjKT/LhWMV11cIKjgcbSigGhN19SyQ
fblEwvBISd8/pbnLarzv2IUZO/+CEEObiK22BSqwSEgOkGPBSaB2XXK03rS4IAV5a6qoChv83/ra
BlWBc2x8fMVTk+aCM1qa3f4hTaAeaQ3jLD0duIuRhKRCtFNr17Og4XctiMRdUja7BusUhRQctwIt
bzPGkf5aj9mHEU935iOLDnFKYgAPsx5wgFpdpmew2eDBezr9PrZRLMLqj4O135BZtbMZVTFoWpQw
WH5iXJL4WoFLE8jmpXcOtQvulR7UnKpptGtNk6pOyc4AowXoFAuT9wHCs+snOJtuP1GD2B1hjOkN
pzUNhG/Od6cSNr0Ppv1Ojft1x+Dt0uUbnIr4/PNXn/Yp5aiv8KtVKjzPZYUEt5J/BxX7FA1zzzz1
hJIPH+RXOrXeTQzlu1Y4DOIssdEaQYCg19ENYgrEU9xzD+z6vvFbyQc1tvEO13VR7yjozcfkqRHQ
0cfpu/KEYWgdtt77PZ6Am7qwArvJT/99pV6Y8lk55NlfRX+y7ekQIYq/JhZPyC87F370gvSebfCY
pf237iMN2orjvAAInTK9rwiPW1vErzjtgn1Tilh2aHc4lMrtC79yd6keinekjJ1EBcOQLM2M3ARt
VQLH04/OuL8B6+mPbf83Psseb9sh8Ibk0357Cm1IlfAX/fkgLrKV9RiCTUMzAheoWAhASCIBUCVJ
vW64iGGtTUUf68fvhlQWE51U2wXQnTM8rgbgeffx/HxA/BYUF3xM/ZMlhrTyKlEtR/mHWSnZRsDa
lUv9TTbrl/q2RyQB+iJLiWgt41rP6ngdnrwzshfBe1I0EbW7W4/HDkHd4olpszfpTOZXEMYZs8Tn
nDGt5bwqXGxz4pf93QyMB3uoyt2UMKNnW9HlFJoh3z8laNNkahlCC9Tgg0+DqXq3SjANXdqaORf7
krAOZNbpGMNve+oeiR7V/gnMqWxdrM5vM1YEOaePMRnFBeUgBfzjZ4m5ihopENzXC0QR+csxteBH
gBx9t0uYTv3AyqwJuNiBr/fvgSmCVuL/h8twlKBNDOKIvetqdBuSDlh7ee32pqkS7aiUTaWbqZrt
b5yxxVFQ1nOam9Hh0ccxDbRxSvAMV91E/NO+L+Kvvbw6weHkFmqJxlxx7jq7uPArHkaCZAKNTIDj
K/+T2lqILI+VbPwBIGbQyCVBhdvMXbdDr+NtpVk/h9K9yojZJ7Ve7TDkZ1eDO8dV5dDQeZrCloAn
mo5xnRTrcuReem9nO43m7l7OYI+UG4OEgN1MJCQL4SwaYrQzX7ABJby4A4bgmadrAW0iptoPDgi4
W7fKa/ZrU8CiCU8BTXSIGYYsmdh7PLWyuoC4FUdJ64ddCkquZaqHsOV/lKdS/B9pK4Rn8mpzm5qw
wWXoV6eS8ePCixEfPOwefbNzrhkeE+1dpC7aZffeeYOwMeiBGbUcYYcsbJUcFQ0trWZhzUhKSAc4
fckETnAhDrqTZhLwypEV5sqUZbC3RK6NWnXhgr6ORHGzk4sq6eK+stmTWvtlJRgXH9O12t8FVfAI
U6FR6iQV/iWWFcJrStzM1+xsu60Rupo28VFdYG3FSbi7j5lnEOMxO4Wv8IXP/D4xZB4XghQb4NYn
Oc5xdAAfHtcrRxL//sECbT3qZS/voL5q0oWQzA9Woq63KCnPakdH1dK540vGYfi6YLBLir8i7vJ0
9DIK1hjygMsyH4ZAQxxztt9JMGq8siQCkDs7M4hshiu3VBuFC31VG1sXuxe6UdPmQ32fiCRdVjaR
RTL3LagTVSziTn2NxPHaj68RusPCv0w1HgKXYoa9OcyAA3VHHmQsFShkmoalHgg4c2vuOoto8YVp
i/YIXv4U7cwJ3G3NV+UvTuG2NNZcnwDx0E70xLhlr1m6YydYDgCRPZktELE8nvIMZB+SZuMZaqTx
JWBvRsSdNmeS8BffXG2gDePv9HQ0GmuJEkVr+j7ekSatrftSz5G4LMXFXLBNMJlsX8pTedDc7NZ/
6eC8iVvCh153+ayYSay8JInbwWNTUuU3T8TEWFyrVpZbKnJjdESFI7at2q5l7xYmkyoXBv7RPnY4
BLwUiF1Y4D3zrM0XzEmPACyyZ2yVqsoQJrXycVNJGlb5Sge0PQn3DKfvZty1cw+AXMg2ZCOQqfqs
s+f3h7NXF8cEY6FS4g1Dt3D/8M5adLNDplihpJ7ollHu1r23zwvDL7gXS33ObHrMb3I5ENZMfeSI
6GFJMFaAS7SMCx+C+QLOxfM77ZXY13HDJCk490SN77lem29pr7DsJ94YaA82K5mmsBWo//B/SWkq
qp6UGGS5pFiy8wavI/oB/MLk6wbTjqqJNrggdJFVICS1rMBc4TRbVRFXXTl1l7W9c1yhe85/fbHf
zEi7hB+aZ6zkt0JQDaV/jaPCAHHPk8/qVtnX3XBDqHN5NtAOITLefZZi7YU/gljZP5AqvweEtZh8
sbBOwWukALBHOw2W/KJ+yW8B0GW/USlqNwFLq6QyN/QrIXLbuBSGuMqw+qpkCpo5yk/DRUJ/FWtI
6ByPVxad3AL4QsdRcpIMMnXBkEyTuQz/rhLabtpx9H50poVbjd5Kg1oYeLUyWyhUAzfHY09WHfaj
MK2aqnwlsR4blZHrYh9Xsok6Pj+raMInwypjKH5o8xfeARBx+kCDyPCBBc0vgc9fdAlf5vuXIYni
C91HkRlzDXS+iQyN0RwdzCj9gyo8E1hDRjecwlfssHaB9Z10DnrNp7ZVHD9rpYHs9pWQrLiXwzoN
PNRYKOACNY4qYj0MgrzeBa0STai4B+ETC51/+m//UBII6FUaYl/RQk8sHzss4/pAI/8XCgbQFVGs
NCdstZM888hIDhIY7W5cP35yb451EC/xdZoNrWf0proFGFYG7tKq2T6k6cEgJIZ83neLYZtLAIHG
UlkUvpcMcr+lu6tGSJNlKSVF60Jps7sO0VK+ayEZRWXW6cPU7gfS++sZQTeaGExolCdqIB2+a2DE
vyocKxgY5pcf5SYFt66VW2CgiHDpwakGm++yYMH0egT28L4vfy36kB3P9KKBp3sapLrVU+GMk7GV
v1rqXdqVwgJcXd1YIog9ebXlHVIghwRqBoN3Y6OTBBQqElG5aFFZaG4Ha5R1QQJAZgKIx5FzBVy7
1WrUtThGOehtDsRUKYF7jd4CtBbYWbOuL6jeuAzwlXcppQGbpQLeALvdBKz6757tsBG0Q5FBmgxa
hIUmG2SbOCL0ARoyhNAuU9pobJF/fUZAhMUKk2gm8pA0ATZDk5scyBogPbZj7Jn1fGaGZV3hiG4F
Qg84hJUV07uhf1WoFPA8TqDFyVCjFXWDuYSYrbVxPgbLSXEGGaqzseYdMYGMrXzYSN7ihQE4v6T6
tAP1o4whSonGND/k0O2DYkIT6j/iNxtNrUfWN9vApx0Kbzfd3y1yNeWpLzQdhb/eRMbrph1uiXKr
I3AEqNTqVrhXWFlxvBqv6/NurG53votXZpXF3fRIUMpaJSsphhYsnfdkTDNfFll4m1u82R66kZff
VqixB7l/hbR95KQ+JhPY6HVnMYT/KBwYkifhiHJ+i1YuQ7Nlbs46FeoimeDXvMkQuRODQkyfoZVV
AqHsM7GGB0Q4p6IuXKuREF+/oK9BI2huNsJ+3p+7ZiOUjx2qYNjOoEeg5IfTnRH2Yt8Crja/GlCo
rVp7Ql4UDQPfTPDOiLeFhMZQsyaDdARSXrW8hjKNaXx+oO3XODLzUYZH72Z0G1IqWAQBwYoeVRY+
O4HOdArQ3qV0Elb8xCw9QivKaEEcyECkXn8QDI3ctHitjynp9W0BPRHkrt973JNOnrAhE7Z/vp43
c0oc5aIS1/ZddjFyZX5X0DfXWFf7kmkSHtWVTiW17aK51t+E45JMpVOn83A8wP5pwRN1sLK3j0HK
2dMW8T9wcGQeNf++KuiNbSwhyY0v3cEdyLenJfEX1iKFOwIScYwaqA7IRZF/Uih1CH8q+G1NqHTN
y8dNqpSgLOmPouIeX6oqdCCkeg+1M5VdPQsNNF4aD4wgNClNXV4YZEwgt3qQ3Ugu+rgoruC0/L8Y
/sC1LXK6FKysBUvqbAYb/seXe9dk81kuY09lcZwMQwCksVYWYR2AwLafggNAXqpEQc9GfPvZiRso
q+fPWN9E3j/g274DloUyhQ+lMY+NyURoJWhHr54ie0eedXPWHz047p1bl3cOXcuwQRWDjRP5+iix
rRzpEXGRfXC37aatSDSnsrH6YEBOFkC7kD0/G9arJsQf+PJhTy7r+bLtAHih+zNYI6SF/9WbtXKm
fNUf3LfMQEbxp1pG4NWN9w7m+AuJHK/mApkRR1dqbFxQXL2BJ/mH5Yypzd28Ip91azh2JEQuU56Y
b5mQt7Iz3Y4NB0YG+jwwBdJwp7eKA8oE77NWf+O6dFfJCXD1AzEZ2lXJc2dvtgMvWtC6Y9t4D30F
xfeOwFhk2H3JmShaAvU/vaWuOjVe/2hQuwdbxVey1ExBEa/sBekW12qEb7t3WuBqJyWSZSsXMIoB
cYbE+xS2QzecR0OSd7FGl7v0lUY+OVtimlDvH9/0IHH/SV9NS8BYnYAPXYA4oRneB+DDlyaAx8ea
SHTISMkhXiM1/RcD8hIY92thgkExLUlu779J5xH8RmDn2kPNuxhunYZ9hcg4hHupuYHTkC8il25o
288pzjdpjrO9njXIOHL+C2xHLer6tyAeKDQVfYZ9rwXUAW3s92kK5L8T1dGFRqTFyDAWCjeu3p7x
UHo9UYotm0aj1yhhg4m8+YwvbdzTBeElIVlHY2/sPKiA5657Xno3D3jW8DPGJ8q+s1GWczf3bbKm
3D2+gehCXCGPI8cKuleCxZJz1WQ28S9C2GgVXNc/1EoSFFrinhai4ME7uvt0RwPqgAc/YTv+cX0Y
2MyxmAqXhlV0dBi6gP3wNfW/0GcCx+OpWgkoADtJ1j3AeMDzav405shGKlyme14yqhAewPn/rsuB
npfSEDqFhW86aY3WlH74spSW1Fm+cE5OFCqycYhotM/kUW6EUIsnNCiWpl0vg5rZr61TeNmf5/FG
jMsEmo7VDuZ+XAdCJR57l67MYi4bssdJ4KAuLbVzVI+jSOuwPKSTRM7nWNhdUS3Zy+dAFcUAmebk
an8jwuKWvfl6J+TVIM4496EZhHj1h3V7rvnqQ88DUEyFQxcFDDpfB9o0avvGnzSQwwJacqS9dXeE
hnF0eTNjSurFwiosIzh8jADYf1rE/LVM2DxbpM5bn2/GELVJSWDaTQJO76NefXyDuN0e8uhUtYcu
RSWXhQDMcDhlw1s7VBu22VDt2TEOOFAZQeso7bhhxYrLAWswm93yoKxFe88xjfLJMHGComTJv6bu
6nR7e9eVE1qJiZFL/FkcHb3U0k46R2kr41m23aIfOmggQOJJntQv9Vdk9gdRWnn8hWPmi31zVHwp
S7RE9ufHpLFHAt4ensxIWwkajldCDTzUFYu9ZSYr2tEARElGDBHAx4IPltXvWcBTeUetzzqw2KZq
/GNxoOiv/WQiLRRAohCiXx1iNbzs5z1vIkJa6lzqVSsEtT24Rgwq3me1p5F+zsaZzyROGCxmc0mS
UqqiGyYaBv1VQ2jwYNkSLXZh80sMbpqjGmu1EAdw2elSW3t4t8x7abzQ7Dd8Vm5jxWPOx1XLsoat
BHVIwNUJidNFTiZB7HzAfTFL6g71D+ijdvawNVrX2Iq4GJVihuN7McuPEv9g2eitsLT4E0t3nfti
zYm1GS+fsq7oFrRnshE+coijpfyOblA6WVM0KEcZsRrgVpPgzC+L6TXfk0U5cZVWEUw3Jl8wVGfm
JrTUBEPZ2AvDZ7U+EF8YewiinSPRLeEQXGW9h0H+pRYzOn3qVcniqx6GjB/J1OQsRI40ws9XwW4w
eFGQskcnJGarZBwp5E0pWf0z9u7B/40RBVD6v1G/UnhpErTfTc06cuVqr48n9nARF3iCzHYM9lNf
lHYuNoJU4+92+/bCz3yCOHDplUYbgi9y2/L/Iqjp52CIZI+0CPRFJpRJKaC5J6ekC6KFZ+lEr9Wu
QY6wIOFsdgqTYpT3szicPIAeXKS50q0UBK4oLV5f68e5fwPxu/WIUoWS1GNqbSFCej9IIZklwjwK
fzJVMF571XHEK2M6xMGqh0tWgrJ4bG3PlMDpXiQEP5dRw12n9ijXdlXxlS1WqEcPA5zftg4TyYbU
4DvhdovHGy9Pa9O98G4KKUmnf5i0pG1m8+nCKq7g16war7jnYm+vGiaLoetLR2bsNdyLyajECAVE
0TJJqlJBa1NqAVkW8dDZpJl1rRaewSMTj9NOSBpktfZNzf5AK+/+pFRlznMvEdeiVaEujDuTRXNT
O9PJpdhCtx+O6rjWt8qTwnAMgDu2k/AM8qooY1SBxlcf20wt0TulkqAiMyFf2XzDBiohdf3r63uh
d+HVBqY9AsHVByy1T7c1nUvQHu2+Y/ihvJG5iYNGxPDNEh6yzv0slPZmpcYZNVNrpmuRfSmqMie9
Kmvgt+F+enI3cqwJ87NsTsBNXc171mwJcqHEcxTZf9mjkllPxzBkxNm0ma0hRaZCewwxurnIvu5D
sWf0p3DfdTvVqMcwyE1oxcJ9WcqSsqlk08CA9DiA7Mt1R7LPQFWcLevrGNsK0GygY5NR2wSiQd80
0foFOMS0eCgFxN1zDEzpiO4FrVGwa3JgkmDIL97S+SpextX2jrrHVDrIC+/K+iqG55UB73PuUrsp
KhOpFs5D2uUPLrgBJNzXy91QHf6OqM2kgbBVZYBb6lLwx2Ci84prXbMhA6kg8PUBrr82G2N52TV9
1Cz9Z2Zvr2XYwgIpv2dq6ugGLyF9h0kNDIkMHIBkReyycgW5IJLfAN9RGh/9azWqV+3saaTBFgNK
3hlz1ti21WmcF0xJgK0mGNpEN5iYR52BlQobHoZ+hsHuJyfBiC3zD1d+peGS1GG9HG6yHTVdHNLH
exAV9Vz8fHG/XvJbXID8yqIRHYePplX6L728LNYPTnLf0F1Nll5C+7lvXKAd0vMUUF0qWSL+oYww
ZpfR7TCXyPHuKuB8fjr3S1l5otzgavbDSb5ZxHFZYKcMBDMnlfDD4VSqY8oPZTRgLhA55XOgseei
nCdms1ZsJ2ADShEkliWBhb0NXKETWi1TC3yiaQBltFhhEBRbHwCkOJhqQ0fNRvqq2hmJhKw1AtP6
o0hJ3JyhxfBz4kMYBbmEGUBlmAko1EGmo7rnbd3XtWSDGgrRRJuNgPCg9YsCc2/BNOqdAG9NMHn1
pbmDXe2kNze5KF3LEeJl/rPSTBgD2gPtQ9WxKCw5HTj4L/Ld+oN0pFBqJzsPq+wxS0Zbj5y7ZudS
vqO/YYrY9rXaH+RkXS6lag2IRwGsakm+OBJW+h1s4uaYSmpt8CLw1d8moMBdMD7ZCQzJjNl/N553
g5RnOF4EyackemUhq8mRwpb6eEP2ImIsQth+boS7Oja/ocmsEPQAugJ6QjzR1PptvK5/EWEv1yvp
2NOEV2w18Svg9c1rh7d0goec91jpP3H/F4+CBwQ6FtiMxjGPPLjM1DV8xmThrNGcDK76WTpXEBLw
daEvZ/x2MQQEv10eDNQpURLiYGdtsAYkdjf0UlUJQBUjCptt5Ieso+Zagza9yJjz72use3fGS3si
dfpq+kWPFmr3A82zOIbxVRpBuZbJWDZ+qMxkojALe1tgHr6mqv0yIyJP2dP/TbycxlMfl4qX/wpA
+SnLAxjWu5L7Yt3x7ogWkkiYl29OIokv3X/EU4qHj3Vw07eJJrXCMI3IYbtGh93NWJMzQHLz1NKl
Ho3KHFpIb2d9jWZ/HxLhwptky1ydui2+OfBRfYAB4UPxlbJFynfFKhHjgPGFMsI6Rcr47L9nb9j9
LhYl+66ajy9nscWzJnko8Mg72GsKCk96h7+pzFZ5o+rAXhuDpSHihfTG5/T9hd4DfNFDARoW3za+
G5oTgpSccmBtGRMngq6u7vQ/0HkqsAMRY2vaGzd6ufGuKsEUnu0nFyu4ywjLxpW6fEDDjQ5vQn+0
uy0XKDmRnjI0BF7aK5Wce6i8CZtBtIjyQR83zZyDZpRciFWPkKsIZiHGmN4543XIUEIXjVnNpFek
h204g7VR3h3okAN7Q5VqlqdmNsSi5KKTJvdYoBD8LAUCRdPy5TBHG7qviQ4oBfxGFIVgezMhXjlU
mf7R6LTXN4bx8b1uEDIXx9B2s2ou7I12LxNvI+KS+4wsA5KtFxdN/Ba3B9sKqWdtSGwAtgxcGy2L
93E2g2FTtT6Hdju9xW5SB1FwvMtkp+t9S/mbQpN2O4xXhEI8kLVSO06/nTPRUR/PJg6ZIq/mrzQe
E+ssVHms25y5AnG5VBpnFgAnd9c5/v7HODv8o3c/5Pc/EromGo2lHdHoA0vUwbNvX4Tb/aWftUUk
tktSTV/sAfoTlTadzfty39Y337+kzjdqoCgjZCSqz8aY8E3oG1Rklf5aQ0wtbNrVvGYYbeNJg1b1
+xa+pm4N33Pgy3dMnIZxEYeS7OPdKenSLZMdmqxVc15sqlSmdH74Jz3HPtOvGS2+7QwP6w8hxfOy
XH6T5ucbfsNSG/oZ6NRf8srbzwQc918dDtjMt9mOP+vRC8G7jWQDQn5TgOp6Qhimfl5DpsvGaiQa
areLdhq4LsFZZ3X5gc926kEKblD3I+/tUw0aNmhdc1m74wDecrlkOTqlXFrDnqquKFfyfUuvWd2K
rwcDYZq/e3L8HvmQB8S6+BLBx4JcHOe+dUeOJfLHdM4CVWTPyyIrpt9JB/oneKekjG99K2f2jGYe
NRv5e/vcVyK7LX13UFjT07A7pcsNtanBb0dsTXUYIrn8NILEOk5q7u6gRRKl0NzUN35E7RSDBM1z
c0WPuhBMxebA9ODRmUJYjfUPFj1XVi44DbNwq6pmlLdsMO3he8V0lgwB11pjJZ0PXNco0B4Co9Mq
AYEj/ymuD9TuccqR0TnovBZqX6I+PYbce0y6jkmaewegQfE4UJ3yft+E7G4EAV5HYtakSciB+LVb
r+ZF9aPi/yAhb+3+7kABZKsvti+8/nZuESQvOVCHfCmRjE+yv9qjL9AXVHoFmxH3abRQdj0IiNgc
g34NWh3hK6fhVsVBElkLmYkPZvPP2HN2EwjqkoN8TTH8A/mTbsZWXb4BpBVZWPO80tguQNfGNLZJ
5rcA0Ku0j0Tm4ZnYFQwdjZqGwiBWDL4fZztlaBouIp5RJnLn3FQ18eq3obERjCiJAmczcerHOhLR
ZA7tq/LDSsnAduCwXFvI08sAiy61bB9kL/Z7yy6SDxS33RPNKFutWla2OPwgcZFleoQaTby7r0ZS
yaairBiC9OyjZ4aAXH7Ly3KfkxUV5jO7bm/yX0ljqYg/hhakubnndwDjrG5Ru5FZWro3l7P/kQ6m
yU2KdmcgETjAWySmkYbbMMqrazipCtSTlsSVriJvHL179QtvpcZzMVzrH38VXlUbCDW7Fjg4Q8s+
rwnpqYq02JnCEMrMFBTNoA0LlyD8E0JjDIUr9CUZ1AJ9jEAgx7sTJX5z3gVea/mhJJ45590Kk2RB
eSeZfM5CSn9nBn77guS/xHLHQhPsb6TNJnKjFndrABcS5MKCSRKeU3/pWm4KUMTsqwLonDNVABn7
DjDtaVfF+1po+8R4InT1OwRShWDiYihpWNbJ14D1cc3wfBOIKYA/3Hnj+ws/+Mj0ex3ZjqrDsTN+
jM7RAvf+1C6Uyzh2dppklDYCxQ209QTYtFbobtK6QTlF3CuvSljW8MtEshVMHN8mt9eIEBAZWOcJ
rCHKBKTJTeY7BqXDz9eXjum52IaudKaMaDvvfPd53L8YyUC0qg815e4SSfMDEap6aLLhTfSSRepR
VIFFqc3UwvCT+yrdHAi8lO/BTrG/AsdMObx2AZ+UGl/fH9Beix3muYE5eruc/SwRLMMKl15h2K+s
koHhDrHNsUuLT3pe9CpAmjAB6i33DrVTArJbRUSPDqlrKO0l2PGOR9YiN8jis3TbP7GBt1EuLJW3
kCJTEDu5HiYLrWFZ+tDlje4WIy3W+1dvXCV6ly/AN0XxR7l8J0oV84JD0qZU/FrvIA7oj3YVcnDu
IkCKH2b6jKmMmhvVpbnkwLM4YFFxVO7B9tb9mEpTHKDdULyw/UR0gbySPulRhY9vV3uStNgbStJN
1TiE+Xy9ZrZp/j59OEa2nL0aAsLMW4tgoONpCUQcZLNMXFWH1uNRjL0FajkeC6vhvHowtCA6S0+L
aVD8LlDOuSogX/qW4vx1QuoD0H9m86AyRb8/eoOz9Fn8FcmbG5npftfMYNXjdK6StWXyBPeppeef
Q5h3DeemoYFJm0wbKERnQXKXWPhvE5q1BgEGVCs+Tn0100fIkioVD39V0awo8SYgN8p8pDG4Jf9Z
7K7uEw+MpYxWUpOUDJYWqqzFbApfk9MHZCoYz/nMGg/o5oiKoipJzIfns98fqQtuYoG6eZEbtOtT
s8sjBnmDa+/CJVTPfDVRogUHL+AnPF9/Sj8oAQ5WrP6YY4hQPRsjQBalzYXiS7YBeh8pKkYmMvnt
bUAGULqb7Hl26h1hzsSVPM9tFcGris1VPGsp88Smik0U2V9j913C0VRLCQnL8VS0Pa/J4T3YInh0
k/PU+ztSRx2T9wNMG4tJ3U20UUtevgbZvv9+VvvCqhjYGObt81nwB/jpvUSWy9sMwwh5aw9wxwvU
uUTLqnngsplmayjuFu4KVvV7dmp6IXRF6+aytNz8eFubKvU7p7sIXPho17Sp6Ls+3GOP5RC5CDgs
baXq3M2gULRJ6PmHlYbJXnHStiPc/YsGUgalVwTpsgx3MJ3p5z9DB7Z76oPVKvi0iI32D5f2JsXR
IOtAK/la0FYTOKylXgijPlvuq89dcMtHQkjvQxpLTPNwiYoJuJ0HcZDh8t1wN4ARP4tW9e3j/0zp
2eEQIChT5hezjKNDEKwu7dl+k8CYOanZQIAnbd3Wy4IbDDPRe1WyeOnOq/K4MtHqFcPvC9tp4QBk
+H/QZIMvLaevTeilSi3zST1dSfHWBfltit3fq0GKDG+PpzSLPY3/GgFePVlYR0pPPdw/2J3IK5Pt
i64aDPjrOdrzoXcN6LEm3SkEqdzu2ARWOa9MLOrrkqxMyArBwGGve1vhQZU3Zf9h2ri+uFnSE27u
pSBy4xNpoGa+QUuPjOZCQVccQWzkQGUD/d5j3qB/QyHIGyDrbZtImfzpOJcAR2iFaIaJ6jzYT/5e
iDgLn7Z4GsKQTHzC5P9Ns/QA3NADhVL641CziBiwYGua9J+/slZl7C/RAhOyIkOYkbNPt1+OvNPr
ATVMDRl81LDEk9lca7VRM+iNVrkT9Enr5zhNcEt+ayV6WeoPSyBJIAI3sryoDsX/0AXo7mx94Wro
h1FUeFuV5xS/TDeK11ScjR9J23aOEnDdTkdq4rbvSposRl1ldrPWLOBI7G60k3Ofd3s2kb3FUpmo
DYo7nK0Q3qH7FqPFIFF7exElaLKt8Zlm/BvR9UEm+FHnw5p4lhZQe1zQ1/dXeoQcH7A2k2ree4GP
mk1rG05UHlCcenv9PnawazycbGH2aQ84d7IK3YReEvObosJN4I2TIIxxosIDqBmdbR/7d2/Z5owG
+3CWqJWPjZHRA1IKr0u0a9W1QfOErjsY6L21RcvKDZQV9fGqPkuG5Zi7cU5lJ4vaXs7Vx0njaZwo
RQrQ7OcDWbCWSxa84vBb2n+1CysR7s4xHOdOnU/TruYg7YrTBCo/GlWa3DJNSKrSIq5w2NeWJ1Ka
mWQuOE21Sw39SI7o3Kqdtll2Sg/FeX1ESUfV/+g9u6OCWsSmkQzoSeYQJIGmqYlMzHhkmdTtpnTQ
lWdjxSahnRsAV/5AY6hlH1bHEmW1ytFJf3zkH4dKY8Ta6kL+VceKPTAmNouuBb9lowJ/dQa3v3MK
FgtRPgk5nJ9FCWfRz0LPk6HP8dV+DAAWbhmN6tJ4rBMkB6d81WGyVGHZEOr60w7JmuRbTWFmhIXh
5+Ivg+B/FPAk3JMhgeJZnTyqbx8S0tFwrgKTqkNlAgI9NRtfrzKVgPuUrVSTgvGrVql9WUDqxnfE
I8V8Q2vqPL6M81O1Diau915mZJAK4wx4YrZOE705dKqx6Zbm9ysAekDhmPT3JPj6lBRVRyGj4HGS
ysWG1yIgqHcxtMN7ovcv3YuGPeOkBSDy1fBbn83KU1v9q/KIm3gDMZ5I+LJJVxLOMN41k+Rx615K
GNkF7xtVuuo7nfociFgxTIhzxEnJKqq8ZO4qkPElvWKpedQB/JEpaNz0dMPGhvR3IiplsOYFJrUz
EP0yD/D18HL5oaPMl8qIHPDE5Qu4iCkvxemMPUMomvOwYBGpUalxbQ0pofTWlLbN4QKFW/lxiK/U
+HfSzuWQLC/Mpl/X8oQcCtRz0wBBdXFit81FcBqaqUW3LbNsR+cN0s58shTFSrqzSuh4ITZt3N59
b3Efp68nD7nhyMntxAddIC5NsWKB2Er6xHHTse0FHvnG3SyAp8feK6Uf2r0MshyeWhy9RS2KUCCI
VxqhVFE/UzeqWFSwOnQUEtsO6JhY0HhOMx5FDowyN8UpsDli6/4hVoARG6DmkqrtRf1H1MBH+3w1
9KXhC2/dA0q/eD+qkTAhuAN8oyOp7riK5G4k9H+ny2FPsY2dWOLfUkSjDxHte6wzlIw8qPbXDDTc
ctDqGr6RJ0pN5MjFnWWYsn47qNV2ebdphUXlI+J5nXAI0tm5AxCMcL/8N6LzUpAgWq/zOzEqZsvf
JNXtIHEXEdP1dZU1bhXuQbYpHxistz+TBGVwHyHKOk03+p8GZjGgkk6n87nrvQOMjhEi+5hEEM7a
TFyXTNFqZGGMtTuiEH0UXJnmiV7lpmqCk4c4gaI5/430xNjFjb3hR4FIx7jYNHysqAsM4yABrYL7
nMbhBChp5b9s22ckQsyGFGqgztj/0y0Hzcz4wjzyL6MLah4NpEHYdA431YDXB2ANshs3uGW4bQwt
bdklHL9avNvpaQM3F67d1DB78RLAXFIv2gBybf00r2UjJOTxiPLRgVyKclnFN6fhOgbzPhzZpnlk
Uv5+tcMWk6CZARxfD+qsoNvvQFGzPvQqW1iCVhtW9CW2OcJywzn+tE6vtQ1Xe/80ifX51IAFimWl
ZsrtNVe4odj51loIBpwfkIKycfOQWiXsOfKmf7MKKEmrq3RpcW5H9T4eVJLhwcqgJp7YpJHXy47K
QiBKAEoTEU0DQ8iXqOcd3Kjx3iL2wV25NFtWVRUsRXEqw3eSVI7ann8Krw6Ae6Oc8XsBjnk9Q4Cp
zskEsPXi698SNiy3JnWrjwCImSeF4FzN069Xlr/BmjzCyq37znID5zDXRxe9X30lAsLYMU5Ty7Nl
4REnwcaANM1gKpu5sY2PswkwdiY+baXwl8tE7izl1jx5VH58rONRps9H20UHzhvETs+GP3FapIcg
/eiDBGBJCoO872DufEch4+q1kBEy3cFexptm7sBIRowF6h+Qkr0SDSxKZrvq/x2IrEleZf4gHClN
q7czjpP0+kxRSiEs0122clHz6Ehuni6hA09b0wTGFX/R/Kl9hBYm3HPmkel9w01z2pO/483toX4H
FPV2R2BZp/t6G95qbqKBZ8KI3ZF2jsmaS3JZmmK7WVNQWTBRs5GFAMeXGt1V3T1+AwANQyWJsdzO
Z6UMr7wu61CXlYg2O4K47j95ew/AdV3bQLNsbE0OxUt/Zd6zkA8vWbSerOlOIXEORd56GO2qBffB
cpgMzcIVrmjWH1JycJ302+MCxQvWADB24irEm3rb+hSWd5gXK6ibcaDqlgI5DNEMDl6ojLqQC9zV
7iMOoQFUbmL37HAY07Wh9J/kTG7r10Twy2A8kXZ0hbG07UvhripapGnvGbey14ZV4QYI/sPdAR+d
fkkxXubWuPr80W2NCqcDGm4ylqtw9mSVEpdhrww8X22+dlSqBZDpffOOWiYplhRRyhgXSHResL1L
NuDm+Qt1E0wgpdNxV8ho+c2xWQMu1euEeC9rIJqQNcueuGI2M5Nc+vc9JLkkytmemdGD3CVsHvvu
gcbev6EgRoxZ5KB5GGTCT7Ta3a0Pw8l+sSKHLqP4H5z2ABZK8mnhIeFQPDieKhVs28NibWSuO8B8
oTj6vGIk//Y1bW7gKta1T+G7NM7IB1XlftI31wP85IHF2f+gE2CRbljaPrllIPicwgLwTDxEZIeN
J2RCpTyiPLoGrUGqEi1Te1YWxHa3Z5s0d1iuH+98TGIjFgCmc3o62UvFNRhVNyIU9xeItgTnIzUl
u74mTLHiRVOdOrveTGjp2UDTD4qthsgAakHo97a9Z79N2Q14zrPJkivUkbe3UWvKD6f5S2B4CNQe
kJeNbvg1Qo/N9N4tsk4AzdlJVDW9zSQsNFNagfNxEoFcRsh7TJL5Xyzlczti+bC56IC6NHv7QzBn
iz9DhXxkW3epan9tSLuasjKI63FQsQilttUxQeM0UlCU7ASyDSKFZSjBb0G51hV7XQCvJeJ0NYPp
Am1nxC4fTQBYdR8YUG9AZ00gk5r5g3RJbIDgzct0iFUGLgVN9deYS9HiPdjT7nqPMLuz18LymZsR
ZnMXpqGuVo4tLoM9mIeWXXxnYt/GP2grWs1mFLRJ4WH8599meuTLeSGTk0xP6ZxDx6tAUjxHnn+9
SvgHvmDtKakSC0WZI4E4RKOdTHIDFsMDxBT1smGkgVIc+/DwIexF2YvxN0vtdiOYM8IqJQ846hZ2
DERW4hRcAw9PdHZM/E56AJPF85kHhquPZ/VwT1buuhWtcYGXvnx1BXOhnQZrBV6fTYExCiYIh8Q2
Hf1m9CLn2YNxd5SWwtQ9BnKi7YOVzJJokafOwZQZ8jUgTWWKv2Ba/qUhifJbN0Q1wM6TGqffV8Zp
oltIjNmOp3oMWgdhdE2sM8kq9cppG42/yQ2oOYVTFcsPpaoQsXSdc29RtHHmENNfdFC6AqGXOIT4
fibFkIeR9QHf4IvnqMY++7t/EtzqR/NzBxeZgG19gd8D4H0G8i5/MKcsy1aKpZA0T3b2lGHyODOE
5m1QT8IFDYucrQVbbOpjYeD1wnOTfKKO978msz+JydDSNvwFeNjydJUByt/UPwZrjLs8j4DD5s+y
nzCE9F/oImtaMCBoqYMdzrfxPo2+oQFD5GXjh+M+j1oLpZw0S7NNKkF1ReO/+Iqg8QqSCgjvG7V0
L+mokEGxJ4qD6f2EmUwqUiqT1ZmTn6MUjobXIdH60nASogUPwRRbe1CoyRgT/6FD7SFWBtYXzutL
LIGZLYR5jRrUOMjgtG5gz+xtixecVm9jjYpriVQHq333BDt0hPb4/GvFEa/pXxGAuZ3eYFLRe3fH
okv2cMcspjLSjBTTMuq/tIgQMP1LM2Taw6li40L85N9uTxtsLChNiMYwU0MIAvFFeLLzxTOLVheb
jKN6dtrjFlcj3zShC1nuCdrCPse5HkVKeaBYbEPALpcpSXAypxFug5Z3VpKZgFFwfBzMRLmlFodU
OBJvU6xwSjClboIWM0hDOxFTzwZY4eqO6PVKRDndzvfs7o6dIvRxqqjGyde9zA0i1dTYF/O02Eua
apg7AJoVLjVI8TDVd1JJk9XZSib/cRKmBYjRyzODyxE/DGvx26gSPVdPDmzvwsDhPF8WzzX+NB6Z
ikxFpi6kUce5dN87B/bV8CzLCBS5pPqRIeiC3jMV9VUcBfKifdKt9qPcXTev+vNBoeAjWrbpH0Bf
I+WD9/oFIi6VlgQoAb3i9qjHFtrGsOnAjYjLlJAcBumTrwz3/fXHR5tlAmB7rE3nwELnxEBL85o8
+jKNdmAzikbMTqjQL6zd8X4DgCNzIpjW10liO3bEM85vYSGuJgmWBGJFZZGf0bNxJyJa6NN9aiHl
pphq3ZS7NUr4s/gr/9aG7e1cvoPM/5kEI7LU1qRw/8OWOFxs+bjvHsbZFJs1MuAJlkmSE+j8mYgJ
Ndqug+226qK7/TMpm0Qe5K6/ZNjWpBC4M5zCArv1efXknf3Fo8ItsdDg1/CUY+Og0ojkA5dAUvjg
F71Yv8QPWn+cH2kKvluL7J+u7dNWj/cVlJ5iJP9EoMXjzs3e05dOxJCRkjBksyIygMBeWJ6JA85v
dVPxW1nwh1vvLdBuCjz0KkxQfS9sEDXIwxHN4EbMo/X1+rqo//ryV+S/IYY2fp6HNtplSn09pDdD
JIjI85mSaHFA9kkWZLE4qfQbtnK2lXPJCeaaDm33dhwlIgI7TWUr8npOYlss7xdguHDgHm2X4DTN
uZ8lAu+9EQsmQQ9/9RyjvL+7UCA1dytgNOYwfICzqwlMCNRx0XkPlQjEmA2HP+HyugLgdJoMHLhd
IRg5t/tyxTFzlrCzE6CjWWVIaMf2Edcy/3eQ/hw3Q2WicBBJVpETvivWHAe5dtiZdUipbhGELS/Z
KaiGBX9B4zOab8l8dWnV1vMD6DGsj3A+pklL/uWcJpBxtgvJkKoNZjlfiissDHj0FuK6PAu6VxNu
l7MU5dRzKQqQ/que+aVOQ6lyRvl3YROSlsABAq6F4+JQmXkrxOntQqe+9Pls6TbMwKVNXXowBRL1
Jspx72R+BxOUDoomEmGcl0MzFRdFjd2N/A8bW31gatT6rfGdXNLgKNwOjCpzfcUWnY1KkKJ0iL4+
FKFVffMpWM/6x20sQlOXt4QwJQtUkQ/jdW1gLZZ7rScXZ1FHtVfC8Ue6suRdZBcF6SS8qIiJ8ihA
MFcYNmFoGZLqkbx0wXfC1eD6BRi+DkGeHhXUjgmJqP5F1vk1IWhXF8jsZ7VIhn1XcADHaxLaYKzl
vdLQr97m/X5EbnapN5WniF7ZPt0GM1fWyz2669kHXKwgYrwKoi7dU6U+DFLfUKjWfCc+XL97Cgi3
n1o/aYcgYPEKVCTdVFoT3ndsaryOp4zzECgjJOAw4FemRF8JbXgwo0FuEnGCFsrm59anJNu+erGH
ANHm2SEgoU6vaUu3ax39KJicQwtP03a2DALUKaRIauGl1QS/dAcEYrvb2iCoqYzIxMspT/oJ/YGL
8uAciwZLkeo2MAMn6+9vUT/pvD0s3bUoH8gnKCp+XZPhC4k8YpxHoqUq9VD3NHIN0Nm46G4iFJ4T
3lM+t/iiGUeNiHRyxrOWvaAO4VV0CpkFVVE/+/rvrVAiFSQrxbBbioqxIoMagh+Hjmxh8i44oAja
N93R6e+iFHn/g9Babvkw2zSE0N+1Upc+Q4XWokAH8+KQNmfY95/4jw/lzl+yf9lD4dbdE1tF0Ivj
Dw8goJx/sPb9tkx9ZD4bvxy0k1FJ7fG8Ea73s1C1WJ01U97EMOIB4RnjPrHbt8E7ZMKJ7aI1aQRl
wnVpugqIHjbnkWfLVqPJWMdFHXEtp6SnMTeiRLSKNf2I7T/FrIh6kvGl4hT5BF8LUGmu+WuomiaM
SoZJLE3Q8Jo3zDE9BZGWosbg6WExZAW5Q64/5f/fhSImTF0VdwSvEKQkExMsX8GIF5hpdaeyVL6y
Ygt7V2ofmaVt4u6Al4668kv4hITWl1wKCgn49cAcDHo3x9l2qS1R3sXJK/EVi4Ol80w5KLERyeAS
DdpvN777DejsWzDGsFzM/H47AYMt6X3tEh9oZBV5EYRKcRptQmwr7MSndiirKbXFZIhOIz/Fv9de
2QBoEcPmJA4iJPQQL/g65682V8cH0UriD2tX/cEKuGjv5RtlwdhdnkTn4tTX8HOLjFeTuIZcYHlg
i5rovFud8q5+bppr5ybz5fqub6J0/GxujRfJikRNBviM64L5hChQRLmOREbCq/J3sArNxl9U29WJ
Zc7dEGEqiB5pxR9KgXhHRzZxHBs1kVRO0eNGJh/WBok/Ev/8/MaKpQmw1KadmMgp4NrCnUse8jvF
3IdDzk7KEg+WV3kLGeisxnCUL+TvOKWlfpHNP3XRW3iisKphO8ACGLgZGZnRyleYEdKpUPq1qQna
MSD/fw8HaWN4hLb7k6LVFOttJXdjxKGHY3BwoLgV/8yyDx4ZV9Rjod+Z84RPR24QRzeVNziT4d7G
XiLW/exuzEfCevundFAvP170axKHdXOuon7Zc4xCotpGPR+MSodBEiHGtZGaeQj0veHJewuW+8U6
Tf50pa4Mj+Pt6d30aDWg/Q1myEZs95ZAg7l/Cc3NBbSW0/l5gMbU2+tft6KSRNvYfk8bNO4zuRTP
RZdgs+PLm1AYLMlcpz8cb/dUYTwjwAZtIPoqlmn2hAiSF/GXK604Bh0/T2znQaVShRQPswDJH+lB
kM76lHVa+YQb8Q/E5CZOen3/xF7zQSJRbxPOChQ2lF1SVurE8D9Edtda8ngaVX7BWN5VUD0i1GN4
lAXj+Ml6gRBgkbEX+VWz4ILMmSl4ydzgME0kYYTQ0yoYK1cJcKI2+ZOxaYxQMY+xlQCGAsdnKSG0
bZk8U9K3flYKJk8kS4Lgp6KaqpoH6ySDjU6hwbTayzWB/QF0dYhTQvu1X4YKhmXiZeeTL1ynrNW4
qswkLBUssla9tbGuwu/c/EfzG2vqLoOSmarecPpmOPi0l/LTmU6bD0sbYnU44JPsbjJfb6u8Dv1h
GByFAycFaSm6wYD2fjWCZeliXPHP6QkVsUwtDsskAzVwNu4B8UfQfHkTieUps8N2r48IlsvedMSl
AVOhnwdL5rjhPa2PpR4wpuFRa2ryBXzHxyL172zK/l+GeDqdloDYJQm4qA8mpe0rBHOjn6xxeTID
LaGsPDRFAie6OOvXxXcf4N8hDOUuwG5SMqO5gaLgc3UaXH3yhdaQqRHv0AIgPcldVsrxB4IIKnwP
Cy833fG8IfMEG28gY9+xtFGFo4JA0h2OYf1Ga8zZc0XPlPpiJIjV1lWBUh1IoNBtwVxJzgLuMhXG
bKH/oHSCkAQ5wZR8MNYxkjPTuksPz08tQ+bROmykTqmlGFnQE2QQH/pwWvIIh3CTLd0zOTIR4Ou4
LUiqp6zNBw3jbSikRSw1ghDdicuh42DS4gL6Zo/bhKHIMQquxmQZvuNgauSoQYrAzk5O+NLVPKvj
vUMN4WhIScWmQTV2Mt30nfHHCjkT8zrsqtygHgg4LfEaVMeYMiFAou22DlNHx1TUZZlJyV2tDqlt
B8rCmQcbyhvnvuCW0dfThs5e3vwCCLDxuVtw1WmsX1qOUaEiM5Ia1VINAULe0N/18q1rhwbjMyvJ
J/2tJSLutbBY/QjslHOpbofUEyK0WskowkM5ZUYT0UTnhyNFkqL9q26/5UuBBFE75kuk3ncffGDZ
f6s3wodiqwCDnBtVp+Q9UuFp5lfgcMAsA010Ujm21QTmqQe48zdFGyQeL5L7BJDZD4o3q7gDHtj1
7CayiGJcfYrAUVaW14RP9IKG/3nJ+N1tG3WaJhuLm0suW55OJdb4JHavvRhNCmNGEEZ3kb8G7hnB
ZaWuq9pkhPQBTyA61xOl5I8V9zyc+t9ftMthWLbDng6FXFBvkSlYzwhB3TKdZZ+cqOekOw0gbmMV
mGW77ZCG7HXyBF167ZcwpepShwSQLomXGbKKLiDQ1O0VrIX3gebIP1Rz8aTH369QWoK4qJJcNwSE
PYImzc7K2W3Wndmn62bTvwwes2dHvpOioem6Yj0TgBu/462C6tmX08gSuP4t7RymPOLpcA2sMnIH
dMewfV6/I4JgwizmwXYK/H7WtfhnrfzbdFNuDOhXsjULVI0oC/ybO0mFLOGwvuZdimpKvrHRcw44
SpXYIfLNTsVXXvqV5NnMoY1gTBMxntK07BecuxMllMioHIKzQfZfHgHY6u6YUcRyLGUrb5wMY5Hc
2SKIzSP1WhmVX9WciUstO3ZkW/S2VxPfGl0njIv32ZzjeDfCbim9vvqVNuJMqfpkTx4/wV42WATD
XeGm4c00NS0c623LQuPg3dbPj1Z607dhHxXcAOYA96bd1VmiSBtC94kDssDtEnEclyHcqmVGdfNK
oatVo2WN09ZN4uILdmiRw4Bb7awE6fKvAOogKHdkGjkn79t2RLTR4knSTflZuZmga5DliVq5GNwx
qafd/5Fo4MsGYCT8WlsPijCenjO60QuO94sYe8fuHsMqt83MOqqXI+AKIem0U7mgOWIc+2FwvnuZ
c9ynQA4xg7wZ+VZu0dkv/mBvoK1NNLk/HfdfvSyQEtwr51UQoXJZA1QulKHMN13GNrfWpu358Q0+
jKx+T3kpmQLPBUw7DjII6wxLmgLFCs+4PWkJw67yAO/brYz0nPr2sWtzmYpD36PsuEDfVMIYfgQh
R6LAS+UxHcpQxlLNT6TsV8rlWAGwOc1OfjInyFzBFmBLutdPcOBlwRe26fGcZ1xLisUMzExg47OY
uYfrf3gCqbs/AUNIfBh4i+gFX7ERpYOPYr4FY/VqCYq9JoPKc2efmUWxezIpzVlPa3dWbudlt1UN
d8e7EDykVc1TtmCPmIolH7QcvuljxS3R2b4Ln583PeC5ifZy6q1Br1aTUCFQL4nxwn5ytzEUVG2y
lKPpZguSqVTk9XoZQa2RTVrbp1ooBsIgWZCBKn5JmYd3hUtTJQCXbyZ/IL0Z6PmdTvNJxH1kNi4l
GZcjTo/eVr1G6unGE+w2d6KY0geUFw/7/1MHxeh8TePQfgg2thfCGYxxNrTDYtBI3ShtWKr7oV0k
4ou2mqzvRz089iJ+uQp2eE4E3OEIxQJbUph+ZqwGyvh1zxiLp87qcr8YPInwxDw0nEVoCPFQarUq
HrzdwDkeLGm7SNtHzabrzq3mzxRfBcZh1QPssJ64OH+Myb6zbD8rPgkqK5oMAVC2aIV1OsMv5WdP
Jc0LZydRtfwmm7bfslYdf3rfYjkZuE6HwOQ3bsELR4lzIG6WHQU5EAii0j67PH/wYR5gMCKo45BE
b4RMVP/BCRH8Xfd/0WmYnRHmPxZSBa5LJxIrkA72FaLZ0/Rd+VlgaU8jaIv85yOE9SpNxIxhz1pM
RvcIYCjLBlqfMs7dDcmNXUN0U0F0DA5dA8r3Sq1IQ6YsYA7HNXAyVxmx+vYp6Hk+nK73OFTVYbbG
1p2rBWzg1YINcpCXQe/xPEdu2ZEBaecD/69kqn7yuTp9EwuLQEUTAO+gg+/hpMH3yH09UVTlnu+6
Xwwh58QpzFlBHH5jSq1HLrEy7KPSZuo7eydPNthU7BrNAWpHCMeSTa5A0kP5iEPVfwkpHNGozw5a
eGZ4FHcx23om2lOceIW0ycfeVveRQq1Ku7fW6cdk2MBzJof9fhN/mxJtgrGs3gNXGZXb9ctvD5uP
y0oaSqtxqLnpTGMNorAcWzeEZP6O1notzLpS+JBLv1te3mUsoosutCoaZXEq92/uV7KRi4aigBgf
oXpdhg6HpcPufKWUXE3c++WhWzE5fEeqHXliOvZ8uhc/TaSl6D/rr+Bmszkl8iANO2kjzuFH0Zd+
HJZfs+jL1huBzM2U7t1eXOxCgfvqolQYeFxkUTrXP+hucazqLVUJYUVjx45deoY2JhtE1DPfEc6Q
w2wjJgY39HVFNIw7moG0/P7mM0heLiYX7Yug4sd8vNQM82zkmGwGUd/tvVY+cncDZ2cH6aHKhenP
Pz1PgMpV0+91QQor17TAkMSg9E0iIxDw6F+6VE/CEq/3mbCAnhTm6YIjz62FFs5nndGZNu1r8Eci
WNjTvLg1VuSKxRYNV/Wc6/OYwO/YEubRLQjC0Ou7YbLq0dAcQ5Y2QVGVySUiVXeWH2+vd4G4UgWJ
3XX4/5eOuRMhzSom/gr4pwK4ALBNHQR/Te7vaFzSKNrKiC6kHSMp1prcmocVf0KvylJo9QrJel8z
4WS7uia+dvVvqA7SFU2QCkIQxwxkv3CQHHYmJYFs2CaN9+ABK5fIOw3MAuY4sDpD0r6m3nSf3DuP
Pk6BlFfnuKIl1Zuzpvyo4oqcoth2i8DMYtPEaLTHd3eRv8A/t4N5e6sRsK8vVQnePMn+aTtk3K6u
HTUQ+CRvd6EQ+F7kg68G1HXP0Wb4FWEGf/uoY0C93vYTPI6Yi9vQqDLcJfwyhlXoWg4rPm4RkL4+
N25DocJd0YaPt1n58CEB0d7LDJyNcolxj16CykQGGmn415K+Sa6i8mlCvC5c/dYd7j5lceWFPeSe
mfHoVZpN8zhyNIa5GzcJ9rYpocoTO7a7jF2vH5NK/qmZi4fUUwbxxV1nvjAsWwh8WQtLcYY3A0Oe
xWxUuxy9I7f9cAYQTOs5n3oG8Uy4hEmw7yr86rEQLVOi3F4CiNVyoDj+HXkPNs+aCMjNRLuVo4cY
50LyuiK/pjr/6Vz0/uwh5iM9MLyGO8uSxVLv/20OV5q58kAp7qx0hv3KKa44ZHEOL+rPBjStcaPj
fTcodJgn+XFWb1UoUdcJppl8iGdNiJ8zKJHjTs5sIa8AWPF6vwQAE0PW5byABHPuag+M5LhyIgl7
Nvn5R2uV8OI1ALKffTUDIA2dSfxe/3qkKnmFpO8D3xKlQipn58hqREtDpO2L1cMMDcosn+5RgCiL
fL8a5WjVKBa7ciE5WeMOsIFlRL2Lj5si98jhPYrZAdRhJy2++B6N2SvAERLVOxlfkcTFm5Ypmak/
uvJzvSe5RA1CM1l1Mh0TJwqLWRnJCi1LhIadVi8+4uUeMWQplxNjPmyWOddw7Pu9m3VWucO7Hm9c
bMS0mosXFjPAS5W31940AsMxT7HTLW8W8EfhyDUUuw2NTffAlAb3q8DbY9eTnNGHACbeIDyvcWTU
cywUqBZwPqgYVnK/VL85M9rsgHvx01vsWT9FocxaTdGeWVDvVbFkS1GO4pN/NE3zHilNLviSDFjY
XCutMdUG32hB9WoqTzoOq924Ed666bznd5H2bqgbJuLAfCAbG4TLfSbDPV6H1bxqWcqi/xD6TFBp
flqyUL8jjIl7e6GBII+KpDosOO0vvDC+/GVjgLHnu0JlkAKjM8QQYxKNZAW1jhojkBbGzIYUZZhq
QV2I/+5OoiNp28OeDbDqMI2/qISOfeRlfQNMhxVR5WF3wcbUR9jJwYoBUGYrD2lM780ZAtoIB/aw
mRu8Pe09YOQq2t3JqcYOoVX4rdW12t0XhPFR8gdkHM49dl9rgsQYfm1IEYAsaZUEQLxPFF7Ty9dN
1Pft62gWTy59zOhWlhHS8rXWxqiKI3bb2Okz1RMoe1zVr9oCJ21EE3xSsCCZwK/zIyvTgrB4xdh6
bV7jVvWl9JI/KkJmK960z9laZ6mVMYrCiNNhEiJZHulJ3XI+h62aN4Ruj/8Ol8OddvZH1Xht6vtl
zCNp0Q7jLmFMWhJxN8uyzpU7Vm1q4OCnj2PmssLVepzvq/kYPNuNaU3E1dflZ+QC0+HoSpHYK1x/
ZblAwqxdCj8sMdyEKnRokTvPjGSCh2fr6YcE4FTydrqltLNSUuB0qC99SdgdqdsLveEhDKYOuTBR
YoUhtd7qilVEo7LBcn0udTRzp9m2Egcy6vmle6/7QwMNrvpMNAPFEnuV7YXUSa4CHGtJakhD1UfB
abo1/z2QU94bBB8yx1Jfic3pTit28OsQiqq/CBVVjsSGuBETbBL1B43PIQYmSUIl3jUyxzJ4XwUc
0kGOqSWfcG7XjZDZSJs39pUzJrdH+6XNmEtxfm0jwaQazrKYZt5qQ1X3eMntaB4rPnSNgGGmxMCX
+Uo8gJNJnd/aUTdyBzzzY9Zij4ULJcDrB6Svm3BvSbrh4FUTx02tNyROSGWnv7+sDn/+KF4+w8+/
VgAYTq6azR5rj4KbzyDDnCNwD8/GHryiPpp3oIOgiSQFXFw2p3yzbp5wpLiBHKJ8tSp70MY2iiOk
uR5tSpQZw/9ZoulMjEQqefVPUOPm1VbY7WzVpFzGzIKeVOcaAiBTVtZBEKxRCKxPuLWBUpQkSD80
snLcla5zjjg169y0bn6pKf74yq/+NJJbCO+8aJZ9OMgYmbp6uHab8JwmCtbAxi+RKB/xVBVgVnlm
QKTxgaV7qQ8muTXtNcAgxon0tN52VIMNXM7ucZMgynDB6kNczoHOI8XdQFhqRC775Wq4Rm6dCIW8
xvHhE7NBIG6DFzxN+OgvLCq2oGOOleIjCEnQFdwNI7PxRe3WXIql5zDv72xjFoNf159EtuwZcz/P
wb6RF4AiqTDxAvl/wZvXWc5baV0gtcoJO4vOZIio3qJ9fkd7TtYZWCBXQfNXPQkVtSsbN++qtdjz
HmbEF8AQb+eB0AWkTv8a2UroeAmE3pJqApS/q/QyZjuS8sfzzT+1hCiO+JFaeaKuTqZPgnI4RLrq
GAq4/v+XwoIjQET0icH4eonxZtihZ6bXSjs2D0a2PcrYSgBJRXN5xVdUdOPVOzBnyrcU3Egb9YIA
MtwKY7jYZ2A412HyCm9E3Z0wr0E9OQpzTfduWG4I0JYVXw3QZNOOkCQrav5b0mJED8tcZ/RRs951
6PJ0Zt+RD03meox7jrIfKYEHHOENTC6gPui35OvvTCY8/hsa0xU4fgfTxzkLuORwGN5z2J2MfSJJ
NY01RTxhS8HBKxcuE/Mkdx+3U4jG7m4fPq5qW9TsO7TGFInuehp6pDHI1uO4/DC1iUJ4eEkLZV3u
ZDLIqj4q42njaF+DyFtYY8s4C2cVrJrAOomxFsd5lBk+jG2mZh3t/GKo/ScikReGD5rAuz+itVti
X0nZAVage1fv/xCUk9iXnMNIOeSpEQBtKu7mun8lDyCpx2+K5S04MjtLFaDljo+TqPtkIvFzMbJN
p0ZZRkh6YVBeSDOFqFmmfj01BOCuD9PPFwiReZqHNEr8eCsoxaQ2yuSAhnafEFn58H6y1IVOLOXG
I5wseNqYrjetL766INDRrk4xP3IY/YvpN9DXUDBGW5Wn+l92dGEj3EHSOxW8PpVC8eFOjA08TBXT
6hh9XiVSduEFVP/gnukd8ccRnf9SJXhd85gZfYsx8yPQ18P3AyaeNdMNHwXV5FL6oZIrRYoOgCGX
bUdBOVFipHHHvDxELE22h4iIqfVZF8cy/82G87pmzFt7NTscuW5iWRWKSstGMEtlSO0hCiwQwB+m
CSIPbi0+ViqsOLHGZAO/77ZTqfJqSrOivXh2bhe4J4k2dngCyJ3JGKo7+wMQGOyjRLCLrYT1IFLm
YNl1dIf8xKrQXAnIp8Nc3iXfjV3X88D/3ReOFaGIufGkMmejfD4MvYfhcxpAylfNKTIDZlxFRwKi
1ANcPGn1WRgm2Du9d1LBcn+j/keCKCEQikhOg/Ko2XSqo3PUa/ftk+p1eBRD0KDR7T74tV0QC9xu
N4FEff4ZZVvu7isunFv7tdfiWnj7JAE7Bx/bNajnkCSiTK5+PHsozm8aNjKmrOzIk8ZCjRUkQCNl
bX0S2dpFujTyM+DmZDjIATww6hFSBp+09USsmDJjHsGLhiHOzcZl/EziUcmKMvKToa3CytBMxxFq
ws4JnWuZpGTML0Cta1G1rY7R1//4otzQMcsuqtn9iOh2rC0GsnPSS0vePCVZ6hnOXHEqsr+/TUAM
SdvXIe/c5RTJiklD9kD7WtRcod3YAjE2YiNMs8Vvt8w9LsbfNTXHSYPqNAt/lK79moQOpm7YGZPH
KZxNCRbdTMwMi4P1ElNe6dkwhAqFPZ3/QnQIem/iRIydMXEk6lc5hcMEgjesdGHLUy7WMYJaox3X
5VDS462rZcigU/bIE4MBEFeJOVfiQMCRu5gzzYVTsICE3bnlEbJJrKT0FLt/k5/fPJZuvOWDJfDf
RUrYqPuyXhutYFfBoSni2z/dnUSeXcr2eFee4oT7YoZPTgW50RyUrJgBwApaqJg679wEzVumzyXP
/L4eeV43zLwWZRhdL0TUh+86woMKBCMh8idfop2YfMYFeWAFLMzNYXsJBcsLOzslIpPUE5zrzVF3
HlpwH/RHWKFImZjAto1UmwMB2tJS8GpMdDsIJf0UjSMX3+e1S6047Zjj1U9HWd+oIDGvAcAdx4xC
lyDolHBMYHY8bS48GxB8FpwE1bTD5dKnUw4bN85e1OWn9JzIkdfDST+b3Y8+NafDBNP3BpCqup/9
5VOxTo8Uyl3bJRnVTlRxjfrcye/d4xVhKWtElP9hjGZwrmExn0h9jSE8I4Y3hNfjV3m+BqONFQWs
USRZXVYuq4O7Awu6NYmlkZn25QyRogCqyOZLIjLwYBTCsjP9gCDKmFqiS7KlIXSoaK9KsiVrv5vH
9YfPP8o1qItaXpHRE66KbQOL+eX+OmEc/Kdge3d4ZHR3dvP23Fzb5wQQUx20bVx3Oz7saasDhfaV
VyfkWT9uzSomMiQKCoXeasPjV9I0XyW/vTaJwvRzKIVEsM/tYu5U2mQ5eu+zR6xGAFmMopvA8bxP
GpomsMkHH6ubOe/zbVxboojpXx7y0AQA3tocURdhfyUItxTYzvrZkdw9nGx2+9pVblyW39snHbEK
Vk2T8rzetOCGr05O0BWBj+gxeD66Kf5yJ3MLWhYrt+BH0hhVb6HL5zWXvVcqZKXVtEkJ1lCahR0q
ld9X95u4Hy1sOtwHbcxJMCOuer55UVlYt+RZAuS6Dcn03II/x4pwUUTwC4084RAuszhUo4chojDu
HGj5VtYPxqIGKg3gECnEYYpqGU9ltoaxEcHM3Sb2kQTFPJm+UD+G+egOHlnp0rvb1DZTufzHn9rc
AqvoHm+i1omPiOGA3yUVQftJ6Tvc7gA6VaYs/zcN24h/KVpz3CG63lEXK7NcpiLtPB+yMgrc7Vjp
J/vKoOASd3Iw+mzTCipwFFY9BLrcCS2IHaHjJ8zpr+5EGgYUoxhwHuymo10DsCj7kfO9Ks7TrpX/
8Vqlb5w13OnzWrpHl7SeWG+AYF29VKRFDOFw/zAiDwIbq1wZFtuE9i9W0C4sH0uHcvrDUMD/hssZ
JTn06otP7qtPTMw+TMjMcDsmI7nWGQkmM1aglQdtT9hbHHmFEEH8IEaZ/yawPFhPxl3Lqass2i+C
n9h98ULxw3nO7kjJc+oJZxluvYSXCQU/3j4TEXrdIDwUbhayOiQXyI1AOB/+2aRGOBfV8oOi+E7V
ewCgnSDYR4+Va0qzJLqUum6LJtUXYKyG9VJQAV3OjBKaPrH3eBAOg9IM3kUW3ips4JpVmQ3FzOIk
xski0qIB7EMKfgBWtm3DOSsOZisVceBGM7SrFxtd+QRDZBlq17+bgKow3LhjXRHIvVds1HrjHU9n
mpIOUqD6KWSaNqWlYez9pjMoi2VTvvzTHJ88uC98KdRavacRq5xfdcFfwLgaSJ08tc/wCtFSM34s
bMoXgr0aOTJw9AbJUcu3sBoHTx7A73FSgN4fb36RojZaUhuDCFbZGCkYoQ6OPOoZCpOHXVr1Pn1V
Dzj2VHbdJ/H2zXVP5sSX7GoiJgno71RBeGP8DLz6TaUo1WngXZZsMuTCp0itPQMLILuV4nNN+4xk
3wDG4NxAxAZW5Vwk13qDhzcr819BWDJAOFKkqO3QzzBXdiFu39GZcQ0maxAsxm+2Qlsq+ag6Yyxi
BOMebosAk5mb+lIRVH90vwp0CcOOxBmWz5qrbdysS+hW6tXdhGdZUuzOvoPWUDHh57k/MVv6tgXP
1thTrmGyMpOSVk8j5p8xqBleNgGI+PdDxqwjWKv+M+VlUYyLcgWlLL/JwcR06p9D4kMrPM93SQ+7
I7VtamRdZnExLefPamOP8OBkOSa/6QeojfSTI7XxL4uEQRlRAJUKPKHO1+UBV35Mg2977EQIeZK8
nP+Ym5Q3O1qVG/FSu9h2XSGYy7qxvopuyii4+NH2bMuL3DsPPrucZ7OL4z3ACOmf1vIi8RQ5TZQ5
7YFLlrTWRJAsn3Rv7bs23R6nyyz9Iefyoh9eVQSRAUMK/2HmFJIGkCROgaahQ2YCfNAXjpjU5fgO
hpZAtEdx57n2TST6vagVB5+CatBqVvCHK384DRJaXjcROtxw3JY4G7HZ1rG0NzKGVWpzYo0qS8uO
3mmKvJ7Jx5ck7upjm7RfhgubsDO8k0XzyQo1groUA7T+6ZIRIXdbFaYbNV9keRR0/ogPN0rvINXj
CsfDrtIPfYfBWFNNITNUwZvSBdF16lgYO+1CsumDCgc8mQVVP58iID9nxf3qfMpfAT8b2XC8Jovx
zevjn5fCAS/+GPl7wucwH0EFeA9eocetsr6EaBwT9pPOejHG3WDmnX6yXZ1gycraRpUH91+9G2Kn
oq59/78vM2VYUmSnLD7ej5RkoyWFmIEteOjZYmjEgpSLhpQIcRE3DzQO7d9hKNnoDiz9IK8LK3Jh
OHXHwHo5tCsMcJufScy2AkvWNS5KEk2Wk7LEByWCHFAtnyw2GVi9u+6S3nAWzjTzO+6VEdVv6dyH
YuuWimVj5n58icnIDvZp1xvHfoR6dQMLR9qkKNBHQLIb8U3t+CyRx1JzKeYVjHipFazoVKzG2k7u
mRkISl7x9Qp6kvyllVcFPGbWfSlGGNtKEKjOsCQFS4IsyWl4o74XkE5fAxOk1tyepbT7giNgu8/m
DzPBuG3Ps0P8EpgSWb8B48qLe4654emPe7mPFYsXAk7Fe36DqEV6WnVBvyhor5nV6ppps1Nje+dx
Vn3OjjmatzkRBwOfX28nBXuudnYrnVyFYvlhOzYTja+yyJ+VBYsRBQhcNy5IdZzreWh/61+IypOj
hr4GC/vU1THA2GxPqVYl9Mt18Qh8VE/v5+TkesD7HAjM+QVjS+DDt77X4SscuwuasOuWan/0uNJt
1atKBSJjtjs7n2SsvY6zTK04J/dS9fVmupdcTZmrn4PGOdnKck60VVw0Xd+ll03pa4ktZavPj3rb
/Nu225B0qCN9cj7d82GreU+U5+Av/YwAroMxQGr8xKi2/G4BPVUFqt9Dl6eTPjfjeRgwT3XD/e9V
aQsIoKqMLUIYxt5ovsmryV6bujQINAkAcU0GECB8Byzi3/Axp88RBa/ejAXE8nuY5j6UWGxxOPGZ
+xK1XaBvN5zB8WF4fzcqBtjhmNp68XVcVnAlT0012nrBvUG/U2ne1nNA/zLjsfE8QTvFo5E+bdQG
s+Yq0LNAvpSulrXjEwvjx3FTf0dWdehGg3W3NkVyHOUBVWpVSB0Pa1RNqGp+RFF5DEZdag5QS0x9
EDPntOoF6/E43wjgtQSJ9+wq12HQ6u3kHjE5QW9xSDoEMtZ7BHeVXe/B4DlDsYe7dyDtbF06LZyI
4O30nnwjafF0wIJVJQWlXAgd5iCz7jOpAgCQIijHjrbzgO68qaN7xOIVuufNfXdbFpvfpUbB4V+0
SdtQXoMAe+hXZ1lO4EO6auc+Znfg/LVNLFpa8fH4xkMiKYES6aNGxyPV1PkbnEVPXpfmInjFNsbY
zHzictHNKZvDpnljLCCooA4QonfsMpGodWyb8gZbJAd/oEW60BeClRm3cLJsVk62c3wJGqTmFnmD
rPsNEfPKsEbDb6IH8wK0SkR0kGtxeJ5P5zDjKtTaCM1lTQ3FMeHqLbx7KgeuGMOm9yC/zCeU+aGR
7ya9o0RMpbYuscZLPEfH95hWGEs5zmf9tgaxJuh0eNxQqaGMxUM0W62PxorinRmPxuDcz2jYCmVS
/BGvCCssVNpVs0a/q7KYctPOube1qq2YGk3BoLbPqcuO2voDfy9owfCwKyAMDUEoZLD/oBi193sX
kQCJPLTclYl5UYd3YKHkI3sCWny0R1EBFMUoEsrRLyjNkUsuBSmtmPktnYEafGb+QSVp06vdbhND
aPCphOP3AdUNFaQpTIm1cOXCeh22aQea0DOtvIbpJvnJDBk5uOXfkJq0TnEmx17oeAsvC0vhwWaT
lVQqKTlEqW7U7OmDnDUUm/uwF/oBT248e9qOE4VyuuhBOCZec+iqkb+Z3S3pzV1MJJHBMxHsSx49
wZq0gYFpMSsnZfRmBv93QsOzMrk2GCoTePRc6suxEM7jwiCw3uDURqUDJy4sh6tEWmb/L7TG8pR2
/FaGUDLmSogqnzfcaN7hb5FjcwRetrrdRV9rFKkn6IF7H60Xc75aevY5EBEbcecVTuGHXQxqmEzn
WEQF0Kz4VSrSPoyxYF0MpQ9+91S+U3gtGjBrWXDmnHuyDT2JeKHGxEm3nbKc58ZVvdfXKAQIRIzr
aqfCHMmokV9ObLJGoLTLbYeZZstBavy9FGb/EC/8mTHG1Cez5Ug8skwCd1WHPstNFHMRvqnWd23T
X8XLCzDsah6B9UF5dljmevuoj3/Xa5u4gN8eRVlWozD2pEfzCeTHn5ncWcNM0F2QLXFvrkW+nmnp
3cZyCgGp4tTOC3xhZX8EkcMOpzaAq2z/iBpBYIZJE+4wBaP+fCG/lq/tCHsmn5ZV2NhsGRgLDlQP
7VfQDTdPEobQrnvshkOPdSHCDuvFygHWybWOXPL2Pe71LKGr49ZtPYetSbAW80ZwtLuD9DonO4Rz
MGt7wGQRpVegkD5JHtYMlD3d4xvFKPN0PXxRzkpUB47a9gnFr6nrnoSh3V2CX5cBOFpQGZrtROGR
OFBW27iodpw3h9DwiJ8szuCwbQZ8/HeMGKW5gfIj2ur5XNefV/+mG0dbw014WF2MsgePLtMLrJOr
8jyAwMSUBTRR2bmLqHWKjerj54c3s3k2K+Ofqt73AqzW0fZ1/2izQwrQbGwt+yuHW6Mp1pw8ZzDD
zwHS4sqywMDgOy8Q6neyyS9emqdRdo+7GMDgCaoXXxRFqs+1ljc73B444j7YuTQ9kbS5Tew9uLVq
RyEvJUoJ6jpWnDeU9D5mdLKq97HJ+AVBwn7eHzYiTjykovl+MeusaF/jND2IpTBf5RLxcT2yHEiV
8WHqmupS2qY81Nxi6sPg8JQQN9iFeCKGn60iwNMiYhYb7uERTvduLOkGJq7JkPExihd2tmJWtrQE
GMmTdI+1N0aKV1MfG26LxdnMjRgeCQMZRUu/dJPHgLaprxj8PkWhI0uPEMr5GDwUBpzp07yc7v0b
f3v3yGm0PPwhsGkplUY3xiDuRBGMvSnzV0S2AhxKr1woiRQ0pdiK22yJ7WzECodDiK9+skbzE+3W
6921VxnLZAb8ZIuzHxIA7jGj4c425OjnYBKzAW3QIb7GsdQsVEQVmd5wpGAsPDMlVV+zAoMV2Lex
VTL1L2wKhy8ePdkjbD6vEVgZ2lFw1UisVCX6FxiIQfZAzUmC6ACFdw36kLzZ0PKTsH3zd42cZ8+d
pPSHm3o34+KUxp1Ckp34+SStY49yTBGG6U8i61rHu3bB4WVb6SfeB1E2UkGG1LL85OsULMKsi8SS
ZVI13X2JBJTWQAOLhrVfAXr6+HlKi1SUgfOiSVEZKcIhncoRRp3esEgyKndQWToamCIvQE0zAimr
ROp1+5npT+tW9Y1sHOye22mL3rpJRHwC9Fb2c0wfObcINVZyRwUR9pbbACFKYvwCSME6i7xU0DBn
91QorOyRWmM+u3l4A5xQ64jR6OKvNyFZL2DLhIubsHHFv6Yixp0IkY6Vga4ULc17i48l10oYOjoz
x7JR5+ftwtaG19f8gON0pZiSCf75TYl1VxE6HGCwuqPh2WFlbPwiQ5KILLZO60CMjtYaaCE76G0i
RL6/Cjk+Rds3t7AR0WjyHgOV8+Fxos0uvXNldUVq6zq/KCuYQOTUBeZfpC/u/kTPHIemP+1byvRY
yKyrgdG3Ma2qBLuzMsTdfE45hImnwKFed/8A3e2gioj3DH7pFX42EYrFAYvBEdkifyqmw8JGfLge
M4CE7zOiCERenaGAFAZE2ez+Hgg2s/UgEFLf8P/zI5SPEAsDLkbl3b90Org7Oj3qn+HVY6tM4G23
fb/hLnTWKWE4RdbmtAqllsmJtkQ2rRcNgu7eBlmd/b4IOR4V5DkVMBoFFsTRWQJVE3fkHVPE2C9G
SY5V8onqxFYXU89oYFlArVqreweSyUD5MHKs+P6YCVrBmjLE1bpSYD1+1UFdczHtY5n7Y6XRRhe4
GCYevMb1zLCRgEqTqComJFAv76PY2YtCIMOOlAXy5lgHYmeBKa0o+hzcnU/Wl/Z0h5IbAonni+Pq
KhkgbjtemflDHzJJqQVbheQb/qgDxZUrWk/mgKDAyyWOAlvNSNXAu2gRkfiMDal9Iv4uQUp70P5/
IkOn6bsuH56LlQDfIDITJCKKXUcWB1OHwBzM/YPkOO0iW2FLbzT2eMp4OQJ501wGsUxLUeHCSKpM
sFv4fse09lf1DgT5qcT9vhpGiQ3lstHfAkdy3dcAOCvZv6p0NUNlpm6MSqtFIJneZB97fZJqWxe2
95EIHijlBlJrxsqKLlxn0YFgYbP82rrpKweaFXWUUOvnT7351s+oeN2JPzUKhEMjEUF1XeHqf6oW
yb2AMU1BC091c4x+jcuojNqKtWNLEimW+T1Uvgzm/ULc7Q6LVPW8Oq0AUPv1l37e1WANaEwEB7mH
RvuERxoXnj9vTG9653O/S6w9XyZTfaFaOebQpmzRme15o3vcbi+i4QtobKoKV49+5ScL2RVcFjyN
Q9ucr9/meP0jGDvnvjOkzaBzS5+X8ErP2ZKLKIuh0gnvYga0Mc5Qckz1KqwTQljb36mkI5M+9kBu
0xKbkJ6paKSfagOUbfSN5ezIFo+Wq9mxUr0aWWIRJs5sya1KaFcxOTqRf01Z3QfTiBma6VjnYxYy
C1+RoNKu7JHmo/yDsvR7EURtsyEQ8tSjUw7haqeyWjq0W8mKgebe3F2r9CN5DM3LB/UHXQDeHgnq
SHOKY0XNnHlLpZVt0YODVbhg8ZFdnUHVWtwrhOI4VzwdCIadJkMBdfl0wXlDypz6jrmA2WYQqizV
IOSM/m2W2/Mh3sLLNn4VwcWivOIKrA/jM/w+QtFwL8ktc8muE7sKWHbMCMosB4U1hODFtOkcwztQ
TLOf7ZENXQR2XPLR8bHjTwpL4WxwA4ELffpNqUcy8O1Zwfl64U7gbp6MDLhXzmDZB5XYJCYs43Zz
rQlWzvaOk9J/OZ29abhk6f+wdUXrQWs1N4/oRFtLvqCC7Jzs2V+6GMqjQRA65dUYsaN8twVeEubX
gXYRKIFtnN+ddGKFxyPxs1SDgy4tYRgB5oEPr32hub/4zocgl+3eG9fGc+A8/wZxlGX0lI+yjQUr
mQDuFHt8f5IBQ25mVEcjyI+NjtxvZXeQW276z+LMXiKzaIa0wvaffor9Dh++Cu5+zPb2zgDO3UUH
HZNUH+TE2ENDNcoOKY3CBYskvev7rWe42xL7qZv3YrCvRgnlCqqBX1o8lyv7vSw08NQQnXionfls
D4jftO2ieokdLH5RSjYZRcBGBs+oxWpLJTRDdhfl6Eb5Br8P3F0MvYMGhzYsmLl+sCWQg+iOLdKD
1uRpbUHO1nXLBTF8iPE/CvZ0ZOBr5VtDoCaheaIAh881crn+cYPZXMs2Dh/5w5xwbjaTw1jpovA6
dIopWkZBU8wT073Apc5+afuphntkiM5k9hSKRLq2ASmi1rpGVfecXOqWY5w1J2JDZDJkpYXvaDUl
nBGNM/J2feimjKDYPRIyU6M6osbPhccX5egCF8E/W1DQTIy45NlRe6+lS+mKIF6BGo1yumkX9LDD
7VPOXx1PjVRgqCawlzciB2+1iOVKPtBAei1gzCTiP5HiHSL3r9uAPdIYcLBwwhuVvj52uqyDptDu
8M9U/WOGIIf5TJPQ46+33uO0PwLmSHjBENVtGD0LMwb2h4+SAslZYHNDSaBv20MgVvdukU3klQ3P
NQHerGqZwuS5ztbvkEBA4zavTzDMAQ2Vmd+e6TXei9ZgXnqDA1UTTRJRKJqNJ+tigV+yN1gT7hJx
kHKh3iP4wNq1cDXuhdC2FTBbxHGcbuQaP6ka/Vi0HKo4L6GTpCc8zZsrvHsZv298fLdlc0aQHmNm
4HChg4tZ5BZmHAv2vNhCpuXSxVNN2RiFYDIIiMYqakHgo1Eo8X9kKDJOg/hAS9ICdLU7fNsEawqw
un2tDJ+KbazTIIw1UxFFEXPMckLkSe0zmD0/0OhSWlkehquUYtGsn6+0poXk/G2D/H4SCOdVvWB9
3JrQd+Gdepaw7qsY9dAVyhzhT06hWS9gjY9V2QomNzoNBn5QTpl3+uQujXZZY6DZOc3oFKnYu8uf
MdWiFZKQ8hYtBi3GPyArIsVU7z4oWyPQl0GNLswZUcEB6KupqQifLWNToYjZWU8fcmFIgjVoOQn7
eFiYeTR5xlBM6Pn4fBYRA/nhLxsOCLHyE7zMxEgB/xDZdYthMS9xVGYX1ABX792pwJtEl3kUDRyD
7HjTiSQGcRHNTPIQuHhElAKrQ97Z8kht/NTucpQWHrYi280xRnoZf0TcUafyObME4rYcCU1kYYY4
Yt2yEd6Tf9L2UPo/lYeR9XLFxWwLF9Q16pw0mNl7HcTid+CXxxIVDLSSjSfWMYF/qdkZEf9nSeOr
Bg2Dma4R3PzEhWOtazE0jEynRaNJjPTAjtJRlLN9Vv21h0v9gWcBuU2ZxY75389XAIhaDvcawjCy
HD84pbeM3yCMAbUJp4aoHvjsGiaf3P+t9O92ljh+/wzHo9Qerv8iJme+tE1NjPgp0YGlW2rpqXSn
tVy+JDhc6BY/+rFg/k4hBA1uzg8hIRKqfd1NRvPVa5C0ndxVTPUxltxKz8Gqu9c49MGikTv3o6q/
51ERbupgt3beUNYlZY0ekAdNEOtpDHohZrvrh6s37OK2lGkhmcD+y1NM29TXCRdRnHtS4LV4dHMr
4RVDbQls5WaBapdzeSwU3qyeSmMJPNybQBNrg2sTrtWOE7RlKNp7rKhiP+cQUGmDWPrthGnGY1kk
ZSMqUUwiv01VUZtrT5XmWi9Ad0IhtOi0D5mHU+MfNryxdah2cbUdioRipNVOxL7rHAXXO67VvKfD
1YxBy0X1wn8k83Y1f3VnWCvKU0SAC8+lo2xYS5JBECcbuwTHNSwcDvvK7/IOGoTUdWsXbQY2SezP
F+b7ztrdi2qpZTaB5Y/OiLCPbdr8E249sjciKgg91/q3MWfIWGd75UJ8liRuWNobyy2vGgQTV/uW
duLWUEbo5i4ibIyP8Mli/m6Ze/ynRf9opNzkhk+CB+8NPY/qAn9aMOVUyXL8JvIFbsdcmphkz5sU
XnOvwarOWQkAm9GdpaT+SL62TqpaywDwbIrFPJ4XNYjSyJkZ3pTEAstBFwdtOQDk1H4csi5luCpG
i2BxTIOaAK8rNirxjF96WmmBIbrOjna5Fansi7qm7J0ER9bpRtY3o9ylzMW3q2IVw7rylzzL0DdR
Rop774svPaDbW2Rkhi5vDrdSPWhqqYNMijqHaTUhj/3gPBwyoTiL0+e5M0+rG6gIxaN9Euj9Ky5l
clq/glV66R/UzTguuxiaFCbN8s7F4ltJwILjNGDzETkpAMaqDNaF4kXjXyqeSm8Y1RKAFpBiEH9t
SNL6mB+hTOtr6ivSfyN3nAgdBTuf2sLvhQmwsM9/zT/Igji705Am2DzHhQNKN87pyEsAUWqX3B4m
7dW8vh3qJbiKmCYn9u2QYWl/EuEmpnxKoNrd+xI6cmcyfugxsrvBpW1Bsu4kS+iUGNY75Wr6oLwB
U3tXntTmD1SaCaERhW/qvWI50AnSGoQXOZg/S1/x36U0BVncBCq4U70pfuw56A5ethwJ7eXqyetq
vk+kMBRJc47vK5cgp4pEoc6C4Y5a4rZiBvDPBEheTlq3Si9NdrKOsr3u1n3wsYvIPO3BBdUj0A0q
etTbNJ4hz+E2CG37Sg4DhDGOPUsce2nZNsKIgl+NaAD89v8cwnZ7+6St4yc+luBsANogHlPK5Ugg
Pwq0JkEpQdXngBgRrPce/D376lASvGeUAi6phej7U726Bu6G53ee4dHAVX+1bh7Y74g4eCbxWdwy
wKcXxrIVrPBIA2nFAkBJxS7SwAzrBuaivkINGr2OaFOP5jYmniu3OIGPNuQO2PLAP6mY5SiQBi8k
Dk5muNGNQiXFVl0RqY74IH/pG+Iym0n02IlVolyuhnXZaTs/4UCWfDZHbwx3yFHskXTCe1mXPpjR
rmMAO88cst0teYgtaVIVtYC5/4Zbua4LeWzgiRkwwAMJxRWa1f4nKUlmc4/d5/xk01Fc9yKwO8tt
cFoUXQzZRmQVJZKlKjKXoM7HrTHf5N93BlPrWF8WGTgBmgfgkFIKIqzOM5BYjCtMpJjHZi1RxCHD
jCFPpR34MG9LBCyUSuMpU4sigSFFXdJOPqyKoO6zWAD7ZWir3naGHnYXODcA6unL5PGC7rZHE8Gt
xRyppgb8n/PGMDKDzJJTmuREumJ6R99OJCyq2EuCKAyxkYZHdg4cxD7UvaQPpby9tjVA+ng5SNWi
rXUWWrnig98VFmCRoWxJ4adzAgHxqLWHqOywbotIZCKqu3qmxUwOQajRdcyXiiEKNwUXfJqsj2ev
36Jw2BmXktNr1CglpTodnUpGW8anWCVVvkuUN8VSz3lD6fYHRfxOYsJgMEqjat765vYxOtyAREKW
OLabFoP/OE3fw8Ox9MR1wfczkEQEw+BTthiYLM1aAeBUVFSvzWTWbh2pQfqRn9H31SN+Ez9RWOrX
I/RhSQ7iMb9e1g3pbdFP/7OuTKiCWeuLGhbbaiMHqlBbOkoAgy1sp+7mDKic+Uo6xCGVSNgTU3DO
VGVEUNacp+8c+axnw0dTHWwEjcNk612feq9FfCm+CqXzp/Rup8IgqrT81Y3waII85Z1lDST0XG7v
3sw51fB673VF/EllYmUoDQnX/RA4LaPJaG1IBqB22Ef+BzmOaDV9mIOeoaX4W2RaXHsWC2R3qZQq
lWCl/GUMJx88VzcDkU8kwZHF6EIZwm4a/t6ee6roJbwxehRLy+o/h8nOk3m4h3hh7a9wnJYQjiM2
R4L3G+Pf1ts85kf7ughPUzkEm8bf+k0FUb5joXO/cre0QEj+r3j4mINsFtaMDPdFaZYs6A4MX8Hr
+JNGVKsEuM1I+JTEm2kU+1gkCQBcBicmf/kUdNQevOyXS1I0q5KLOQ5QDDOJB+hwb3u9WoUC/Af/
CY4sk5sawm8yc91ocqh3j0cWv57XrnFzk8RFodkjx+ywScj9QI7K/SW5sBi23V6TIEd6IOErs9Xi
wOpQY+0Q0YlXPjm/Emt79O2KwNwdyAx5k9WF09vyi6J/kQnw8fc0UG0ab7zMdDy8p6WD13f2Xna2
FndcuJutjBareiDvAmQYpgfuMUpJ8Fi8Z/FBbQ0BWRhTXlgoOf3OwdjcrEUHt/1xHY3nHIxlOEQr
XTjlrguuHkv1pp3mpUUq2igTvXVaQNtIZjj8zSM0npvClZvjq4RDeaqlzCaM8UuUzU72qn0ftrzy
L7j+mO6BT+y0QAts51yDovm5LX8jwNu5iD0pQY3D4lYV4U2baZ6ycWohrfQuVkaBcJ14BJI0HhN+
tVv3aHVsD/IYz8vScSfCjOgdMDvQ1J8Fd/37rk1laVdeY6wNsU8ffar+cQ5RSfCK5Pd/bxsfNz9T
2Vrdx3cERqOF079Sc3As9IorhPNiD/zitHs16RBgNaIB0Va7lYOsnIbj97kdrReLcrjzBSmEkJMF
bk0hDLTVAVS85AvFvsf8eM66aVVj0WgNDSiQ6JBS/krHpxAqbygJxA9O4jrFKBi3xgkdD9Fj7Iq7
Tr9MDtwgewRjSeEX1RmTc3PFfGh2abW79REj566Y7dDXENy3LTvWrs7AXcE8LTMbkmQ8ZlOiXcZF
W3sL69SEq+Mh5siZnWXxYnGp6aepLH3sMuM6NXPGtCcB6Zj1x5Jg61j/hSax0cRbJyrshB309mje
4nEszd9kIAZ309lrGs8p6o1k+7XBZkzRXQHuy1GMLWgJ+zRCHRMfjv3QUMGgKBo73zqyTdS4dLix
8dCp9qYAA2so+9SP4KJTOl3on6I1EGwr9kXpqOX/coabzVVkuHMB0QQkeDBDJlnUSO4h/Dzea53u
wYNVMXznwlSExKb+UsF/ywP3/hZRBnUTk2+QhVxvGC2DA7PZ+dv8p5/q+YrB2WsoRYRSsZWCgNzb
x8SO0JCHNgiKQ74cyZb9gyVE7Af3MDoGZ1iK7vAyunOCU6gghCtpFPpm2pTYpby8D9mgblzMMG3p
TvxDzPfjx3tpy+kF1tD1nLavt+xTV9T95c/ayjfQh8igB5s1XAn6GLOrinVjgj72WcrMQrdQf45P
Y4tTyLTbbPbmcjanKH7RB6kFCprSVKr2IaW5wpnDFOO8N9LiZhtkKYKF4KnHC2F4HtnhPEqqWJq6
DTr+30djIyyFwgwMMlHAEFq5fMqbOrYq+ri/HcgBddTpiNnS1jTwCxYG2bvzOEeVVyyz2BQNft8A
al8qSZHZXpfBsX+zW3H8J11+I+fbW4WGgk6nKeffAUd3qVTIfn/SB1VKKeLUDw91IkZQscQl+OqD
kM63Rn6NWGmtef562m47jxFsgDNTCKKg9A7s1yeZyRJr66lJNO2DARZ3p7JtI4crhsDxoxlGoqKY
8vgLbiLpJ6E4JVFgWLsLFAyINugDYS0yjH82jVtZmaAycj8twl+BNLWTiMBX/EJs88orBsUM10iZ
7PqYE1UTFl47QeKX3oLkR0YmJVzOjj/otQU5fVRwhYqfLqPv8AXCLRZvjujpr5NgWbEgNNiA2+2J
tqvYRv+ZrrV19/th4cqvvOw6wc1Y4wuX3AicYX9wOsaIadGJHNqGIJ2tiHMYSjeR+FA+17EvP06d
mUSOMGxP966GGtnvNPqZGaK5OWkwQ8hIZMFt9EoKLhZTv6OtA8U1M3jUoJtZU+KNByCbKmyd8MBo
y8bDAYOztxq2KC57gMDa9mM7z+vL9uTOex1GX8bZz1yg0FcuM2GzewZaADeg4Iba8N2+kT7FRp2i
n286e2xJtmH62ZMM/RdsqOZ4RY6f49mJutQYmpKw/wn3LmNNYE0Jl7W7/FMTVnTmip7VI/KEq9fd
7tBUY4yyjwbuR3npbJ01AzsfYwngH39wARtkuqPOzAwZ06OrC5FG94+AVrRg9ctcJLmFRgeH16Bi
q5/Tcfqx0my1K7kIIZACMEWY/RdiGrEh0IhA8YM5U+Cz2planL6ztGdI7N4zrCjMcIIFLhfMHTJQ
eaGgKI6MP443t1qjofDvWhqIiAHcpcf5azjACqdkxO/5K/CsbMPxQjQ31YDVdwC/LJ6awbNXYrFX
fm4re2buEApMTFu3MQsxHzWyfGHq2kvFyVDAf5MLCnbfxG5PB0TVM2rcQp5Ikz+qyCmv4x94Cypu
sNH2ChIBGCaishNSz7tFnFAPIkw0JG5khfuU73RnNGAf2DCmMcbe9at8znx4IDMgEPUMDHZaJBsv
8Lk8mhPn2yE3GfKLBk1c+gv5wIYT84Ajfg0TVjPFBDwmXKK8TN9rU33ClrERBgkKKIPmVA3Y05xO
Ju2WDmJamUV6MuBXVnaO3OaklI3bxFXiNS4YXpTBxUs9M0g53cGTxeR00hKN2US/FKJ/A3zAgPUv
8gBMu8IV145s5NOvWqJU8QqbA+5PDErd6SUsL/wlLe+NE/8sl0/ejPEeUQYYwpKtmaohExpHYv6T
9nXtEZSVAgkAVGXTwMq39C1mxcEa99haogtjTVG7nPkK1AvQGDXXfHBgF+xaKjpoXYEwV+pZSFDc
/qpThKUVYXb1xkOxBTxUiIjRuB7q5iz1GlVJrqqZrNPYkBz+nPd4G6SpSh+BTfsbHsmThXEFn0Ws
5JsGGzktnjEX727FMKvjc4NUT2I/nfD5is7Pp5S+T4tYT7+Bo3u9MFGC97s5lEbvh8e5+aDacJI3
eTuHwjw17I1UPOh9ZMEtz3qUM8zgMNFhcJVVc9IA16rfygzFrhrMiRuvt6CmDoVQBpuYimeQEj09
aatL3zgQuvi7vX67b7rPchjpvEmvOkDw4nTegJDJHh0mLRtuZadfA/FBAOPdBRtTc6+KlFqppf6P
ppHFBHLJZ2lPHxBQNXDbwOvGn63nOEmXFtuB2YhfLxdzquh7EVOADFOQ/NxZNObBFitUJrnC2Oen
+shMytLBldDqctkn+hkrhocecOmFzSFaVFMBe6CBvJYOpnhE1s+t43a2hORcjXHCCl4tRfgrpDJq
jmc/Aoz0EEGQel8Y+36zL5hnMWf582TKxdVCjtIWbX0LAd6V7f5ImfeF8foJONRrn88+0hC9ii7h
h7QMvRQOnm9WJKsA+d47mGatRAqyAW530L0+Dqn5c3Xp8QTxO5ZSBGXof96LiiY1udLTIv4pSEiz
ulRTHNyNc2NIHYO16YKbuQFUD2AMjNS3FEbzPM5vZheO9YmNeiyKGsuUGRtK0WZ0fyKHi4tpWqOV
yDUPuVx9UYrF5xTlRFO1ENMO6pTkpjc+DMLajYy/Mqy4rau2++8wSIldlA7ZfNoPac9YeE6K8tNn
TA55QiBbgnCm+IYN+cjj0iBLjH5r1GEciwtE3RB4SZR2ZdKyn+Ugnq6Hdl+R5Si/TvaWOWa/jhSe
wtKYi9e7IPfcKVCR/fkUXLdpgeiKGRtuF6whUvBIEjeMQURm1kNoec5wkqc+E0C3W/onMDeS1K/O
Ir8x7E4HGhUJfMwNYDwi16qDjdgEvz+kEuBon5F/QXq4D9id0Cd4EfPvTy/kiatMppcIs5vTM26h
4VPENRkc2wPp5s8JhIyXdK9J3hH3ako5Zf0vFgIXvLJsNotEHWYnpVWYgTQbNIZVmtrPfVc4eWId
aRGPBnNEIXPkQRvIfNNAA5vRzUZ4wosF3Rm33s98sDf4esSSlwqC/ofpAd33WL6x4imTS0ckZ8cG
RZrQgUt30/ZlbU2Tm6fnmqUxGMP4/yA1L6Chjfy6gaSCB76P2qr8VZy3q8hVMdjZA6Q3ty+RVxSt
UlZEwjqXhXWqvNfGiae2u6hACERpumfMvNxLPrbrhLHqmaevfv59NEX6aat8YFyFvh5dGIflaXvR
f9FUUpBrV7Sc93kaYjOkRtvWGAbIiodvz2p216Ii49L/qM42L76bUwl44l6mfvc//dA7hayhgi6G
D9KYip2PB+539rC30UkrrKYQhPWte9ViAZnIAp0/vZ99DwwTyxEAO32ugAM+EH5nYDgSxyrLiVn0
0JBqK1X+aeMNz1iTSEvVcvOceOjFwrjyI9GXu9gb5x8vPAXlK5EuZf5ZKeRkvmiIH8xubHNO1rL2
RXjgwAwsqvA440neifBQeiE4hB9TmFzh5+8gggXZo9lsby/66Ly8PwLBQWow3bvV3osnO2MBvfFN
oz9heMc/yW30SxWMkA5O0VME3qQiXTVLNcOgUIXBTIpq2Xj3fIquN2i9RBClB3uznQ287XcVXYbc
s2yVQZCjyiPMBbhpJmpo2D/+M1wY9ksMgtqOlL/xqF0o9KT2HAGCz7GpA6m5CrwOSLyVAidgHE8u
2CvNbQUR9cQqApcDzGzQ3gURC/DAwgMts06hLkA/6FJJE6lStpiJwff6ysFN5ACoVQcVMREh3J/J
sqtZUaJ3yhlyht/nxfmy1Em9MLPDVCBZJY7n7dfhIhp5TifwfFG7nDFOCbGENrvsOUu1PSpng7aC
UrqnPXdm/ug1T54Mgdzh9NL63ADP8NHWwLlt0ZRwL60d2Z6LKvFEhIESWsMI7gCSccJHnNp8K+IF
XB6E3xu7cGHiQaFwezGaSGtYug3SVAPc3W7z6JaZGEag2ECwPEe7eYjN0L99L8zgQme1U1i93PYD
F0q/krxUO2cyr+Y/OY55zLX3P7VPYrWK0TLUEo2LCEdzNNLKOiwZI7CM/kBE4nJWOzOQqVgvEREm
9gRzLTlaQZJRblrbgnOL+zgwK5qDifu3aT6bmeazLAz6JDbrsyg2uvMMgtxsJL2zdJo/G7CrWGNr
A/JyyAXGhRS+NvsOPtj4+ioz8ar2bjUd25ZaSM7okGbGnz20o/ikHwqsZuZ+weXUs3IsfakBWvPO
0kpuJy2RB5UwkDxPEJVDr+tt6CWyDrvkjz9WdUcXeseSWL4zIgrTTXyAAEL6oc48M8kwDwfmYOSI
hS38JjlcciGMyh/IkQF4KycQT0XhrAQUDSBZYOEiXzLuvexoTlo3M3w3t+V4/qbhIvJWhyVjnX3P
Tz7PCXqqKujwkH+yHS52rEbykx06KtXoNr/z5FDXxoHEK4y45MSaGzXp3tCDvEKDhAnu6XbKSMmz
Sb2TfnFbfylFovWT7NYNznUpGq2IuPrVb9jHKI37DDaPabUvHt40Iinp1vsWml4ORbvpzkTve1Qk
B6ngc5AW6sOQiYRP52PohISZ+rO6PzkTE1Blg8fN8rpo1fZoVCbEpGMYUu/kTG+yavfORbjGjsdu
TnNCG/yRX5aNsMMPs2X+qbfKpFOZaU7D3HS9PvkHukJMz2y749w1/ajX7RsjGmRGuuKo/SaYCl1Y
tRNxZN6U7ONpX0UzzLqJ0c5P7iLXlN/PVeCBDMv+O8PjVHKxCkvy3wZCFseDnI73OO8u8GH3NGdQ
IG+b1qbiogmGDKkP52pesxtlN9z8RVP87X6dyQO1/2yciEB73XblHXD7LdrdVVj4EVRvVF1355IQ
8ebYOm1BxqEALtDUB02rBGNg78oN6yVUftAQ0/juZxEw/CGQa28Ud4X6QFYa8D10xea0MrhJKZ+V
DJY5gjcwUHx/3w0V/zyF9waZoftChxK/N5JVCM0EwLVB93KnmdqFB7BK8CGZbt/QckHoBg5Pxbfg
9aH6Hq41mxSt0mDu6HYSv0BqgYbWqEAN4oURm1sXEdJ7f+kOMgmbV7Yrce7BZPbchfTKvaRqet5X
Yr1wiGbRNJci1kL6whtsdhoxKiXqS2jHc9oF+wo6OU7elS2EIFExT21gLlmLMyAF5qF6LH4uSbdV
hMUHSI+tc6GRRIubOgNY4uZfL8ffzPaILou2Gz5eMj19hWEaBAa0BkLu52/qykI3JQCKObDLXyv8
I/oLZ2yaEMoyFZWoQ6OHv7KGMfgKj5brwkVDTRxK28GswA6k+68BmyUwx6VLQSK/lLorJWFMp2yP
VrhCrKMQWuypQRN3/ae1TiVsfR7z8hK69rEt82SgZ4Gg7+/bDA0UcNAHSmS9kQvwvrjceVWwsgsq
3WmEDtSs5V2Qj9PJGUVChBdeG5JAravR/dhzB0OPfbAkv9E8F6gAxQdINDb9zC/3ovC7HDIDRoEt
8wvU8hAzdZs4Id6cGQGb2qi2lTHzZRakpCCGUAyedSFGQIXZiZS04y5ErIxpc9Pb7sEBcRgleyhn
9EiXfyEvJKuLuUd6aLmREIZPJKBeQaCrYDvhNMGUGbjPTv0Bydol/uYuF6HMTdEVyj8mHKpA9GN6
rc6dlN+WXRNtZc0LhcIgwkQopIWykBNuDismAPh5Z9f1Ao33un+KX/WTSq3AXVx9/82YHBtnq8yB
YkFx3C1GZ8fU962ljeF6wOfGekWkwh1ZT0kbv46/Lnhwv3DY7CmJ+czDg0O14s6rMEnVkjSsF40w
vT7LJ32u0l7nOcns2m3hsjtMTR6igMrLGTxKsLP/LoTqdHQmpH5HK56IaXN1qek1WLmRij1QZdig
HKcm72uTjRvkXLkdYm7WFvJXpnMVUIq6goO71qNkslX8+XZwqxomDuG79Ty0Mb6Gwcvw/RiFSk73
7m5ZWd1kXbknTqsJLe1rKT0snk1naosxfwUt8Q9JmO07obyazhJsDoYW+2wxaYQrcWGvFCvcck0p
Pv2wIqlt16kY2019ip0hJQQ5dT3/Q+iQgtblPcWVu4LSaHFqjAN0/SsMIvkW48RI6yFE94PdF2G9
30CAVk76x+VWopB6QDk8nFilSy3kYUG4QvkTc/4IesZVR2hriyZYMcNTw8cW5X9sM+fc3EDDZnRX
1m1yh9FFVzJH7N4rQkUtjx3D0l9QbX+VO2WWa//cYdFOhAfEAxNL02Ib+NgmYHHgrZ1/y3YQ2SFf
3a9VnvpsjYo/9ttnKYRDPtsaEr5eBKS5Uvsk/dP0C82beBbbu+x7l+NNkBi8TSIVLEdVADE6tCOa
vETbbcxDBRwmWbJ09APZqH3sK9AGbra4FGil72b562XvOlw6kK/0dUphpVFOjxKNBik9mylHS3sI
S5RogNYhLfStMvLDxav7gK+Qt06Hf8fnK6uGIZjvuv99IHO1iMLp3UUpv5Ic1bE7yGzPqQTT6vXx
QFq7+oKXm7FDXjfQjj90M6BsZiaQIo363j71VKifPnOZg/FJXZ4HxwJSUUnxZkft8urnhtUcpiyq
/8rxgR9Ln81vtDAUaW3Yn2c3HiyLlT9t0oiN0ljVfBrCdaoH1hv8RIgD4TVTLk79umO4YwXtsRis
YzqnMGiWIe7KlhcZ793U1j7LA+y83hrGSvk9Sw1MkE1iGuZ7DSH2Y9tf7CiPffJftsLoTKQVtjvr
Jl9TyuIeyLdUcmVlzQ6UjVxJgIF6gU8Oa98EgmlmUjedpseIlzJzw4WA5SLGdQvT4zeetf8LIfBW
TR1KO/o2IJeIdPzKNknfYJT8bS43fvQTX6teFJhAAemDJPVHe8M0X3zBp8rQWrnN68wujhpQFtBo
w5CPrZ/iwyIx0t6P2LIyJ9L12owipPBfHFnicXvYKD9dvQU1cCP2FwjCDPDkzLGfpNe4m7PlsS07
Kn+jdmKw27PRn2vP1xxxSDQdx6xDs/9a3fCDY8EbdqaVn+vCObWFVl8kQXtQf8+6n5wWDWn9Uicy
AjDZXAQ5+zwWV6EGq49+890GNeeMhPmlsBcwHugbWibATQfnSN5VElqcpfrMm/SwIel2VQBXlDM2
F/voFK2JiT0E40WAPS39n6F5lxzNVsCb3RSQB442Be61R50P2Lq+FQMoQylPkt8AurUXfN8yfGRX
zUp7tcNUWifeaWuiSIePlHvujkgB5vBYnWEY0nRVC7LY8l/5LQmUQP5Xfjz9QOdrdNy67n1sUTH8
Vl06m+ZlUraCgraNudzhITcK2r4pw4U9yzcPsV/CBs7xiK9X+1CEvhhG22EH/hpcG9/yOUbORbwy
mlUgt+Q4WhaG16OtAZ7X7uCWnzwPglooZuOSRAjy1ZSgmX6lmkCOjmzWDzexh7WzsWgMWOb2c5UQ
mpPUnc6jetCyAdtJ7NeXLqRuEaUh13CxX6a8TPgARLPrLBuY+UnFOTp24icysFw2aO5g6wbsUNgt
Ymv+IqY+4QCuhR5axOUSe+NEVWbjdtLU9XeEaXpvcJJTWjeZHsryCdtvTmvxy6RATWWZK66X3eAw
c3bd19rg9rmSpwZRa47fYoEno0m76F+1H8C2npON7kzSp4ic5FCxuGs03Y5o35yvLOrsCrWH8l9l
ffJl2wv1bhZHsV5YGLK7MK+JIslbRfphfFZZ+ZBAOF2IQZX1zp9sUSr1mwV7nstPy4ipPvtZSSwh
dlg5+qLuXZ5cCcs1HlOouhINdLOh1CGWMizJfdFwWtRLt1XFKJJAS1G6WsL2JbcBOIcyI33U+A8c
Xukb8Ma84WkNgf8OwuDvaOij7TFIDJWxFi0Y4AoYXgJsiq6CnDw4VRiFXNMIS2W5sxZ9dJrVIhGs
JALJ1jWjxScUCZHgp+ScYZ77/eUyGBq9iBlUIepWPFz7sVWfqInCsFDuyLf56t805ZYXLQoZvhfz
jyIWYbNA8427YvYTTZnES+/Ct+n5x1ktMi6EdtGHHnmVkmX+9lV6C/MRVdsf/Rj+ng7/fZ1yHEUr
ysiAN6xjJhN0NYtJPoF0wjXZvBAdehYMh4UpTL2JoReVqtV2NlpTP8wuMNpaBfLTcojII9R/eNfC
YF3RtPuSbJotufnrxgT8NYudEna+nJCdYIxK0ahH1w9lEFeet/uoQv8Wx7Plz/upNddYIKfNifAq
Xbh4m/t+4WeCybgiTrB6DdgxDcyQnNiZqKDWCN73emPfwH0Pp0swP9fG1h784MYVhe3fbSEdNKJ3
Jwug3l5hOvSgo5EJFyWGk1rc3dVPiVr0VYJHVIQuyGvNbZjXAbrAYhiWYNm1WN7HhQC8O6+VJWL/
gQRgzeVQ7I3kLDoDZbqKmZbK60x/svfLspIZpjaPWaIgXlNeCv25mjsKbjkut1k3tVKUscd+MiHh
GjVgWRM+FpSww5zl6MasEBVuGxhmmBGw0w9s/40FwblBsSDuT7VlctIYl2MfxWB8wR/JlbrFqqkj
boPjWmPPtTFL9rWIdLv1jeWAisRlSiov5BpcWYOyzrX+Ka0ZV0150lUEvxGc42mQv09MbDXDamT9
8bnH4DM4OyQZP030jEAy/8nlOvtzOepaMCnwd1pl/Zr9jccHsCUG4WuC2dLhYJ3tZHbESFmJzq9U
K1THGeU9mb21b8swBjDTIiQTv1lxveevLveZnaUkRQCXkCDzM37VneBfRx3Kd3zngulfU/SUFB22
ZksX0A1VHPmu0M1E7Z0Zsye5myaDu9XuztRgLeJBYOC8f31QeSWkzpHXx/L7iI5B072+v1WBLFyc
rqCBleM93x9Mzz6ozmRl++kQDK2UVcWxeOBVpJI3CIMKanOE27PaY4khUl77AvpDurlqiCoNg+SV
AJxczzghN50krQ/dZllG3vElgHLc6PZk2bh5cppggGiFfWw+Z7P75aPzelmym+ahZ1fx11XgyeSf
v6ghPMLQyGsUj08QOVeGMOD+Y6vtbOvguN9QtGq0gJIthhf7rmmTvIMUnGXm1McHtjixOJKn7Q2h
tra/ey4DWnTTmOiRfndxcBT5Y4pAR5/9bcFqeP9nOeQIB5qRuBdM7j/MEnKtGLIf+Bi0lXI1F/18
17DtHZvP4RU3GI/sRpDilUvaC4pR7Xa8yJR0iba+T6nMRoIICV2Wr302qKjnzeH7NCP7+pQoQ3pM
NlT2PArkOfFJI6lnMZCp2l+V79eoaQz1KsDzUQ9V13AYVWsqsEryrdlVAkmB8O6xlIjr+4IGmI9q
H0rITC2XEDTZXb3srlOzL15hz5mfUOXgkvUeFtsPj0/U7qfIvzLNfSd+SJ6ezmcayD5LqBPKEfGY
Zq921/x6zABh95cckgLGAXLvxiesObDwWjxNWKH4JugSEjVS9QrVZ0eN0V6VUCAcFwMETCgw+BS3
vaPdtOFCGK1X9Fx2YyniMPfZWmdHPHe2UqcJdCEVlKtuWw2BOr41+OUTKQi4Dz44+U1c0gXZ012R
gZug8nm1DW11wRlyH40/TDc6kS9r7yl39jQNAtZHUf9lBY2HzR5Nn1Juhq7NL53lW/MwN2KB9jJK
hnoLW8XKQD5dBLJRsfEjhf2h3VthqIOPiWs+UlTIti8nbYknkkQ9pKBPN6s34C5kxov+EelBN3Jj
9q4Gprj5o/Cg/HtxdmfnXx9ses3zaSF/TNI//OTpHurYhMfRm/+Q6BZhI+i8swez7OYfto5rVNTU
KzqObe2P5sC/+kRGM+VpjfA2i1B6u9vpeLltRgAe0UZ/+MPtbGUpPtWDgyGcNjR7ZUfUbUxGQwtr
oW+B5qCq0Vz+/fpdUgvntz+qYWOe8R4D6X6JwHvxnR316piWpsvoozdJQKvj3aUTxr7pVVajICfC
hDJ2a1BIDWErm/g7wXpvmHNxXO9y2yjuYZw7UyVZFZXWdDhakBbYxetyihEGjiT6FoeQzrKje5BU
ngxHTrSHLnd9ZLcYKeGndgO41udeUaRPQvsKjV7mQV/9AemfvDZ0OlCaSbBBPOwZqKRc8yUdZOcy
ztUMeNMHDj0HY4FKaUsaKtv2JyjFNmTiUELLqY+rIG0TwmhjV+FfThi4mEHawPrdwKTRuYizv8Mn
p7JIcIf42IvmiGf/mIKc6ORf99W+5QO8xc6e/GEGPwNpP7lZKqghlDOAAmZZIfV3fhiE/nC/hHIH
XCXvFls9mwlSvnxogzyIXs3tVOECXn2ZAJXSQw9aAMDk4zkKZXwKklaC9ZyVZmrPA4juBto4iqpQ
LLJ/OtHhlvohrPPt20XBagt5WsRwDRaZ1+/sOtk5XCnW7JZcwexs5rv0cVWoqfVkq2c7ywjLHttw
LSTVs7KfGcE6yW3QpZujbhYSW+PTfp2X++egnQYi38GxPX1ax2Xw+6Jn+Ibls+yTb6hEr5M4ZJsU
Sie2D+tW3i/GXL06nQbdQe/NqMZslxEffhz8aKKHed3FkNrWh0q9eJ3GElXqFV4DL8Nt6Y1KE/8j
j55teTn/gza7vy5A3QWhfwUjU/Q/F2F2j6FvjY5rFRO4TMEJZkb2fU5bXwcGFdLUbVP5Du+FdinZ
nFvgSzd7zmQ4bTj80dghhrQtFfkAa5y5ZnTbYGxxiCUhgnSfcXtr27pxYq04k+KJ6UWw1fIwaj6g
ak4DnuexASfAH8Hc1ghW7hpj+B7ATlZhObKhQ/W8QElY+t1gSV5PAodtIr3hC3FJQzEZu+HQR3X9
L32eMH9vPpxGyvhs6bXkuBDdIvdXt45jwfIf/M/Vw3cjl8/Tu5xYydjEV+LRHg089GlnAudVx4x/
rn6pZMNK8Hc7iGY1nCh7UYAzy893bZwYw0sngPTsy/Db3pWUNm3NkWBn40vbsYtTlq4dHgzOB+pQ
4SGCZ6rdG5CAcd9Lp4SWiXO5sEo/cR1hdkjNOr2aWkzdxisDATA+o5K5ZjkWtHELiFfPg9ssM8Yj
q6D6aajFY4GOWbG583Orh3AVKle40moeqd/J9UyEhSau23Dh8PobxxLpn0BNf85rBkTGfl9zhiCV
DmHUgwbw/5YbMv/CE+Ay4MAIJ/AHJrjWXyZWpSnfswjKb2mIMqbhqQh94VpwGj3klgpfZ5Cz/i1l
KJubiDykDcMZ9GuuqQ4mMm4EcxcJeKJMVjXKmC8fncLQ+fIMITQYSLxojdG5UQ2dzHAoTVz6FIG6
NjOmULxF5J2f2731FxRSxexn3mp25UI62fNYJBnUoR9pOImW+6x51aTBJvo8hl8+y/zWyrVN2M6L
LuBr89sWOGaoEfobZxrt77mDJ6RyrMVyXhxE/IbMpUMPKXvp4dUV0GCaKTAoRFVmeh3rUnNF3UkB
3Kx7rYdIxqrcO5y0F12/eh6T4b1c/VcIrUf0osvuodjIXpx14Pi+524vZKmDF/meuEmHhUUxNdGE
yweXYpAVT29AA6/2kTINNIcbGEhIAvGplFCFzeHNdhfIx0LvjUwe/A/EXs7hxfuQLFjApr0uV0tN
6FX15AvNnbFJjdbPjqdPtMt6bratNG5HKrMRipzYIicVkp6sYf2RSF/gniZ0FCNKp6O/wk3bMJR3
+/WZC4ny7v9AqwmGpVNzS+gnB88ibVRP4xmT7pMCcSt2+E5ClSD0TcpbL3EVfffp9tBtCbYEHp8/
x9gvTwqmqkNC6/5z35GXxSYT7m7rPwI32eASbfwIyj+4CwTVyAs520EAdXym1Qo8XhujyGF92Bfu
PF1V6DMMqJrHclZUGqwEGn5i+juSYUBsIvLYgYpBEbHS5DW2JnYPOS6ApMTCACqDX7HZUW1/o5Yd
kjOTq0VkelxV2tnjTYAqWghAV/DRhtwkeNFmbTbk1FcFqeGP7JGaO6vSpybF9AcRQfuw8EQzL6Oc
a7I0FeIgHWMMawy/HKBiXjuGWf/x+TpVGbcU1rsXAVUK8tqEFltkQDryqxrV+k/bCB6x6CbSNaFi
C4B+TW9/E3dGqgrhHxzhOan0pL39UdruETm2tvF25uIYnog4h4hecxK2D1300E5jsIjJD3FAAhZV
5kR22JxE2vJoia4xASm3ObpHCqg3H6ibRBHejds6n1pGniz1a2jFowHOrfMo1k81NEo1rfMVSMFQ
O0Ra9rlksRUN1Udi8POXR4k5gh8548uc7GEHCRNR63NIZUkPJE11cc0vMK9C+59yH6aYj0ozqwm2
ozSaE55Dp72vfXg3XX8zblzf4z/tjR2douU5tsELgCsOTwhzx6Lun8jS+vWQD06PyJXcsyGX/c0l
MHFTRtiV66fLuT6xRUzQ9rCMiJmlAL2SDx6QIzpJ0Mj1GYUgQ04HDEMzz/xrwfeJD8W3GQTuWpHH
F3cORVMl/x+EA83QqX4r9eR4ehBGwdvCedVcPUgnK5lnQ7qHOR7VQW4nQyDKPHPUOFnVhxjv3e+C
A6RMxR3GZr/YFjRGXz5HBDV0YyWfrVL8B6eTHMKKslsPFBhY0skmbWBU5dXLUhfa2ybyq6jK3o4O
6spwkxVeFkX4pCHIGTSFLif0/m2k21vY9ckPawku+LC5j26son5OG3f6rBULHsIR+2zx9/T0Nfhu
Ye/UO5vaDrh+d77AV1Hvbxuidjp1NsuZYSxWlwn0eNzOKpI6zDzl/aHhafgzVJrDhcOJNPZjKHBt
1/JtClUEcIsbUtxBzVY7VdTsGht97yR1eP8KZ6REhpoRJv3y1BFzP8N6gkid4LmmFp3QkjGpUt/j
VnA6T2wlAlchI86dQHttnMTTg6rthDp2rEGmiSfSOeKizelGhzZgC7A7Q2M0vajm5So9zuetF9R5
FRrgfeYSWUsdr+hzFPKB3T5vr9RNlyd60ztddio7l7TvGdCCqtjaLkOxiRXeu9HYc7ztYLPSywbC
exr4vVSnoYnBk+bEm1MT2NNQqvzpwKJO7gzHcIVW3zzb9nWXfZSlLne8iDrNU6GNNxvQFS+83OJ0
UPNJaC9IlsjUrrtN+aRU91t4JhjcJ7Lsk4mBFk72I2hLt7gtyKHO51LsuGgVIzLDtZpacXSbfMZF
OhugIuRMz93BiPCgy0OpBcB4MKR8CwFVELmGSJngZOCmHr1LQmemYtbO+v57E5lNSeJIlzQKJAqd
S/A3gdjM2uUYMK7pw2eoMixX9x60KTnAaKWzCGeWOmRWPbOIwPmvoATsEE5xrOIKJEVyLKk7jDNQ
eQWi7s09IECqbRM9fTD5z+WetFUHKhZiQvPugOuS7rp09FLbmxLSyDHghGyJg38cxKTlHCNqop5C
daWai5ClGFwckOTaPH4QFljDy6REpQMbDGU39vX0bc5XSiTZcoq/r62G4Uf3tEBN3mcxe/VemKEv
YO0aALEkKV595/Xu9LEO97sUVT8i4how9hOak+isAqe5wewA7P3JuozHpsRwbpLQcBKLmIiMu19b
S8gTM4ElXAnO0qX3qOT0SDIUVItN4PKheQAXGlx+mc/TZVqRQJNnNoIAtbmkkMTaKCYBxcdH2bVj
obkKpfqfz9uU8Y/3fkNlYeeJND7QisCcW031l8/4MXjZnY91BndnK2mzLlMqWLVkfJTcqetCL3/R
ewtzdJKF7jDlcTgXwFwHjYDvAWR1HyIj02mIxSTsmWCr2Nrh3SNoGefagR5X40so4CDUpWUsN3TV
opC9OXmQ0vYlRYeOGA4pBsFOPsP9C1cjn7AD9VyAN9TJAKiOFBCZA5VKfd0zVP7y0EHEwcHt6ww6
/214zpdtOdtyWGyNNI1kjjpE/oyRw7PmNwsvZJE3V6MStpBGPlerpFwgjfx5PxWw8fRQkyvLsuk3
l9Up/xMAOF7D93M/Wlg0v7V3NywiQJ/yrm8YzZ2+vRP/ZfjP+TfWIChXBX23gwUpTltSUbxrPrQB
XdNKeZjnwLSIMmA8lvuWseZmCJAv2yf54CsawJzf+J4hlzU/2JDYLbnJl2Vo8fsnnbRyW2m8lLRA
y2zL3IsiwFZ5gfLmZk7MlWhUghR2lIsNU+9SmBjM/29d5yxoUOgaJS05bNwRAuWtC8voDpu7hGQi
0mxvHzgVojVqM/20NG4wCp5Cix6C3ct4MRcDX7ztcog4GMki+WrSU5VRLtgjsHRRTfFCidkWJwFs
eqWZZHUw5+u1Lc14cuVJw6z+lcidCumFNOhGZEi8/anD2hjJTY02ONjUJx2n2rEIIL3MVSQpppw2
mpjcKHdoErXFSEguk14fBNpqYTNdOjQXAtZ6aMoJhzf8CxAyWZCoCO2GwNo7AlnLl0c4XGloIAos
3tNjA+8YuGBdSQHud+W5eMi2uTqxMkH0m4tTHx81yQvEPrc9dvy/YwmLrWuAyI4WcuEtiTBKyrOG
SiRfsFcAT6tWeiGPyOcbjYA7lNBKrMfPn5MBVfto8rl4A4cJ4DfEVTdaXWDtJTrAG7q33KAk/f92
v1OENVcwBGCAjnLc17afdUzG8hU+ekR1CQKeEDgZLS4z/2mPjoWnNhXMC+rSMpGjrIRi8rbjLPp7
5/damh6KBqR/HUi0U8+ZReAf0pIvEzHDa6p4d/ze4eUAAq01XNOhvEzG+lfYIDqvqojPncAAZ23g
cV85LtM5BraOVaNUr6lqKVKoCkdzfY/MVblPN3oYBGDmID9nnMNgZZw4ChKHrdOYg96lRdtYYA4b
jeUtr9JMDGb1YPidXEMQ2NHYatN8pU64BW0Q9PLdOfRvA6d/oHc+HCp7YljpA4GQaXcAU03Jl4cD
v47Cs0iVRxkCU8gPR6IKrQLXe9oSHNEmoJGQK/RqpdaQ9x6gidvVMiUkSwimAMAtrGtMu6kgpyLM
KH/p86fTiCEBYNRkq4ThRy/XEaKExmBeSf4ZkwozxnFRgNqgWYXF9SeatmbB8/BBCjWx7ckYP8Rq
N85VCx8a9WJM8y+zP5wzOeWd7mjD3r++Xlq0Q7rCsef0Z6a8hBRGJf9nveUh1567ELA8HNZ9PA++
NNdgXatCY2iU4/BLCIUFPmbZHiePDQcnbH7aUXxJRikqM87SzTaQlQBM0FOqgjiB/ZpRUJlZ/wI/
NJsUMwCCeBcCSLSvChAV2xUXnc6upGqB1IUu8R25+qnessAYHSWmsEZQNcXGuTsfkvEH/lJmRVlG
GgQKwSvV2gPRZm34OCOVl9lJ4UyzdhtssFnDkImAV6R2g+Ax60Yzu7/OjRugU86Xlh2+/lfRQuIC
ogQ+vhta5BO5GJ7XF5S3inb5Uk+6k0nsNduFfHTJR/NFdv0lcXIdpwevLIKhImHDNdkZnfekqrLV
mfF4ADErht1TBPRqV853OGoulAWDERE2iInlvhr6L0qeu3do6RvZS7Y4Tig25eOPoCoI3HRMXIgW
Md3CLNCgiJrEHCw8BaDkDlrib3g6cnnM1PAJY9G5dpS6W2P1FgsrfyRLYcxMf/7bKUtOfb8CUCXI
tgMusW5Xl+EcB3DAwyNw6Ua5MvTjl/VDM0MkTrSBx5F/5qP5iwXqXd0vYXAhR+ylbPGFdc8GxNHH
8v2PnV81EJuJoFsr/oPVhLq3avvRHRKmwWUGvF1cl/jgBEJ4vbDBCcraO5pM3fPpONpsNXmggYSo
do3rDZHL18JIxiWBs49iGAEsrJbBvz2XNWE1J+jeat4+K82ytVQjBjZQ6qwJQv3R7lL4taHF+8qi
AoCV4UobmDwodqu2PmFtzYLOaTX3lJZEcRfQi3ur0ZcDEXWKOThhqTK39t6cCZJ5FQeWn/4O1rjH
WQJrmS4Ja38toTBpJeiNvdn0vQW0kbXyaX0lvZlxrrv+jbH5asj1PsOT6DVEPr26Z1PoWdca1SCe
HE2qAI5AqY6mIVXyPkG4rFE/ztC6QGykWvVmrw1q3gGu39PijquM34Ita5Lw99k+SgybPFbyyfOK
0Nqp4mE2y0tke5muFSb1wcS69MIPfrbxWQShXjL4FOYeuAsL1sAReew568svEXnmSOkrJrP4MTRj
lvgvsNaIZmngsIMzgbGBwNYAn/68XGfB+OOiedBN3jvskdqj5MJ7Rx3eHTT4b0AHoBxLDX/mK5pm
MP8oHDGdmPn57IoQHX2306mpc2ni1P9H7VJx1EYcvZi6I8H76W0viFTIXpqK/GaeMKwJ37gxqkFb
OBQpbgEzfZZbn0h6FPgviF36oXlNT3GBKzSVSIKQVohGvNOZomh8OKVA8rCIccUjbEK68LajCi2W
njqeZDd6lZ9TaTbg5PW3e3m7ZgrgPI6vfHrIupNSMOtMazEUfaw96KJd5Hg5avresRMmaOfLVQ39
lKQpXaCcKiZQrkSMLapdZbgR5miTT6zyayRM997dM3DLwZBvKqcDCrjk2eL38/qjTE8VhkVCuKdG
nmE2uIG69iIravOzOqqnZOMLnqo281wlgKnWM/nAi367tCGZXnhzqJmQbp500H/YcOv8rWie17Kl
9ByPqkuRiPHS1acMvWvdeuFCyxOqDZ+2vfRApcFTUNoshcmViWaCUdB93QgHvkjXX9xjFUfN6LmD
N7hiBAkTv4wUxq8TmeZqmtwoDAgzIT9ZIYwPcwCVBAY40PYSpR3fzC/jJqDuHoDzp0jKsNTgZMBm
vGqsKR7tGcgJL4DVlIuBjfSBPV7mwFQClisDJ+LXe5G4PJl7LFq2IEpTGYBQNJRzsZ0twA35jA2R
OdkUXCqpaQMLnqTfytjWtdTVzXsRKp8End5nlOQugxEt7TdXXGtm505HnHrjDW+mFKpSDtM7VivW
llQDzVgbUL3gzsLthhYr4OS/JZe+jSx1FLbb+oC9JhUB8YWfVCcrfGAsPu4lX4tFV/1c001yUPyL
2QYUwPmKTWImWo+vXFYZFNgPd9WqRB/sVHsW7aMNuWc2XEZfAF3CkfaOwj9LF8wGkBkKf/XYT/s/
hjcgvU0QWWDFdiBgHvpBeXfdZ553wTiE5zjhvespY7C/wYViYzMMECSWtpugNpBi9Idb2DSqsdW4
khdr16cADzeBGtSic7S2a7POLUq5KA6B1d+Z1BmX2cOIhAz4SaqiUCDWnEDBDT9AyZpZUTETEXmh
vAa0WW/CVbvkCK4Fc2/MrnUIANwWDT47TRMfnmJiMlC2120lDW8bxEx/3db3fV73FHry9tuOYDkh
z/42NNEz0zFRkQRy5AmCzemL73sKQb9S/2Ih+U83Wd7Pwm+HK92s4iCGjH5xM8Qwq/Fuw7sEM4f7
rCxEtzTlFedLIQ/Q1whY4t6Z2A9S0MlQOk+dWEmH0hsILMYZFcHdZR3B08HaUcTIqYFHpLUyVzzV
EArAUXcYWJ1zzKjt5s4jBox7+M5r1jAiZqYaTewlElJvTn+28WyQ0VloFcbc7hxDiYuiodqxJkV2
qEYN7SZ47ENTG9bBgNAzx3hOSvJ6JdUZGSBSiBOODOBUPoiMURGGvtHYHn1979bLXnInHcAH92oM
KT6TSG9FbZeKFF0l0f6Vb5OW8oGiYrZ/X/F3krfznchbqjc+BSSl0aZ6NcDfyxWnRARqQqqract+
FH5kbv+icXu82NXklO8edjwhpL7+NMi/1J0Sink2i0RToaDox5AQlaoYB4RPFX0DmudBEx2qt2OD
Xi5dpPSfbpo/CzpMZY5h27Q07CUL2b43av/elStpA6dVAqDDsWgoij+NkqWGs/8/oy2eDttSoKsY
1EetH0IuOFrhCyasagxC/nBBM/ghKHlSdkNfGQDT6jDSJOovHYQHmnMfHJlfhBtcITQT270gQnFn
CWE7ZnVCyjxu5edqsJw6CHVX/tBtP35AYCbt+OAlId30kTNKIsQicXLpxhjuoYw0bnc1C+uk4lNF
EanwgbhPBJHKNqNr4NWvnmEXEALhVMZZqQs+dtNOm+EC+ksP+Vsjt3Gn8iIxlIOZxx3cWfG6ke91
O+3aQUjIbGSdBBSL7omH2jz1RRrqD6sswPM55JyVvqpDke8iqkEzHKmHtn2jAax5EhrURxTNgAn7
DleX1SPUjywZzibxoDH5GvTzpL7i9o+VnNd+tas5snT9X7ay9BT5bsT5xpYjw2LN3/TC/WKCpz1l
QquEhfILjKpKuSD6aLpgtwHYLsPZRs6ZgPqplMB6crqkVcidhH4EiFwBfelKcOpImhMYcJirAJXP
1gJ8lF9shfmD1QaQok/EBwGa65q7zCJtOt5fwPx2W9i2wJFWlA7PrcG/FsSSpUxh2Q2vLxOv2BM7
QulizfThDoH1YEbj51ssvObGrE4hIQOLwphjgtFillWBJ/9uTgsD4YeY0x1O2UlTFR11xlNxH2H5
3a6dHVGT8xbF2DwkASUqwPQr1YCHo98KhrBdMopB9lrXrmfnW37Mt0yjhqBPu/rQbdXb9blEoMuE
7WsIb15kXlMBKAVzdTY0DpcUtirtg6ockJyx9gl9Llt1nIO9Mca4FGNQBUWIoxE/HwdAJUh0DSmc
M/zttAaDYFeSNtngrf4RisUzh375+Mn4ItRp1DiPxctG/ZekWRNHTNx4DiHdoSgm1IWILa7SWCHP
qj8XkEY4FmRnQ87yBtaX8VPz2VWepmAPv5Kxh9skxdG2kVapTncrQe4PJGE6j2CCfH6P5mbOvuNc
1hEuyfm6NGIK40WkGOqBJVmOzs5uK/TC9Qi0pkPNY1XwmJ/4ZyGuWuYzEKdDrhOq4nXF/68IS/TG
lnwMqMZsN8ALxNFF1/w5Ad+Jvo6u9BUtF6plt24hPTY81y9FWE1ntPFuHWsHKjZNUoRytFu5Xk/N
/9UhiG6o8NNLRNFFfgUTCZZxPRkNtojne9q5m4+p//k7XZ+s18RFkn45sl9K4xabDVz77+hHBU8U
TJboLupD9hKa6IfLRsGttQ7gqQBK1jmkj/6ud5nQueU7NfZUjfY+Z7M2Pao4LOjlrNDDpHzR6Sz2
tth3CiU4Hul2o6GtFe+LaEHX3vpwRzvST0HUN5wxog7USyMXJBqPdL6IbiGk8L4c9ac9sYIXXMOL
+MrBhV6dVTVYM2+9OCS/DfXWFQTlwBNCHV4X7ZILC0HrmXITp97zOQfiW02bAXylAgqm1vGpFeXp
NZPxdBTJrlbmCyjq3Zx2vH7sQ7ZCKYibQY7OChxxRPKehQsd754R9KzAG4/v1CV+ubMj+ouYDFVc
g+NZcZnVJGUHNBfyn17wqTdKRmk8gmuHH44FJfGet0+z7mjik7m9iHQtmlVcy4YXN2q75hPg3SqT
PL9jdKotsvb+zNhiHxaNzYXj/6zx+vIhGEIvxeZN8iRTByrzucenA6Ww18heUssYoLwJS3iWGqNQ
theQom+BoUijKWCGni0IjPlWlX2Ezs5+SH0B4DJp6qM2wVP9zLXi94O8+fsR688KWI5P6yO4Ueki
8Fybul/tc/2Duj6zxYalSkE+kJoeCNp/ah+tkWRHihbqEaOBZ8GA+ZVBFLVTyYmkaN7F7mJbhYDt
lg0xxxA4Xbn7FQ2cSm9TT9G/d4vOCkkMHZnzJpVVDPP0Mjl/EPMyG4Hp7eCLvKNnfDNRlKpcrlkK
UY4rI9r9R90OXPm1wDZYdXIyZiUtG66HkRPxxojJfFAFn8dW5zq27AwZBSM8cILLEY08XvkVHVCV
NV/xxVnVMmvXxTxgRQeFbU0e6nkCRXCwvCEoEhBTVMXHkexYMTbpCLCruzkCg6FGBuy/selEpULr
wSPdKayGNvsVF4dgZ50eTvpEWiR8/pEhDBx6k7FZ9hMlFbZR9FDHFbtSrn4BaC+AiUFwoDCTtM1g
+CspcQTyWF8DvwIUKlV89sjsJN4rVbTTjMstGDYKjdvnDsO0NpWtH8zMC4l5Sw34GWRG4BRlz6g7
v0sp48HP023KjcfkXIAmYEIiaaXGniDvc+BLgt8GGqQ/ZCDYKeeNl3ZR5po4WvaFzHS/im45NhPJ
TF0F8dNoLsdVrSK1T8CzhI0UG2fz7EL0CPv0r+wjEM1JGQEw4VWQTtRqtVvZkO+dM3v90Tpv0srG
ZYmA5jNO3V2YlrMJks/JeaxXOEE8z7PBQYrgNQ+6sA4sf4FP8FK+GzilVTpjXVgG+8cPL9l50owt
2dlkHCZ4AptyUHvG7yeH79Z5BjNnRoVBZzKrlD8EQS3j8Htw9LDDLVYUt/e0jDJEZWS/ws1AQq7s
ko4i3MFTOeX58Qxn9n4Cr5hzJjigCp5oxGeDK5rLISYChc+YV6YCuh92cOCZGib7Ue0as6rcW41g
DHji2bhFI0x/grwZMcKSr6o8NLpSBCO3kJCyorOicQxIH8+VArcm+FSme/CdNUnlsKazFsPtUvXL
dsP0dD28Iu0sKx/bIVHIZ9lOldh6kovPHBlEwCW8OXQYll/DkA0Tfvcz7o/E2gCarYeAwscF7hT2
xO7fRV7iXSceQ1ImK07JHwBV9VIy7BE+AycsBX0y2vlZtMTvUijYPyaBDmEntfWj10HovH5HKmty
GPjpoPlM/u4s9JTVbUPFCEbwyvXine2ba3jn2l0r8wx6EMgF0uWXvaktEjlkiPCl5BbLsTFS5Bn0
BM2V6lfze7HOgxlYJBx2IhfYEZe4qCs+kaQGXS/h7X27vvKJQtxgeQSik3gbsOkjCYakemjo9APL
Kt3yLltVzEtHkjfG3kj81U8l5R2sbjmKRIz1CbUqM3PiynXhHXyUNMTajVdXXDLUbUxgYHqCPSli
K92rIBjuB6Z91tP2UhBc6GldlS9yZU8a1cU+o+baqu3Rx2ld8ApVsKAGxLhSLBeNWBPFk9FhDn16
sH4Na7PxtamhwYfVQvgX6Z0c5DhjfKCs3LeXvV+s/oSINfXCZQSrLoE15yXMkuxpOwzoWapU41+Z
2VjVhV+xLl0xabmR/S9oyWUZA3eQbfh7RKN/N67sh3ES0edaegzag3DYC2wynvL/FMqaWsPYJu86
+plM7oaBAia3OAagYqRmyCcjdcGIIpocMfanRtO68VzsjJux0cszGa5+4VvV8wiUjKdo+pLdBVBp
M46i/XxdyfV1yB3uFKvFgdKt9cCYNqiN9rJ9fhzypXo2nlFitOTALEH5vvNk0yu+VFmSeZ2ndpww
NPX4m6+9YeBkZqeERj/N2dntnnGTFZ4mNDs/egrrNJg1UUPXRHkLPWmYd+aZKOoo+KcDc2Wq6/ug
WqVd07aQbplDkqYLfndwJua084RM5xeoPb+NjAsx80UaC61yqugun3ASYoQnXrprbIoDjbnjhli1
W5MBmIKK4uvmZ8q1pC6Anm9x+t2QYP4/4SBi1GO9/W8RBHSKfqQqeQ5lLUxnQWNP1b9kpi3SBao9
KoAtwgUVcfWOKkTKGRVwqNmx4lgzamIjElI1JzK3wCSdfmoudYuiDQX6Weze8aG6YJR2WUwM0PHJ
mnc36LvDqES4eVVa2D90aBWRMFqpt6vDM6gMmrCJGGvDpZYrzuugyIM9Q3ATV0PFRXjNHCZwon+K
KFmwD/Ch7no2tjQje0qQcFT2IYky9uOYvKkC2ljGVllPBbF6dgZ3Wk3mR7BgJYGzHDwbR8S+iHGy
g5xsJHzOe+KrFyLkmD3bOYkNFs509pPtiVqnGgckDylUIMZbnMonynj8NWVYkdikNwMpBlC/4ySj
RdFQe98/mSD5j/JFsDDvPgu06l2qmEiUztIWEnDTcG7FlyIZHanTL3981LktTrf1lYp1HfJ3/yk+
gOSTJNJtp/4du2SK17vA+B79SJXVzt85Jej1TU7Z5dX9zGjPDO7ehvJGAhbk89CQzljHhCjYKtZL
bcTWM/uAFax5H7BXfP2XueAMg9Dc5pyGnyJSBq/0XDEpZQEyVPLWS+fA6NM0E7qr9lOphTvU7yBw
Z3wwILMMihWpJI7Wq2v1S1gEzWtW7a2/h6+9/GEEZEVxVLwiXLX0y7BhFuPwlbwE/vh5wKsYHBEZ
THeKg0cjStsUBajvVK5fjFAg8eQz5YB24A4wNQENY+DaLkx8oLuFR2ap2oyN9reyrILBJTIju1iW
7wbEb6eNgF1Q8FIFRy/m+kTQwMIk8wAdLFZrRcCvnb4UJiww59EqXoMeV/rpd+sapbSIBO/s3gqF
fuxspXE2i+N/mPIQc8a9q2lk0K1JT5cCzQLW9mmT9ZEnsAWy8Cb5XlrovUG0HQfKVmPm6GXkd6lS
LN501HtWCo6ptZxkrjlNEOiG/CcPzxEQ/vN35KkibndAbdnq64oiqgjWJmmpw/4m1xwKJYOU3ZKa
feDhB7THOXG7/2QbqzeGgww7Axs+nGOAjzFfu2OHdCaoOh+rMpNEItXlylId9LtOfuAUz5GhO4xk
yHTRCWRKpDsUjIYxueEsJ95ufwX2yCb+zHHGdTh27cAVin2XAjpoYdayB/WqyAuyWFqZOp8FO7On
FzZRr3nf8gJtfaFEUYeauZTbjFGgnfOIKqp6CzWVRuWxUikWXjXYpDHb59q2sfZTR/cBaujxTbob
RJHSP8T9rHQ2kD/bFaUm8OnHfdxJy8J29Xkh1vlyKzLm3on0Kksxc39bdEO64wVgei8gAaC1HP6A
Y2EyOtfaeN+dxgAa1FeVAXvSNu8YS98R3YZ7QhPP7geexxDmEfrhcKcEtXK87HyDXb2WIWkoqXkq
lWFri4oUtIwun6zZwLfANvjDewSTi/E93/z7qHJlpHPePes65dINVVx4PIm3aPBHycbqMH6sLtb+
x5+mpUbafpSN8Me4RMFtKnaILoDG/NzAM5xTYB0Vx+62rfSx8h/nZkgkVIIphzEU3nFUcjSKnc3i
gYHk3qko6v6b+w+07nQMSBJ+62jKmTHhpAHR9SmXd3UHD2YwxtIibwBMz25yGqI2h3MXSmDyq++a
u1ciga5ka071xvt/Z4PbxlkpUSZjANvi7/kikwYqVYMn+vtFavlZbuKvEx7nQAo76c5XsnTwsuwl
TkFh6FYJnt/daw4iilp/j+0HNY5U9EL4ErRzKmWZ/WwM/yNOjtEGhPvrWaGQZQVuS3pmiu2HqQJ2
afadshLI/VLmfd+c2765A2nenQVqfMA6/zjgwHaGSwa96CESg9w693Nqvq/KUMxdhGZbeqBijzir
gsJm/M6n6YiO5Mb6m6xC4LILtvUlSxXr4USiQW2JUs20qw9psbc1w91bIOX8MLCle674B4rm/igz
kwJC3VEP0roLt2t7X0G45g0C5ge/DyTl4SEdGDwAfZSWflY+/vzEgFwkWt45GdziaNyG8noLCdkS
GKjv2ZEGM3u0cRabZPytvoFDWeWYb/CxHOsHhbcN/LbH1qAIx3oc6yCTpUOSR/8w1F/eu95K7IUW
jTZlGfDk87v29gK1N2MQ0LR//mV8N333w73lEQKJ4TLGLBVPQXdHXmgMxqpAMFBJpaqxsMoWWny+
KA3KOaiEotwf2gsZuUn4CmNAgtVx230ojzOAP9m7sMdOAjTry8ovgHrelYj+qpQrhxXBt/v5cWdM
WcGWY9Ir3Av1UHd4sFzKC78rOMJiNXu/J98L39Z3z1+TsPoOS02SuHFe4xtjzI7s5tkHv2vwy9aU
zZq5md2mOnPk8H8cIykYL/Jb31aOudQ6xHnPEwxqw/IhyRlCBYrhYoBSWLymu2KsHyANGwgn3uuH
saQw6LdJbHGsmJ2FP41aRz0WHYXEA4maJYNHKz66e69wJz4pNwWrvV9xPHnxcVYpp/kpK8I6cASp
YKCtyR1qj8bqf+u4NfAYQi/Xgl3HPXaokENxfhr4XotN6evgXELsf93lvbIeo1VqobRGZDoUIQII
urxPb9JpTRX1mC0m8V7pakNb6fxlnvPIjpKgcLCte06BbvTbXYBTDpBQ6CuF4loELW52itaZZw8U
wHSlMMqeS36pOfEFgHFCB2rY7ZV9eVVcRTXa0C3q5JBWOUnU9L8e4oN0Y35keZUM8oa13Pt7wcsf
SvjPyJDTHSXzMsQesbjk5NUGpeGAmOkZ9dcvhnbwht28/He3tHW88URykceLuXhKy0nNZaA3J29/
ixA2ilzHCztjP5KbuGlm1S16lfrGOurJA8AoOPIWW4CEzUmhHSOt04vyotBW5XIj/51kEP327PN1
TCoAOxd9CrYuchjqxrCU29iDL3G9t49DzK3vXc+Xk2gNNXXETbMBEYpnG7dK/7hLs7xW5jZ9XUkM
9q8arqltxM/RagSS+5seNE8rslU6B596zo45oyQi7jmQp/+l+H6nfijHkqfBLFAfYuykQzGFKigy
CeneWkOUE/YfRN4TDMcwjdLqR11B3EY9CbstOPciH1X+U9gfPVaAzCXO57EF+XU7N6jzEQrE7h/g
9SxXGlBYAcBLLHh+OpD6CVEL9e5XIj9w0MCT0gDHWH+T8P1xZwY4dpcAg1wJaNX+rRXNa8Hah1Y0
+OkSfKlTgEK4QKe/reY/cqKEtgulwsfugqS5D1YA16IiZKBGLesqX86UcTi0XMTPuMPJy5sZYs8l
wtmhmleB5KVhDO4rUhVzTBPW2D/rfVPuZJ/5vMJ6T3zdyBoFR/IXdr4uJMIzvqwAkTo9Lybv+e8f
aOWt2dumdEtoLeV3sKt2O9UAcoWn36EPZfm2hLuUFdUnIcJ4MO1pLIUqohGobrdjr+bnXvHL7bdB
j0jrYwkMYmtHX4bISghyXMkrn/OWznA24xipgCBXA7K89JsSJdZpS6VXKZenKcqnTUm6q+suCXhT
oiVw5KwGtT59c5jTrp5XGwLP8FvcYXF72ORdl0pFdkh8ablzrHcelcRoljaMcRAPpO4QIeJThXtm
Ayumpa/+IIn5gXMl8/YWFIEu9YY9xZCas3lPktmDdgw+Or86YchtCtMRmCecKZPv0VFZWUPV01QS
6qi+zrYLKxTBotQWLEFEuYUUHCDnG7CxhEQNtPK/duEiGpmynI0C+kYccjWw8BcjR9z5E5v0zvSp
W2bDY3OYNmRBBjnJgkcmnldGyHW/EAIudxbvfVs0uCU1/tDBFDSqSZqP4x9P1Emkdl/Zd9BsAxMt
F53Td8eXKuX1eLi++AS/QctyoCrxZ1g1/m1ZJK3D8kwWozwxzNRUKC796Ra/SSP9FOL9IrpKDPWt
AlnQ/vug51EJ4hlCp+yKvR+ryM6I+2DTD9S0SieagZC6YWqRMEMfQkPlD0BlEFrj6BFObgPIwjwY
57cGdSUAI44e1YtPHMvJGxXpeeyNJaTW8f4dLM1sQTNvYxtKTMDPvi8V0jguwWq06eMcq6kIQQEj
f3md1ABZT2C6jonLMrJDUz763sTWN63xx0e3Z88hU3PFXiHK+N7htOIWCq80FYb+insOOFfXDibP
ycq8O397CE71cBGGezLNgN2Ok6eYoGNHGNhjMjZ/b25NvLer03iB3U5VHhIeNg6DK2h6ZPXpzkjz
Fw9rEFFbme0Oh8gVGf0cnKASSRMpDA0/m8ApfQlA4wQNMsJzw8h32fCqZyLdKz1jNKsG6whAvevx
eJWGLVWBS6WhbHKFkuS5l5nyr8dlwebcw4rHXGML3JLvcAdXxsMFHAaUcGjEUDF+ZxKRPtunwYdz
P8IgcJ59UkGL1Cz+9sg3RbltLuCkxh2XIi29tPAfaHnivK/4v8iQp+KDOhYKANNAPnwngFkwnFvy
ROeyjOjlC2GMdsMyprlGZ5h1XiDlrw5lPmseWobvIalZtOCskqYrm+6sLZFN5zyS7JUNhj4ocNyg
rgZN1v40DpZfIu1JdRwy6282HQrQtzs8bBILN4LcUoVAWFPcwJRtTakQrt/SXLrvlyv3c0yN4fn8
z1k28u+z51vwqWdEi6anrE5Q45l0vbQyjIEQUm14B8I0xrTS9F4z14PrZR91xtFAagNKmyig0v6s
lcxuz+NdoCHExfRCxRPYkiOM4M/kM//WcmOA+k5vvPCKBlLxWOgeK7uzSKk1iSC7a6PVQt8qOpQ0
rYHXNxVZ7yuheyqXCBa1Saocsu1HsSxuBsVLteIq7bjU9Ero7QcnAm/BJmhjTkPaikXBQcLZyUGS
xVbahPMXMDSAsH6ADMLe4+nSZaWA1FwhLRBHcl9CHnj++vsaGY5xVx0rWbz+6nIF46qScIHd/5XR
PXYr7dSO9NdT7TUvxUpiRTdSUGLZgp4isLD2krYCmbh2Lr27bVLzK3rBwiH+uOBK1gXbsBTC5vE3
bwgAp+337RSr/QqOtU2FV/hUTa/vK7e75MY81If818l3i9X3Cbuiwt1I+06cSnJgYncPMmlJQZ0a
+dswhXycP3Wk8+w7G1QyGBHLIAfy5hSaBZ/a/hKpAi3zHGCemC5lh8xq0qO0uQ77930HF6RzgK30
yzGzS0tQ588b7QDyqoyBTaoexXJ5X8kKe4OZN5mte6PPECvoePsKE6YNutuzgxzFSqKvYk9OxDf6
xYw7sw251yejBb11Tqg1fYd11eJfhGH0dHPyIfJOzsgGy2glSQpEdpUPp3gUmalQHd22VpjrVKgz
wwr90550cOGfHDYueBm84my75WawY2RV8lq31VOQxrJrHqbEkkWumFAgkaNaX/nvAvlbhpWXaSNd
rNJlTdHXmzCDUUNDg3+r1PP8ZtMKivkW2ihEl63lbwXwnkFDYQ6OQGsdWyzytcd+e6izirM5rTtq
Dvb1mxoHvYFIBhaiyM43nflAj1sxtGIkTgGWfMmWCfYM5Y13S3+1hrzB7NWv3WLWPnCPfN2406TM
dU2VN61scZ2rbcFUB5R9+lX+DgoTIJOzoeZKSCxrMOCfsx667SwaqmgYJFZ7TD8Wy5h9YJUHcrZf
M/5GIEATTl5W27oNbRj3PsbT+ZvKnVBojpiVlBSnlWqwHtBT2i2UpN5ORg5Yh5RrddwA1zEq5/JA
KlaiMQTuJfJ+DXz9xhNbRH15mBV7zdgU563wkHw9uxhMrwzO9ZAndiQtks6WTbDhqW0l7cOcyWlF
DkljMcorpmdWPRle0x/jWsHdMHB3gN6NqVNYYoQU1/PzgTvCxOrmltsNk78WGzI9fl1WZPZ1hEB8
0vs1ASVld3Mvq+PaZpgekmaXMoCAz16XIPIJ7E7BUS64zeiDnkMuLpmVW3zE2LQd+CH45pf4C0Ne
qZTUq2upEfi/1ar3/IUHgq7JU5/XqO+whgNt4D4SqFf+zpMCwkhci0ODpZR8xQNe7Eq/OLOxVQ7k
OVq4WxosH6A/58429vZ0mq0uVO449WjHaDMqOJq0hShV/PZhCldIZ/0rQ9iKNF4Kw2SjQPMuTRtT
GEGqShsTFxOH/i7D3VRvk76tyabwPJsljI6GKz3E517noa7PD855XQZogFc7gnTFVcJUoypJiQ9B
xny/oPNJ4+u0fQS31CU7CV3Vc0r2Tj1OzWaNgPpG7BoCKTTbYSBFmpfNYeKfCOEsYE40wDHN497Y
CBmlGGefPHZITdGkmvl8dhiHplS8ln+l+pEPOGv/QiL2Iw73tdcgKSC7+fv6IpBT2h7W8NMKm0Kx
sJhPaFKAMfZrT6FLS+fbvu126aSpFQkhvkEH+5uz1EtnPlcJ3M1kw9+pl5G6IRq6tK7R2iFnx7KI
Nv5uRwzjxKCx9z749JUyZZ67RUJCP7ZjlNTnqbe1gznINj68bYrIwgvaegysQQBHVNNj0LaUqFke
eA+/IgfMHC+xrBynRet2Ibt+pLCo7SWjQ+qIHUR3kQ7ZTT16Se705hJYgLSiuvg+DT83f7HIBZ92
075ynda10ExnV4sRQ6/tqGEad6gcl3DSy0b2bveU712o+JALPlf2Q6x1tYr+1E1a5G2eFcwc6sKI
HrLemfTJBtTSbWzgVjwH96Hk8TLH/pklt0+CBKYc5enxHRozNL0swTgWuiZExnFnvn68EmUe71Vo
rMtB0/ndh+vS2Fgo8DuhsWEY6uDl0yOHV+m43W+jxlvTQ3unnBu8fPUn6Zs/5IisquGZRRZ46vVY
B0JRxLhnVP/5dCH6pQPvcxg7xIbSCOJpJgsu/iGvuYU6HN/4rV9XaJpsczBwSer/HaIWjgH5dnZL
qgdS2Dp5n9Jj9N+hFfxL7QZNYwMnj++6jrZCOzDShzr6A7TB4bp2VBnLiGJUAtms9EzP+59GkPGP
hDu+SmXkoBKx3auFFdt6qiLHPan+N6VgryjxxwDitpXJcFifgOjsvs1h5a1iN1iplngOKyNaWvJU
dfKJfEbNltF/9bFgycYhBojq47UQAo5EhaKa+/gosxbTBvoNE4aZDS9B4GSxeeitIeit1dSBn8Ol
qJP5M/od8TSqlJRudqu+KsL5fQzomzw+JhKKSOklZyzirfWIax/X/OWFCgD+pA4JkfS7WTlEfM7W
yLQJWWC5K7xrrPvACGwIlKni/A6tLU1rVUkZX/Krm99txdI08V5FZahY14GX6it7PmltWvgXmyJk
0o14D4atP9l4Ae7lwBjNPJR96gpmB82MbxmR9MGcpytFKoKP4GgDdr7d0p3xOSh15V8scd1eU9rH
CsatncJH8v/t+YFIbVtozB42Q3JFyMkGjG/WkOg0kQoL6vCuQ8VFfjE4L9dwSoCvu87XQRr+xBQJ
8i/yIS/CJVPY9CBzmIVL+Yp0k5cFxC9vBf/5/6Hmmq2GTiemanrcWsSbe1uiokSP0a5pe3jia/gK
0i6k2+llVhIM/6fLznu8XJ7ew6qka6sQDQhXIzw4jHqBSZMMi22qgGEyBO+3x9tcHUgVX8agmT33
kTGs+hVMSRCZrywNPqAUzmTSPBw80+iWnFMLWDWLvfT0OeMlXR7TTkb0+UETWytBi1PWbM7KjHRH
VeLHmejKVMD91Ky0MnQ7b4Rpk+XS9eLHGVpToAV4HmfKYZWLGdmeotJya6a0kBUEqxiuVSVvom/l
VrvMmJNN0OCQDGa5IkifpNmCWYU9TZR34T9sfc8EAXaC1UHTzqqb/Y/JkQOPlNJmdgLcmrvrfaHk
pJwSmLWAcq7VaMWjA3029Y9LSX/0OPMoLMZbgmtILTWkoCuL4eoZepfqdsnXhkzsh/U3BPjzqV7J
6A5kTbgCrwbPp5+v9gxsVsmqtKoqzVdFjnGpMNuqBmptH1HYcN/SGlXNxGdOeN7CbIxLTpUT4LEO
zJCbT4cQ+az6ailaGA9aQhKemj0+vg14x9WdJd93XCRqZskj93zrqvAUZGMCwWaqaFqx9XQE1ArF
/swSaf6CqtEveDJsQpHlcodKIRgQ8FJFGBvUByax5387SBUXMzM9Wih/ClNf5Rndyb2VZGLvrVVE
rs9gcoCKacBtwXLKDUCEFOHD9Exo6pffPjpAwoViaHMwmwDC8WMcVaR8E2WESKixl2Axl6bf9NSD
2ptfRClgILuLa1PTt4XBmNwAYLsYQL0sa/P0lPoh1Ul9LguXkkmdilp3N4log9AfKbnrYkNEzDPW
eVnWfWUaooXSiUu61fzO8MBAlsWPuxT26WVcC3X6LGiDE6rN9cI/lVUysC/H0XKZHLnSZzv9j6iP
wkEfz1XUdozL+wkTyy6D3kgRYwimTdbmI0Yu0KF2M6pmS/qoARtcyR3fJyWezZxJ0YiS+zqZm2hd
qrvwazZ9bA+ueGCCYb+DRPSOCDyndK3dxo1GNGXwds3+WFnq6xMCjiyIz2F5T/xPa+tKzRJU/U7i
MGrwCEYN1rixiw1vXHo8lyz8Hak8vLt07c4dbdANwazRqpyP3bkrqZB8EauFl+BzI8FGflKGNGIY
7e0FyzoIrs+LMaUXVImkf2g8rkMnBxn/FP0DLJ9upAu+KajcYfAK5qcQOGqZBxqKs2u04OsjwZfC
Il8xJtL/CwH62C/466R3RFf44Y8U3tSsBHjtY2Rb5ttGeq0SWASR1YGudXq8xjys7SNn4YefIFzX
jb/L7hLaqwEQNFsZlJHI+pbJvG8nvzZxP0bmG7pPRQaAmk6tg5DgqczguvlMj/IaRb/BS9vhf7EN
0++hYpqK5x4XJzezgse86Xbr25YxeiuTlIfPl0PpftvVWZ8ODWbM9k3jIBOIVi4ITBYNSvlFjXJ8
/Z0wqA6KSYMMzw9FgHut6e+ttn/1aPcneyxz35Y5L57WZDaDgnePkkYzL5vP6qEBtFwsP9Tb7Ziq
3vHqmkdMUCCFrlAaruD0QCHrmMZ9VHtLGo/AKIvnl3GxtFQuEAt5Kl8BNRzM6UI6wcc3pEP/tBr/
sbeN2HF1F0YIWb4HK9j9DjmvtUeIsQtErr95w7mcErHJYZOlQUXpb0jzqdKakg53pzh+3X9MWjE4
gMpQu91D2Em749dVpe8YAB/dlqxvdw2x7Wz7A4MMpWGsOMkKWboa2idgRwI0aDah12UI0h/3zv8S
+D9QzH45XsxxNnjJXsmYsa+QCqrnZt22k8zn6ni9k5k9+N05J9lwInLJaN/fO1ut0KMSyVt7H1sa
iPPYBe1x9EnAAycOCUcFQ2VeveQPZq/Q+/Tp9iPX7N9aipq7ZesTYgCQkJNgyzuwvK7jEzcFFY1j
sYYXtR3gxYJdAwalr+jEf6xaYn6f843fvP78tLD4tUHPb/Z+VVIHh6eJBMLYWMsjNCkmtX7jEnLY
VqojEKHR6y7I5sFqMuncntSD5LY0iIBMVEr3EAAryo3eepTSfyL2ptVF6CZ3iguqT8rZl+c6sP0I
ogxtb5kDQetnLh0aJnHGDMZWuJuNw+8QjEwzzYSS3QN/jCyeM3dpWd6wteDBByOYgMFE/1iSXq0v
ms/JRnov6h11Ca1eUI3Por/hcbh4+jz5QnW8a7WKasp0Kpf1HTyEiAowMfAxsLXEGITxRbX1uX+O
yGSDUsMnJ68x7qSwPqYA7Zfa1zarkwutLbBy4PFQ0whkeoB0hRoK4fYv8tziSzGt0wlEzRrgni8y
daFS+8dMKLhzxB6rA1awcKOY7l72gPdA+Oo81+NZEk5uEbyL/dX5a/+BXd+aUEURNPOQylOpasST
bOipY2iEXET4exV/DDQUdBF7RGyyEBhKWx0tRGkKYrGkXr5Gn1QNpr+O+UVsQ3XKlXAAzx3OKo1b
2f41LGVwnuRsozJFZSMXE8VDUV1bmLO+OxftfzORUlefurW73MMNH+OVC4NEuwcwPeJs/49EyxOw
szhvAxnCUBX8sOkFZhGDum5K6ztNplEnLTk+4MU0R7+kvkx/ErZiFASwokOtrxlgVeNcniS7EqM2
ICL+zBzNJJSEIvmB3Pj6BQTfMmFihXUSKbIDvzMLlty6CwxIqFtvbwzmfE/FmI2wNUSx7AjN1Cgr
IBcPlZZH3/uup+VCwN33tu9KddO1Y7DPEhci+BP9mu7Xd04/2x2UPXr/8jjFcwrvEp8eARZsA3oL
3bcWtniSRrSAvQhny6q0CttFMM+LdLMj9/vrbaT9Xi77kpIEf24ZIsgZbELYJc+Nxjm9FSyU90oN
6kqMzJUnpwc+A7kdWL3oSmu+P24XpKNtF/nFlaMdL1rnRpGUsZmhbSj2o3TNa+NoRB77ZcUUM5Aa
PRTx6vqeGLES+pQwv1hyohW5vCsx7EivgKcV/PBfB02HNVxz/APTuzDYV4nTlMjyLHpUg+6vqGve
xjUDlf7ZYMIuYskg4B92/bG1ocD4Fe9Ma0S0SiKBLFattNI1tOqTq55pbNjNIMeBILs/TMJMAKFc
EE6JhL2dLpk9l0hGaP0aJcr0QrZc1v4QTfV9D2LHxvgAnXMdJG73GvY/gWXMlIIg2IW/1CKjvZ5Z
LfG4D4MTHAX1ucj22DUWqg4D/p31bXcO398rO3Ff9eRlqjOqlkdSmiapcF7NH0CZZVhn3nAe8Vi5
1f5UGYqIUl4EqhuWJlgRP/IM8uqXLDg9/PyQXZdnNVQcAOlY90ItT5ZF//+dL9Bfz0KSpZ2CGTqP
JH93unADIHqg7LNPFrDeKXyCccTQVtGgZPRecpYjj9AhdvNWzSnh2FWldz23mb2WmgY8DQddcue9
W8WG9fj/J9C5VexBIMMaVYAgJkodKWNq0U2B7paMDMe4veeF87TtBZzXJnCWUPPiPoT+MsudHumm
M2ANEiyFje/iG8iEqwHuK50y4TLkWRrPF7px8oOrHCej+jA2w60vWitFCjiFkzJHbAwbhQziAiGm
c8092KgS6tY5P1U6bhvor3CE6PyFMuw3ZO1Xe9A3B7Nr5tVOJLhHUf0r0U8C68fB0Fw/SFynz03q
bn+cN3Wny6Ck0c3Jdji7QnWnLKOhBl2nAdXDVIM52hf/IXpX+seW1zCcL1pNFnW0yFNXK/ZQe6ze
3Hib3+y8CKFy3VYjYJgrolXJJDBccKncEKCikAfbcxKGdAQht4+XSemvQ4e1ppt9W2MhFCN2R0vw
I6fvBwXilarssBTKpc1l2c2gE40x440ZntL7L1CvuaYjzccTpfWJjT9CF2jfMY0NeW2cZ+WtJhwM
oGJ2hXY5nJiN90WIN5sCFVoB9CyAM5UN47aPh95T9oq4ZvWMS9jBvGK8L60E9mo7m5frDXOjErjL
5EsLq48JerTNlWhKgzmglu5niZT9E0YtdBhw+6HfErc35AvQp33SC4s5ju1J9bzR7WsNvocE2TsM
uvmE0sX532/n4kCiiMbfPxHaqsrTJSQ2vSQUrUis9q8Fa/7jeHRGS/w2uWl+JXsLoYbvF97TDtQR
g+ckp0lqLQa/htx5c4jqvgj/7h3FCWWS+78rKbnMssYSGN75+GoB4ygY4GdtTLaP+yFeoY3HJfn8
JiUlNBferUdxwtj46nKnezTacL4tQmLTKEjjesy8gCM0OffRKbLkby8EyqiRfzPpEPwezdaWqHud
n5WaAfWb8I7iEKdrvrBeBlg+BS/uJkPzbZokFY4lEanvSBhQ/+pDPi8SOjTdbS65u4k54vKEM5Mr
RF1FNtPuzVlkZ5hKFa0D0lWPUu95yYjajj4mC64x8+WWEm0/QIPlNA7Ckrsiv1NRQGlIfpe2FElk
2ICjh0BWOHzlcXLOA51bFhFtjEaS3lzVgOLzELY9R+/0BsmIYvbA6eoJlup4PGiDCTHYdeAr+XmB
bzWqdYUVEoStBjRfICxHZK1b/vNFGHwUaObQYCRK4+huSf6r4OZSgx/51aa3E1yDW6YdOhOxKgOb
WL7/A6dVcbKaXdf1KV8r1UI+0kebmA3jMPi6n5wDwPybov+/sTgBvKuLcHZU1DjWHoXs0wCJ9vRE
c5vi7iq/sXHYGpltfGp+xMQK6WBcqAQ6wN0SHbbRagmamBGlfgAcKDci7EjSq0wXMTDbKU8AJ/OB
/ocZ5TJP1ug7/h3Wdl0I1gNAj+aiN5vQ3UdFW/Q9CtezCrkR9/uNs3ZGxofWrrEQunFyESi0pwT1
9l00txNaLF2D+/iQ9wX8jRobHHf1Y4SydoaY9toVe4MhTCzduq0caUF1OcA7bgfuN+hTLCM/RBbm
qVXukx39pmu/fSFs/vDPXwwLUboz3kZFw0I8XB9rZQrm58toYJS8JLIp6faUeBMcwrqpl7ppmUNg
lpjRCKI/t1B/Fz0eSWFsmYmkpAe+uaupXyh3EzTaqy9imTsZcsnM4iaZFq76HS1nVhcLeHQ5T2rX
OCdoCkBR8DbMbZIeWygrYbagt9mMX6gmUg0GdGuUvKUe9NwuUaE5KysW0pGwcBmMYRkkwdu4Az17
t+ZIjDSTselhuynwWnoUgPurAUJKXhqmUgmB6OwOyrh+v6zBVgOx9cuhAjnIMMI8b6oIotJLwbAn
FJkW3C5beALuoGom41qceESjJ29Q+SbP19LjkeTZX3zz35V63atrN1c6irJwjpfrF4NzOqXH4ovw
IkFL5nn3sZVkiT0mKe3iAOtuLC2xX/ZOEzpwKZs/zv82Cs90P812l/I1i89wFavvj9VsDw0XPzw+
iBRmKOlmmoJsAFl8t/wH9/JXGACxrhU1hhX8P5hmEICYMe/KAONTiATQxQU/CD73R6KbQi3q59KE
UwZGUFhUhi1uf5SA0ZuJ2Esx/5lalZlehQQu/sVtq/OQYE/UaJKAZD+hVuygevmLLmxXeGrfPuRr
jfZhQJYlmmm1xMIB+val8s7VRYC/D+rgqnvebRMH6IGqY+p2izjY1EgXnJuZJ79gXNTIEDVhEB9c
OeuGnm9bphUeLwh28/1anBQPbU4l0PiiGK/YUyeTcSlsNloZcY3xAValww5Qerkn1IQSEwmLoDDs
TUdRsfWzOG2WaKB+d2zPLgpfCr4ppgrS4jLtco4RqNDjj8EV6WoG19gTBFWI9K99F/L/ZLVaGw08
DBwRaPuOl22WIuqfTpwC0/IsGFRislv8vSafPp6Tq6t3tqJgLBp366pI4EHdjXt5yzVf+TWQzkRm
bUgNwRTvKAwH88a9wbu6fGLErNVzrBYViaqRl5orHMVgDJDY9wrk0VqcwIUT3fl0Tgfcf8EKf29k
RNBykCHz4HzcjtwtRfA2/VSMpt/Kla/7k0lnJfOrwunZkyRnOEvWhiTnv1eqqxx6WZuIRHPtgaUk
jW6TVnTBs4blOOdPRku4xfraJVL5OAl/j3n1w3yRccW3K1WqHGDzyme8gOzlNsy1AauRE1RS/4oh
Hy+x21Mx0gu2FGJ9vhoqnhUg5wrMmM7nwIfiLwEJyhkLbvADQBlFtCAPckKKEXuLWWHvxpAYTVJ4
0dSM5LlLW0aCSXNn2VXH5wFVt3aGjHRnALj7f0SusTr3812a0u9K9DK5Zph3ZNQ7uxgywOPbNfSm
RUc0PaXYSO7jyyRXgcwCFrMzjx/mcuj+9l4NJnxxjHXSTzvZI4Ptkb7AK8X/YmLNnPHJ6VWvPwYO
IVvWmC1MSM6djVoT3QFV1GfyvfNHcyo0Gt0wsC45AU0/bQsKD3BAdUM/JCYcJn48VSTRuTcskPEo
El9sqZr/sdHpIUGtfDl8dk5Fk5BhxmBBuJX95Nv6A00lL18c/OFsIx9hXJl8z/mxBhk+nGicAeBs
2TlQ892yf0nN8RtSGG5nI1VfpsxtvboA2EIf5FH7/N+SOQYodfqohFPy3/NncQ7jstYcxHGWY2lR
FTLHXKMFOJP09W9e6DzeW8MGnjX2mNSDsXskdnBCUPG1ECH2wiA1mJDyvH8ns0N9zMtur0JpQ8Rz
rb3CgKPGtWKbcElZETaLvBD1K2tYvApSUudj4diPQmmrb/jb/g5X0k38L399SPlF0cg8iwvrc/7E
tLoS+9s3S8fXzWZXfhmQyqdjtxPShqitERmpESglZWIg3h83k4nJqcuSQ8i84VhLs9dukd5Mz1xt
5A9H/9JF7Tp+QtKSNoVvQp/sSt1sUq6pQO6oEqviKz7yQLdVEY/guYhOG8o7+lCSrdvZ9r6U6w55
w+kDp0qaHM1gijCK0VIX9pejvaoxr1d6vceUvtyP8LBWfG+l3a52aTtFjP/IfpRBI9uxdUpDzXL3
YTubWaPxuB1FVApZtiAB/TA8s/R7Wc2aEKWbjTjRzVdzsqKRyo0nTVisZLlkBaFI4XwYEOI+U2uQ
3Q6gknHmD58jato4U1YHcVGRewfmrjXRZvhi9NLdcp8itemk+17ln5zYobahZqlPI1apnpQKBYbR
eiyQFYvp5o8znl2fHlmkWezD5nGyRGmw9H5dVJ+Dwcs9rl37pLJ70W780VxgaX9YqmCK+rKk405K
lXznMQhmtZcdRRr++wWNraPaMcntv2STZYl6JeGj1ZOwARy0cpCpkOH3D690taqOqBvUieulPLCz
GE31filMhvGgoVdcsMwcQVomBBHr84RGNsiOSIpkKfDP2fp3ud9XoQT12kaI6jJEeKxAL7VCYZti
vRwPjv4SoVgqzC/o4OoWj2Knt4Zte1T/SHx5g4uDAj+pV/rfareibrD7+RK9F8yQd8sYjGZKdp9O
NqRlLLQ982J9Fi+IJCpfjb/scoydkubTr9RzLZW3kWdqC5dbwWYUwejjfZh/uKkG+AJJxku7lLzZ
k9wX5gwqFzzZ9dycTi2ZrkGkE3VxF1l/fZIt1Rr5Rp5XqJF61jL2JxgXqcZdz7iXAP+PKeIwNXAc
3102q7oELJewYDF4Z7muHnFnQNR6pPz+fcGl9vkIBLc7gwsZVH/yaTjPaY94PzUE7AZNNfZUL5eo
KZY4VIlLQPTBZ7WlEsVIA6ypfe5ecE7wory85sP1cMxlfUhyKFcYw522ZZNxxG2kQoGGxS5MyBaB
Eo7eQJoAOlT/Kc5M2576laVRKMaF/tEk24aYxtg1ormlbLK02i/MnWW1gZ4MzjcDaMgyN99YW45+
beeQAhISejqWX/ptX3Bw3fWGHrs9JEzLpky9Kvxvk2LeyJtd+WbcwUleFIl3fVCZkhvxw0B8Dq+v
+IombMemG+5F2ZUuYFNhwhxIpysMuaQd+rAmALwhG/uaOJS1LGimkcFKuNr6dqj32zU8P5Yq99Ht
y1riqfqKwHlPPA4tXXaLGuLBfdu0ZKJ5udAYTRnsNr93OIUSh0GYFU5WrcfsVik7cuxk1uE6feSb
V6+yG73gMACqErsohGS59ezKoPRNh1AH+mTHkt31qC+wnOC5b4AQCAv0LWp9pY0CqL6wEZTVCxsQ
R1Ux0dfzKXvhzCZpRybAgDCYH867I1dLX+chjVPbyJC75S9p3o0/2iRB9FnN0EV6w1C8mT5Ir6h6
u4Rz7qYChTxef1bjomYs8qI9b+Mgu/5zcUyf5f3yB+gAPCqRuW8UIrxuWceQkdqvqjIlU8XYqT5K
Sh/ahMYUVd0URmb6Ut0r1t3RW25DvjTAVU5ivFssZ08ofglpttm8caknyCL9fH9VaFcgz8KmBqI6
USQ2eADNU+8xu7nl/MWiES9mR0Q0y2qyI44l6vZGblqsd7Om7x6j+5giNmZ149l+enhF4kAdr6vE
Fslz5sex//UUhvCcaamdxw1hGmaVeSeHDq3bZPBYGlYNPAkcR0EY1QZFl+HCNLy2sAbUFM83IYQE
5bd75tuD2WQMa2zsuJhz40hkBwvE92Nw22y37LPpSueh2nWt73py80Q5VyAHJq5c5OPITSkMVBfU
YRj8ew9Nm/ZIBuGex9fa+4tYWATdfv/U6Xc16KIsC8tX2EM+ZruYSdaQPzxp8mT2CWuryGq3vcm2
bP3MZ4OWjleAySlBPst9SR2ImBdJkcLFw/4qi/SIM74DpaTjrg7VYkN6Y0dsNxg3Ne+NJfxVBR1R
z1cT7LHBZO4Q4/MBWTHh58UekMo5JDoogHoihiKy43BkrN+s7h1bfAbOqoSOsRZx4WZq6JTs+OqL
VqlIPDQcjlfM9PoCCyupnkxjJWXAIiY/Lpt7XT/lsePuPcCVsl1SKxJGqnxqjUxYV+L5RNSOH3Iq
n9UsUUYD7BrMA1HeclSOF92NrQ0VnKKYQ2+BGSu+MirMB1f9AEYYorn0j8dvN5hkwH7nlAs7FNZ/
U6bl7yJPyBUAAryjLXeTkM4lWfiXJRoITEbeVUwvE7AsYR2NgZrWYABFSKESL4Ss1eIInaB+7POg
rpnYf4V2ZKIBUWtmW9/ikF2Fa/bmZZ+AepTNkPEkqyYN+DSZxsZMFzeTCJL9U+568pQaKEaSNnS/
3Dd+Lx+48d4Ih4xuZNPh3DP9Jg3awMlIeZR/BEifufXQZ/fTW4aPluWwRlUBBQtDqWKvl6WNVex5
z9/IFeCAc9A823N4RNTONoIqP6tKCW/EaS3XkIftVCiL5dbPr6HWSWPd2BdZTY9f1HZfjKKSzgZ6
j1XR3+yauEh+taQOsm60HN8ryE1LhDA8XVzfizC4gZhybPB8RECkGilKIYWNPDbHAsLiEfOziNqy
jRkzUoURrRnLeHKdUrEE/m7JcHyHgkfrjQ+gYMN+siWmnDBJxs0ZUVtY/mDkGNjm741JUYtJLh6b
EqKXuIZ1Cq3ZOqrJZnMLYl3OwfzXkBM6Dqwq1SF5xILwvwqHFccSIvQ7dqly8dXPJusqVtv7Lvjt
HaCSmWKfmHxr4F+zML7ZGoWzgVTzi0RDSoEV38EUtIcIZ1QfuloZkpl0K3QNB090SFzOmKtGXdPO
ajhajK+7bbFDg2R+U3g+eMM51uF2MgG1c7D0YYSxL7KGjAe3bhesOnZPWkzF4XLcW7sIhm8GglpP
sBGUN1D0/AI6jmVmsLA0IjE9m4GIcMPa6uxoefLi1CwQubDIJdWAC/WOdNCugaXFhO8vHvMYMe/F
/NHpYEa4xf2hlEQ3vHjX/99Z4nqzze6QBdWjRNuGuZB0OfJlfZnaoZsFBTJ8bC2vkWzWLYEJLSEX
T+wHnR5PFKvcZdNqhgBEZ3LHIJw0vhoqt1IeYtICcJMLl8ln79EDLLge/C0I021f0LX4G7M9XgzC
lkHj35xsUYjzhYsOLQEGMO6cvhlIe92jJWRv91K7ncutn1ZNz/whd+8MT60+T1Z8VfdBSy9dYTuL
UPmuITbZiLTm5WpvChciAADzP7+WunMQ18hke2K0LktkP/Gu0zKJnE2XeovJAn9Tohkrurvkhk5T
ryGQZ5DBnlJuAGBVkIqGqfvVc7hRFU7fcLHF9C5Wf1qbsMvmdFwqW2NqoD+JkZ0UXx3WWeBCMV/u
C0CVqAm6dHYQjgKDSaD1lii+XhldX0awT4db+0uIEvleDuZJbNQIuBLw8Spn3l6yzozA41SB7IaD
ueAg9mkqdEdk+5IqzRzi4ja/9lNk6g/e/CMpdqzoMJYHpexVJQowpjNKbVMw7yNBpkQkKvbVELGU
2pNNuaOGDw7dZEUoyYuBGO1Jp2FbHVrjbcJubiHco9efUJ+Qod77ZUHB6m45cy4qTnpxvXxaGLiw
B8bQPLVB8XkRzN6BoLGgzXgHwReN1RsxSbI1Oz4Cqb6NXUX/NOXKi9TdUa3MzlTEY1siQCkk+QpW
aMAgKPj+Tc4pV9G9qkSPavvfzTBsTsXjp1AR+bIHiag2Je5mpy2R4jPshGi4xm0CQ+qvwMVBao9i
B77iNOHMAs3gSdLnAQu504z5K17GT/ci/a/ukDcR7SUd77CIx7bNp7ksRBduwBB6aZ87SyDQSOp+
nu3bE8b998zL24JRzZUhfTKJA91BKQCGkR3jNrjF8Vmi+J5QncnzPkuGNmtUJVPtDzgEHgq1Dp6I
AJ9wx6fsO5Z72m2wjFxE2LLqHIL5qwNExDhCQ9mgLWwvmh6K+rgguiq0mekKoWWB1Q5YbccxH/mD
I2HUlvHvVsya28sXUmfnuEv8xFXoxDQ0UUIXTAZcNz3uOg74N6XilN1OfLq/ygmqyiOolIelJ0nl
+b+j49biuWN7REJsV2HV/bZxlCYKO5Epmi7/wFgAFRiNCPVNGd9ycHoO/ZLpcaiPfWuARYaI3x3a
c5ed5s0UFdZYNp/n9Yjyju6NdtmJvts8zGP2uZKu/Tk5wiszDfSFrfshnY9e0XMurRmz24zNP+MY
pmsyPfTdqQnQ1QNwG8HhAenStXhYLb2Cli29vA57VB3dzfaT5yGM7aiQ5LUTtp9JZHK6rj/PVWl/
b+O+yUlbCePYKaPsToExHKgi/1oiI78BcotRQQtbVs/lTCcQCN01/lsnB1ALho0WG5Vu5Z+oinAO
xLYrhpxUrnw5/tIcD1Mdxd3+1orQWIG8Panhjgl0enII7KsctUoa5f0GoTcWxg8YFHXip1Byw1pl
NwB9ESHxCZaF5+VlgUJjj+24A0JulXuitopVmU1NYWcodVInyDPq6eX9P/LWyQsamTyFlbyId7pZ
2Qv2upP+xwO7HkasPnhesYLeiL536fklU+uGu2KpTjMAWuYqtV9whF02dB5DBNobdHZmolkCWYQ4
500hvpksgGfganz4TF3Rfh6D62lvmX3+7ZGpCHNg1253AGToUJewMRkBIymlQDDfX7fTY3RguaMN
BPu6bUCUdLYZidBSCKwwwUIY2BpvGD+hmSlzhwPTbbY/n6bRtxoVWYeAdmbbXhWy38Oxe67nUoTG
2SQbHur44A5J0foI0ugwD2LT1muC4MpBCSv+6pG4643Pla2P9fThfCV4+t1D7Vsho1raR7jTiGI0
lXrGX9+8iV8inOWoF6N9qqjNiuLsvnANS7c9rm8V9F3KruQFQZ9j7HzW4N2eUYGO6P2W5FNEJDyQ
JtvIM84g0OiqSg73h9ZSEv5aM9mUHPaBoAlBbzgtXNO5vk4kvxMRMUTwi5Wn+jhUNyQODL/UIf0T
Fw04XWZ7upXXSQzsIH4b0XbTLNM5/5jcEJh2B0NsEGig+bv/4JW28rLco3SoaExMmwbIQVvG5mWM
5/jQMfPwFGO9UxC+l8u5ttRK8ZwAbIvzDLKCGZrNPFsi+2L/jlRMc9QaiQZwNkSUtOgakf7dOPns
uajcgWUJToz6AQ7XMUHl8K6+zGkSE9F6U8ctZ90IXjbVS0ztayJ1OAj67vF60GJcoyK5XFoR08bX
dE7IQPJ98Lj8l9Z1tVGaQ7SnEP381BqTTxESYeBBf/5CbL86xA2F2k1HqRZbQm0EXHQo1K3zjJG1
ucptpTW849tT97RpsnixpXLc/BsDUvYxm5uWYOpNzqTqB9qXhY/tgv5leIJV/pzkpMSQDMhLH+cf
xDhg5OIXCdCSFaBuuWigMrPpVYv4kvu0IXYZSj2V/JUeoAC5hj4IA3fqt3oyhnp3auTXikYKUzoO
r1dasPTBAqdXrbxKfn2X+Hg7P/eIF7jdX8zZdlCy4T7G+wpVZTqe2u4CTLwHE0UTLY2uv6bYCSTM
3YNdTBkA3kea/3GyPezH/TjsP0kCFpZjgkXfWXkgd8AhLkH5jrel8+8yUM+/IMtDFWzFfXibpUGZ
JdlxcTYb2fn/v6cDQ71jLVDq7cnuFpARyJKIWGA7AXRUNdqISZy09AbQ+ebC6wWZvaIR3oDEt2vt
jIE/hLXbDSeEK/sOWqlgiBPT6NadURbHzVj6cPtrB1/Dlo/J1YwwsEdJOkBeJT7/JNsF8Grxsxrl
9Pbi6wWS1NYuHsv7D0cN7FF9m6u4m3UJwQGhYrGNvz3bVvsllWC/DldmXXwesr8fwuBmqaKKb/a8
tZe1P9w36VjOog5tKMZDNsJvVomYIF6ULn+BIqGTk5NZ+7RpVF/dHo0bvHTAh3zuUaF3KsiCviJo
UlYxwQ+cUDiVtDcha8ULQH9ZDLuCsnUNVUC3yeAcXLBZZRZjWoOIF6pCpeB7fyw3BpgrAINZi1jJ
OjB0jrIBKu7Cz4Q9T0um/WSqEqsdHpWmt99lC4hz5sA+ZB028EEdEIFp7uUh9GeEtuxvyEUMy3hP
aFaj3nLGf6Vm5gcV9JR6GB0gb7D+Ma13DoCrpJc6FmTU22P7ZrTmgMCd7nCwXekwaQflA8aXPj8Q
iyKEYvwc/DEdaYhal+AZF3Wyyf8ESN5JEgMONVreojK2cSYEvOnWIxXJ5xDpXCTTGKbpfr3RyCBO
AQ7ZAWN4RLj5E7tzJtK9b8jdUyLcYGXuuvxcdSYEDWFFZaHKOx1adNnjDf7SKuEKq+l0EDanx9tV
vVtxtTizzCBdrVDKQPrnYKTbGpa05r+FMVKpzVKtgCsp45Lyn8qmFAtPjALs+EPc5Xi3rpzo86Ak
vsDZhxSa1PHP2+AhwWFpTnXZu5LH2tL06qdhnJDzPbkxKHVM39NncfaaWu6AbVHvsd7Z8IJWboy8
7EUVmKh4f7nz84U3BsPBWyhl7x94quGfxDmGPD7liFUipgQ8q0fiK3jzckEXd5zq7Q7SfkpX9Dow
ciUHYHt5tF0tKYLJVfc7OZN6da3GPWKnrAO24WRLXTpGjEL57o0GSvh/P7zohDWP34F/Bm7PC5nH
xM3tMoLgcJyU7c26FHctMwt0iFchcp8GFlwKbnDYvTVtfYv2AxmC0+Hlu1c3ouUYO0GPJyCCgn+g
xcCRcyyJuXn+KRmuUXagrPome2K2C2BBCHCoBYFvlVhASL/ngKURUyVERU9Eel/d9eXQk3E9oHzS
xaQb+Y6kTUsbtvVzNytyySSOuPmd/xRdumJsRwPEcfoJPLGn2g0TVJVl12+6uwdHrAt8eWryt28i
AYFuxvNci57GBITzz46bgnUj8WcTUD10UX/DGJZ0uHqUpopm98q/CkF4nRODNObl53ySqp72QWKG
FFSaKCB48jvwl0eM6hR6f0dKIY9QX0FL9iuKR1wY8XRSyqS+XsA4suu/dlMTSXyKGvascmmEVpu3
90Ivfqr2WtlSiIsVPFyoRBpxSQ7nw9GBVUpEn6MyRSLEy4+DHxtuVvKsF9hOj6eutNh3hfbogOvp
q9HDg6cYvC9qQwfUZRv+cFhLRIMtuOOkspwCBGEj8PsDdwl9dUnuUxVmiz9bAFMxwx/kHztps+BG
4Vnd/jDZLewjkJaR4jPTK7iDcB6VGwcuVp7OhMiSz/MWJOe5Rz7vkgZtm8T4UyygiLDaL+BklLju
rfime9/VqVewBprPRxbEJ3wTopFhAmTi0VoQjFXTLZeF3zLIymuPvMZ/b9+2qbIg+jQdN+FCTZyl
jPgS6+GzdqMof7pkRdw5rQ9Z90H8zMF9nqlZcjngv3OvSp6hIS5Mjp9Iro1QK8SGm4KzeYM/hp3E
iElkUKkCJFoeiW+siDXDdcCy/betqdJpST87ohRJ0bFEBecfXLMoUDLD2WnG3dexxO58/tG4A9o3
XRmT5RJqDjeKLiZfp5JRVYgST0asvkc14lXVGkOlEKSnOTG+OWAqt3YOJMVhGMxLnNVi0z5gKj43
HYzjCwCuxWvhNWZlUl7aNQDaCJ3cKePQhD7kLgmHyGr8bGpvtWSgiDM8UD/uJScN8vCqf70UaCYJ
eRq3XsdgT3c6mUBrR8JtIujZQWQNZgZTrCpOqRqkRz1sSOSb8BAzGz9hzpIujoBu+v4xR9tKb1x8
XCFZcIkxVEFpVJycb2iMo6c5i5M7s8m4omffJzaL0aYCpVI3gXDiS9cD5L2bczg6+yb5i+wqJkY2
crNUU6X1fSQdCvCkF/Fosjg9b4inzx5KV2cWZrpwSbvxJopiQwIl2OdhwV1qHi/wCezSCUY/BvU7
+weuUY4uccfcRWBajNSn5T9KPyMUAw7M5eAU/nVsBKkV5TiHNfxNhGE/UHD2YDo7ew4EngyiiYFv
Bw6fQ3pOKc6aiJE4BMmUe0DsTcN7ck1vFf9vguJfoNLUOoHZfUh9/hECMvkhtBcmbt3zLAdGQKwj
gJZN1EEGSMq1k/RdPw3M4XaXq/xRCJ99lCvuFCBDq/EMNL9WaOvkKzsBl41RH1j0WUbZptBLFSEH
C0XwjLqE2M1ywA2P+K5SU1DQ6Vjo+7Ovl54nT5IBACQTh572agA4/aeTTekFC+6HIn770ZhB8yCh
efrU/CdwrYj1TwnhqeDFnKmajtaJilc2qeVXtX8YNtEs2ryUtQSBbTgCtqo4kvjMS6JqY6kIIFzp
BkCuHQN5UqKDTU1RS4jgW87TpUj0kSsD6Chq0vd22Msk5TtXWYP+hybDbHWx1PgQXM2c2c8muNSs
8izMnTE7Lz9CzvLCUlKxRFo9YfT6HvyXq1JTa7WI3Sms8auNUbzDN5C2gZEmYc8gUBKAklX8/f1W
XevfSdM6bv0Cg1p0lrc4q2FtGav+Z+TKfYJQdAKAw9lDJnnvp4wSpg0544/Dt9OjG/3KSC6DSyNR
WQDzFx7/96d5KNZfgW5CvJJmCPtcGeZzs2L57rxcrutgpiFFTo7KL9FKojgtYcXkUDAdWeNDoVO6
8mztRIp7uUAKvQRKGSxbNATHE2gizscirUOXBmcpmFWK4rubNuj1jPPXeUB94kmV9B3bWN8Pz91B
ARjbCimphubMsyvljdAP/OLzKx2FlRzMGhTNjgS/eVwAwcUnPB/YITpTIx+NOf/wGovRG2HLycKo
aNux00yrEJu9pDx3t34BqIx+Rl0Dx8V0g2d2iBoQ9Vs/WVWD6DivqBGlmwJMW8obkjlrWzjXdSdf
cNqH/cykmPkk1niLM3mrFfxJ9/0bbQQm7BdOcdUiiEJ7qAlm1IfOelf92ByUA8FK4XRvhY//H5Vb
V+W1faLcAER+D+LnBBrfHUExznUWn9nINspqxBQ8Cz4lIW5WjPILhTtVU5U2XXAs3CqrtDfAcbRf
GTcwVw+c+9yO0QZFNkLbllb38sl8bLcZWKarL7DB+AJ2+0C8q+09Li6nI3uaU/oGbZg0N8VXOB/y
lPkDDnTYqcyCeSxzUChFZgmMB6HpxAeu2B4+pqGs6S4leCWuOBLl11MrlHUlgw0Qu7nWQMbA895K
cjIGQaD4pQQm/jXAPkA5mDOuZy+UJ2A0T0zNlRHPMqMyLVv+W6ZqPqvMLKxqk37GS/Osd4rIEhNE
MiUOHhjAni6G5tuTvqedxceI2AG4+WrsBLAf1N07E73TAm9vs+jsOFuDf5EQ5/yaXAWoYbO5XTDI
DywZPiamDpGp+nI7u1OdFeXpGQlCU4flZfE6nCsZ/YezpP/nwTMSsEaZoziVvEOdp0sAhT4rES+7
lCoB5L6CF9BTzP/d9nk6/NuwYZmoXGDSU+BOPMMnxUkMHMiLjlooOd00PZqfZxYDkWiYbsZGBXa3
pPY2m+ocnR0bifwRUNgWSExbRsQh7RVKcUpzt3uSv61OCxqSM0k3DXhXAlAdTxcRxG1mF0KQX3iy
/t+Z+J4+1I1B9+HKIblzpND5zD6HKb2jeqcmrr1F6KGwCB+5I3IeyK9UparGGb3TCru8sxWzTxQ+
uzSjUnHRdY4L0/wynw/45xx0q35F+jJE3a0/QNOM2ERybPTnqEKmFcrss7s12CqaiG7maSl+FtLe
OKk9QxcUdPSez9zdTsYpwGm5tByWU0FF4hZ7GJLkMFSXbEap/r80MB+ei+BsjPZnbPUpC9Xv8EjP
nzY9cjgLuDvxpJnyY+e4YQAM6qMJ64ucPTgLMFz4lTPcAzmH9RYhAft4sGnsWqpxnRrzoDFHy8cu
PuBDFUGCdxPHRd9Jf4c+NOHDAKYb/H7bfKTRRwdBOixopzljIiWSSepdCg7+fX2/oqojptjv4K41
2wGW/Jt37JZhUbcN1XILRsOhoDNInSSH3urkJIagtPJg4dM6Nbm9m6qdaODMiDFflB7NWrbptlOm
dax8pJXUuk6KetNhd/XyWwptMBzChtjezWzkjEQ5nQBTZi74/dZmNTTToi4E26uBMi4dSLob/n3j
JPByTA7v8nh4c6gUP05aK4a8ig2ONrnO5PLeG7nxF+asJeGYr3NezPOFhDlk75V0xFqEASueoRGI
RO1Sy4Afiu8tT0yJrVNAgDWAIHUU6AInkyFw/B8QS/uSB/GdL2pReXz6MBI/90V/zk/3zR3Gzxd9
OmBGIXbRif7XZ+NyorvIs+ZjG5STetn7ppsZzoX/8LJFfrjONZmKsd9AL4ojwQdmEJ/DIyakKshn
d39cC93I9aZTg2jHdSsnROkgxOTX6xmhXQQlEuYI3WF3cFj+1jOu3R15XsvXK4HNE+ZQiuatmZDX
3R39LvorKI+Uv/xyFEWCQK1ZYJ704xG4ftVpXpyNwgnlcwq2fSX3jc28mK2RR/XUet1soAuY7uqK
3KWmQ9TjK5zWRbIx02KGoiE0TOnEr6VdwJYMa2N3UQmK6Nkw99CSCP9oAwgYRZw/51QeCeS5QwW/
pg2gY0lcbjOcYEkz5be3sZ2eephwDTCv6mjMcc6T401I+7yHBOBRRbZqRU0RLa6rJdOeGPPKOfKU
qpLj2BUsrtial9YEb1fFC412ZIkp+4j8a5vqVxwrhrozXIEkTmdwp1EqPmk1Fppf9DlAmCDyiMOt
/kjYIuKJsCu/9B+0WDWqxcuw5Fs4tn+S/72cHFU+canEnCnGb3LktxyVNYQtTWvSfGKSApG/DcKq
P2RHDXd6ViRQCiQi5qgzLJ/nM0erLq2Wa9N4CgTuWRo5/TezOlchtNJh3+8IF8S7eLHtp/cfYhFN
Hm6toqF8rqZ7++ZH/HYGmZ6jp6kyvC4QJK2dVmqNovK9Ab7nZjqW/TNbe4/oEzh0L82e3MVPSanr
FWq0lWTtqKJhv0p46HDVDt+PHvIqRJvflUmfnX2+D/M0aTQDRRDQOeCuLwDwV60m8zsw6CTXc9IH
J/+erd0a661HG+xzrZBtkUIl6RC/YsyuEdeq6+QjqN0mHi3v6GYqZAk7YOw0f8Ewjrp5oCQ6qoLn
ehSjATOxPcJjXeyDnyh3LsS+h3GzXio7wkgUM45fUKNvyWBMEOLh4be8iIq7iwfJn3wgPhFH/G1Q
6xU+9QTdsWRReTo70kwX3ATmv422Z4QnyQakCcA0+6dmq712yNGlx/741SgcfT4HDrD1lJH+WP3A
Awt6E8A3TlQ6r2bTiIt6kGo3DTSjTPOjoh6n2ZM8+i3lf67KGuh3uA/c5jSlH2x6xRfnoIvb7q+F
Ozvh5CHK5kuOp9Bj2kYu1m+BBxoDkmYRLXp/XT7OZ5QgU050vV4anKhDVwxLZnbhCbHQ5UVHoW/4
owpOSu4p+N9VEbiU6PuKGSq3hn4JjfAgwhsrvaRpgnwGexLa6Wy3pXkukg3sOROpvMrCTOMqsF7g
w70Ss8gE96G4b/StQ+azXMlZF/yGoPSJXIyTZZBc20VjIbB71jjYLIg4uApGbqiIV3etGdcPvUwI
oEZ4SEtdn4l1whOxX6HPMJFvUyI/ExQeM4stGXmRHF3eo+HZX3AM5a3tROpfKuLY8o99w8DU7G/3
YS2nxVah0FHBmin0CQg2jCJSNkNJ3r5r34VMiQ+ho5zwONj12TOwUazH/idetV7bQdllAB6a8DoO
D0KcAsXwpiPb5Nfjb6jHtwI//Oo/r7ZIPE30Wyz0qI4/3M6xf3EwVCdRoRHkrFeEJtw7hFHRroxI
AWRpgopIZB7Yrvsp+Uq4PQ+GVq+pqSmuvCx7gXjrxbW5dP3l264zIfYu6OpQNTppmeKJ8FsQmThc
n4RrnBVXtX4+9hsH5fqu7fMR1svopSrurtGZdT6ZQJxvP8YVHnB4fbABHrfL32j95Ek7WPacWBAJ
e7HehD+yaSaNCErcTpqQoKLCvQVoRxEsuBefM/O89d0299sLl/LA2sVw43K1yvEvUSDlyltqejou
RPru4wMuWvUSZCQgw8L1UYxaj9vLCzWwZvy431zKXwjirJ1y3w/9EE5o5dc6myNse3vSXTjJgTaP
t0tV6ffRAGe7Bme9RLmXVhj1dnYj3L/t4BkasI2hDTzrPdxdaRbJi0N6CS7a/cuNC4KDYhOywGY2
xrii5uIPk4dSwX2j231YCOyKxRyE9LXAb1zTJUliBNa7E/AxACTBUbyGpEsZOerPo5t46REnvlcR
CjCaORQfbIve3ZNNTjaj3TyBqGJTkPFhWlR4z/Z1ojNKF/BJvVC6wxDyARbBbAe20Ffk0UScHizv
/bS1s16XUN2qDeGjO+29JaK+HH6DWMchkAVNzMca/rkdvl8wD1oryxxaKhM9XeN4MyKmv2+okbx/
KYUTQU2B6UvOBSSUqIJ/astbuD0KGfjE/S1sKOkmrLV+U1euZrvrx4QP/5vW1UDPQ7/AZ3lsE870
BgFXrtdBuNutzFB/R6nNm3JWIWWY8oaBZFSoSIzureykNO6ctinv5cBuHi9CwynmCCEjC8gVVXuH
RSoCFc23WhWeBcLHo459D91GxqD6X6/4IT4XajQwIRyhTS9LfY1iyTxcJvDizHOeccBHJwKNo39p
erfXt3vuXku/FMwVjklE15+F4fWyq5e+FbcWKEm7Bz7Sbo/2j/0Fj3jS4l8D7y5NII9snf+dgYp5
bxlue/RiuCMYqUbMgP+yFqRpWwPf0JR9/JbCHXitHL4g6J6ZcqVGKXZTqF4/2M5IYFdxQ6H0UDNT
Md4Hzf9/zXhYoqmFXAcpxs0Dgphb6EA2CoePs6L23A6OHBiNtBPVyvky5wqFK3Phl4o1ZILyBR7M
XRze/4ikGIG77P125KuvYP0A7fMJ7qvRsdXuaYVpD3l0sssCjEfTr73YhdzT3VPl72OHoAkAeNMk
kbB7fpouSAQ/jwP1zd2nSCfGhgC+DNF+cWUdH+gZ0w1vhIH6HJDwLW/+fsMJ8HyHHGC3+mdiknck
ySj/6wPWcJC0Zz61QlHsc6w3GkP7V/I+E8A+4liI/A1QuPh21XGfMTXfDCyvZvdiDsVh0GTDQtB5
C+ORhXKpLpVOQiROeZjJNXVEaK6pjhn3QAqOWZ4AGpBiQUIXT7gBiO4GTbxkXizhAtJ34xdcj+fS
3GJfkgO5Cp9Jnx9uDYa+4RwoDdKZoFtp+xp/Dsx/WuLNBB65g2rniYbuOdCLQwJHFuUnINkjKTJh
oahFSzG4z1RK9nzW6mPg1F+QXDz+Ao9VZCl4LAeWV/6+JvB8fEFqaxgOxRzclSzN/UDIoxJjzzqG
NfxuWamqhYFN69H/ZbwX1lqtoC/hB5rqRz7iSX6Boswh0XA2ZBg4YBmYlGG2C7+6VwHy6l+rFBxL
7lsTdTDgrJ+zbZiZUx/pT/VL6tfu6V7OmEzw/7EdoDjF9HsyRucT3QvxOoogT6oU+td00RvgnqVf
1efEF+HFEmpJ9kTnWzV+C0yj0pczu7Kz9vefvXk3Zewwksg8tOilmm7f9iQpy3kbhTn7LN5D2SJL
o4alF4oDo2kCxkv6cf+pRMn4t5DNur53swp7Diyss698WwM4XdFeSz1QyuuRr6LwVqr1Urxy7ufU
NVyDc9OmRFW1djZoz1BCLIftsINF54yx2O8eFBvQ8/q0okcpAm5Ys7fBD5jaabiEDUWB3hxmr/4S
rsTQPo2DiZBjmzXPvgjL2MHU6x/Hmz3pnYK0mzTBwkwBWyCbL5WRzVGoo4SNq8XyficbwX3zDJvr
4i7/TkCKXYHTOu5DaEQHjujn6eaN1YD35zc5NIxv+7mqLMEz0FasYAlTqwQ49yTPfcWMjr3yOIp+
W6D3YTesw0gb2U1LethbK3shx4lIoWW2ptx2BbB8y9w6Ba6jHsPrshrkFlBOn9Lsq8ByV8MuRP0O
xRiJ+AczLSh4TVE8l9giKeOz6B+vLYOvfXZhJXtoOgMlPf84tnASAHYYEXfDb9IVb+gMVZRT7tHm
Ex6fdBNwmXXsJC7eI8GriXkHDxyzWrQHM21dkyw0m9evtVagIYB6h6nyxFOkFIRgSAgDNFQ4q3AJ
CzqK2pFAVnbfZGMzG50TJRcvUvSmP8gAlVYHuVpdkuzZEwLZGZ8dA8V85dEZms09gO5e6yxDEO+b
uA6ym1k3Dj0BimFp3sNuwHdpxai4GJWjr9Js12FxYmUXghgd15bvPV3Hyvo7UtrDrO5KhoIYdq5u
T1R1GqFqcbDUk56VVOBE7SSyqzDcAwYFysPlfHWpSsynash4MISJb6IHNVytMoA7WFU1+aXl6AWT
XHTNPxQcPfoUnnauozR8K37UaYeTPxudHrYBfkbOZsaspZGhOLdoAE8u7nsZxLrvcWqqq8VQfNOI
84bUuLmHOj0+pe1d/HtKnd3h7Lnd61n9kvip5LuS+DtndZSRbID5+tghMgJPvN69RgRL8EnEjqts
CSP3mVjfakufZIt1BBw55bXkcHgWTBJpa4h5ywnLVqwqWEy5o7Hadz3a44hl8fyb4IhjoMHRVDdN
Os7HhaHyYxEL1e+VbHkByVsJRr82go0KtmApaNrU+yg0FMBAfKhURCTi7b/IhCE1RmZYvMf77OVo
PPc5ys1s4vyRsCGcBDVce0eYoFOo1zJHE+7Yu9NPpj6JFXMF6lXudNMwRUR5cX3K2Hvzv6avrpCK
XK+7EZjIuiYgTs8WCZBb6VgFEH/VVjfKQrx7lRMmr+crWhxb+oPMunZsQSeuE3G6rYQGMlQVrzQE
oG9vJcEYaw1FZ1mTfs5tF4wu67tC3UHP0O2tbg371fiPF4RMTsnNnVi/7J2Rz9J/eeKyYg1hc95Y
APG4vLZrKELpx1wQplsmxu1yrHSFI+ZtOm0i7DMnNnUzOAhfy8CgcT6edJhhEUoMSCU33IktKsBD
lJAfL4UhR0ZJ/AQZ6NVr5iwqMGnLdekLgN2axEYVZkBpCit4OVpxy8rr9PzDw/zv7KL2StfSePv7
MzuxauO36bEPHfNDu4gfYPYPwk2Vj3ZOn/gN8wGpTg7Qr3g1QAte9MThkRrM2AFkHQT5Mlggtg0U
w29Nf+Dkg1WPLXE8mgUePupYp2sDg+v3cBhrFU5ISzziMXSIJni+azfT4FsQX7/LcVrG10ukts9S
PQbDvg/E4Kcy6Gi6vT7UGgRRydagDFBJ23Cwuj6zlJAwra+g/gB4UHtQIzIH/17KTxtLIHqKkGDO
4njrKsFyYXkhpVLymHv3HtcpucdUkMk0HXfmRw5e1C8pTaOWyons5tryTvbMi+GO1PRZXvb/lUbC
pmlJKJU7FIWMcyMJoYUWCPPrFLFbH7/wGLYQ8dgfyA7fZmybHGawJotGa0chMEm2Uns+k5OQhulg
6zOoWmgX1RGCamUV4oLHiYGgSeYMbH/BaDAPett5ZbBE5CgsKGXWMzBPBODwUdC4jc+jq0uMJ4kC
nexpK3CunspnL4eUOuxCFXqq17M6NAP5lnGT3mSjM7JLxtVnWSWeyP42aj1Z04dRxGkpgPeExWRl
dkx2n46VE3xvoau3r8ukl28xwxQZudxzU10wjGcSCSftasTYbVgdASups5WpflLv9KioGC7Kcm9Y
54Gq23QeHmNsE6NZLu6jc82MEa3DF8SV1/Cz8NqPQBAklYtXwIHc9WWyFlG8MW97knXJwX8yf3G7
8tdtIgPKV7l5RoB0S50Kap+jzh9hPa1pVbp+PJUXOtwWnTNwBU6PujfYs0v3GEdchUICYeLPe1W/
iJpUgPrj+Tqz6nepSC8wLdtAlnH4bT/b5IhxgZeIA3WSR54asASFj3ZjmHI4k+1qbl8ZddP3vPF4
XAi/vwiHoUePTMLeyKKd+PY6Y9ArOfLPLmehSmfFsZ8ldrr64opJVKej+RY1B/WDJullhXIY1M77
wobxQelwTy8geQogRgMrh6BsmnZbwmXoYJZG3yT87oBDnLOK3gq6XT5+PNQ+gFFiFBl5SQF0nGLa
CBTyq6C86sAsWTHlspkah120uqCmp/f/1AOhQG1pOa7s43LdiCYQzGrNQoyMbglE8btv/hJ2VZ0J
Ja2lG70bAqUCufmRHXTHXV9Q2CdMiPBW4JgsBPbZ8rBHYmGwIqelVKjzfYQ9tydVL1JoGkJ8rdv7
28yb6piolU06RgQaby0Qo4EHv+F2RzBsWJYuc/45iZO8mG2s5p4MnbiAcPBQi8B/tI/dF6kyqAKS
Hsgx6i36/JyYJzI+3LQCZJjQDu9FyFbLlJd+nminAyMQDXecWpBEaXrn5v0nzRkesrpYLleBN0fj
Qlrhd3uMvA5LBaZ9lL0PJYh8RfMYqYlZkidpAM0cip9y4ajKfcJPDg0M8+8Yh1HmyKYSH6xJVEhd
LfS1TRItQmMqXLuncH6RoF34183y1JI0UgG5007DlX+R5ql6t4rkG4y5nO8LbNl4XRnbhtGmMHAF
yeetWTjjl2oij3WWSm7SphpLnSaV9+AEXn6Oq/uqBdrb/X9lpQB9RwFe4lm/blVKhaps9g+K1hT4
nPRAO4V1yDeWbCgGOuhu7M+I6CLA33wrF1LCR1zzOPHCHFz7uDsP+wgf64gk0jISg9kWw1Xm6SK2
JfBt2ipplAt33Fi4W2kcTj8qdze+VJ1cMoRGNEfvaoCCEkQIUuMBptv7gIa7bSMLSoZlOYFyHIKd
TSn68Mup9LBHWxU3w586ReKvDqB9e+UREGn6uuZ7fHiH73w7SR5EUyQNlXRj2nSZlIqQLr7+r2eb
60MEEbnyY96aNYUHznlRCNQ8lFYHclx7Ug5kjLr+aJlePQbQTtUjOmKZtCv2O2tBChSrjHKkBOpI
ukQt0F6BBrY94bK4VJFnDiQNQ3LLuoPaJocqfnjcksR7di1bP3fw9MDPE0ZOXqR9zOwkS7mGHSGQ
CjeQVubVCaordjI3va1MAheDdWRfgnh+lXdh0XHArGVYhjUZ8vBISCJz8oDYfxhfezcHWth4gvs1
EQzys/4BkCynSu5NnC0WFU4vo8b5n+HscDN9NQGXKWR12ZZBeZUzZr0FBOtFRBQdBeTbyDcfExe+
1QZZGyf/JnbAqLuQhUsW0KThDRamnVn8khcXgstRWJNQujwgOxThUwO+T8cwNSNM7XChpuK3yypw
2xNZ5GUK5ji7F7awGtY++EZmej28f122v3nZtmx++w/cKIEQT+yEU7bkTE4BlqDVziyNOr6Kb8gc
zhB8p6mRBoFlsm+TPGe4sLYLAT8q9wSWf6No9yPJnI7o6jmq5+LB4xHZ0xAsO1xdmOcyTrnR7EPI
REuUvz6BoRTp5jlBRg6IxXVfQ2I8f88N5STjQHtsa0rpxPYOHUY83gzyxbikvlmLyagXhvvK04qQ
tUReXOYLpVivYXogYq3E/kHz2u06w3E2Xnzuh4rwqDuSP1oKT0ra7x1xv3tvdvjLsGwJ9jAPciT4
1f2M138O9AWm+ZxXYQuJ2ZF0DuWMwh5Ier/+Hvz0+X7c7aNipG3+Hu5Q/CCHLCWSsOUSA/fuqrnt
wdik+PVCV2a/IH2E7ZSbWDZ3/qcNy39XdWoxFvrFBFEhtLX6Iqx6Xr3RTv9f12cUBx9U6gWoFIcn
ETuiRrBPnNUthqGdiNK6eQ16E3ZOCcu6L/o+SM0iCvz4Dj217wdXNy0c2ovmW5cqy1Npb0tuC0/r
yJrnCBIH1Xf+IxgFl3McYex3IHRTzT8FBJKRcJ3E/TdCb9m2GWOVjHrZl7wM1pvXgjUUGa5UbMgc
X7XP/A0cahUqGsuq6QlDMcM5wXZT2YGBZRnf/n2SxBWBvZZnLkueO8sYMkQpZ4m89RkOSdQWWmPp
lkGEFX8KOHuSvQrNy30cewP4d9wb3FzJ4oT2xz3/Zc0Z+AzThI/1s2YxrTebsxM2IoO/EsTxZkbc
ZUROxnKp52XqVChT5dfTy/w0JvKWE+VXChy5xHrvZEOV21FSjemd5m2Zi8WXvkE0x6wGRVpXpHKa
Ks2DMLCUplHfWxE8mm5pC80n0/sO+j1YtAIIpP9LKzU32oxZdR/eE4IJZheF59ZuHBbfPp4k5mb0
nWQXpsW4NxCZgYFxLf7dxRqACI39AWowK5KDHLgaS4RmKIPsXYjl2WHP59ctqFMX1zgcx99GK4uR
y7lbfEKHW4ZHguxWntT1TJgsCackinDiO0MPKi8+IDfxgRuyE+kZ/xaLZsGqbM1UMRSWBSa/Wmao
uHY9F/8VH+0p+oGrvJ4L+EHeW7+3wdAbxIMkI/Jb2U4yOzDDEY+xBrrRE8UVMiT20XQ2lsNCYE5m
U/bq55PidGGEKxeawwPzw6MLBeoVrjDc4/CgKHGBpH6wd3QLyG8hszn7A5ETbC40Pb98bDpPaPHO
YVpN7XrQ7esFHuFS/Qm6mB1gx/j+Hac3sujMl2reKCmknbLTGo7Cv0Cxdu8OXU29RJCF50TCLlZW
j0P+sbR+gj8dFBtq34CuApkiRrIzmrcTCYBSA1mTn6yj7o09/6HHaZ8ZN9zec3QOpYui1QPOL08M
RotLwhofTv0eCn7m7wmNhEP1IzWfchTyd8brsmj/EUrL8jhs4//0VM/dBokzolpZHu7wdnafMTU+
06g74y4+H8bp9RS1BrbySPwhBQR1O+TScb3vyNKhGMNyeAqPzDjO9FwGEwB10vOYGHt7uHRgffvp
zDMLPyvAXuIZ+jsQJCzRGN/GUjWLUIAIaqKgTMG8blHubI1EMqa6U67whamx7hFmSExoKfwhUoVm
Idtp1MTRd4+rLYx2F/z176pw5fAjV8PxbVDYtwYPvFE1MrdDs+ykZHEmi07o0HXZYZnisiWJvJTH
CbExY3zL1LpCKOTDLo0UfOIaQXnOAZJvaLZBRKvOIPuX2CQVkuxjPiGNi3w4abyt/cZxFG1jBK3q
Cw+2Qpnl8LIHpQCEK+bbjBH6ewl/fGrk54XeanI6Rfp6Kbw5kpg8YpeulE35gi6mQSvUO06tOyEb
uE/unGOnNHpnW1S2T9Y2feZ8fTp2kXh6krqwK7nri13DfaX5YH2R4ANgThnqOl0ogddCrn/Fy+OS
wVKxhjYpM35txTIf4M0mMupgzkG/s3bCyBLH+BD+GQZRLO5PQEpITyHZhxwoDmHJ7oGPGxiIGr0H
cQ9BY+97eVlMqbaiXRyapPtk2w1fOQ0cVBPh3VMBfWdmtpCB5ggAYbeIo6MGisECaeRGe+25/SPb
Bywx3rkABbuIJJ4dwZJe1i8ay5LQ0tWoptRHxbrJGmIad8gFg3Gu4DKIY1kB6JAakyIfRNPAGmkS
XDXnhRP7JdSlkPkNV3KwWQjwsn1CQdrXVzjyesKnYMixlYeEcpSSrFxe3Row0ngxi0AOoceRmo3H
Rof0eis4vNcysvYP6U0CfNH4zNwqEa2JLEt8XN6YhGXHerQTPCtR+sZVVX8M7KGPthqKxdTHdwWX
z6F5azMeN4Xto++auM55iHk9nsLvkGl8m9WajISg2UYEr6YhJu+JuXSbU4GYHAMj15tPwTelZLV8
ByCtUIeRY1O9rWV2TQG9blTDuM9r9Z3nQExjhm4keGU/JT2t71U4iXW0E1+v9WiEODo6EF+QW3Uf
sfybKSG0lktMTmsPpxdmGTuoS9p/UxLmMEL7gMEnqbsgQDesNUxoaWcQdChLGCbgEbzy9JaaC4lK
81AzwrbNgqX01Y/gXSObfFZGWRnSRIa/wfIiPjrPQKYpzKGgoZwXzqrN5XdJxVw0+RPwro2g6yyU
0PiTfgynoxe0Cdgz6bglXBeHD3InxjvfVuWVKCQop1F2I1JHx5pCNOE1IMlrEAMMuIrDbn57cY5x
vNDBOeYfS5nGhR1fx602YQLA8ZAffXgeBRg9GkICnCbCcZg1NHx6/il+r7ClnEtJ82E970pVGqaD
sAatxF7z/WLxrwQRAQMnsfFXt6IpYenHIfhiqX7cDnccwiXIEwdZLzX0WUsJpRJ0JiEfoLdbrvBP
5sPjqUN1Vc+NdeC1S64ewpE+GMFP41EiK3SYX58/8WeWz3cos7MiQfw1DqU04K9HnhSE+kIPpx1m
U3pUf/o/QQ8QiwyGnkucXQgkpFngDD3eBAKKx7brDLHHRCoIQRc1o7/F49eAHdnTDO4rvt9ywbPc
QYN0PcqGLG2xJS4TnPJiX+izneb74l5Fu54Io698PQciRvzahoaj5D0ZjRaRCNgwWQHqkHhVo3iN
3KNhpCBh0rxL4WZ5cUc2IQm2xQsO23F390o0AZ+ySaHOV9G46EfG1ZH6zi8vKzSnxwJ3tV5Uf5Jd
QNnKktwTzYTo9uNCDdUownJ06uaB0bDKEZfWyYroLAjLqrwFsJJRnCsYp0RzHmT9V+akktWIil3C
X7jDkNZfFbZbVRrx0GydRsJivst5x8m1fgLZ14HOezI2Rk251Plbt4Hn8r5pJkZLL5nXBppqXLW2
xkvplTUP6psMmih/BbJvP/dIocIB8A/pJr6treSPQ9L2/shmINaHBCLDdqAVsEtFSzz59yRnZB4N
EL5ztNgekTPcVXzh66nXT4ARaxfcsRUXfwdfsFSyTJIRisI5BF0bdr/kqQgDibzy+c9pY0WAbmqH
pcjHMGjh4eiLHKfl97lB4PUJmuY89764aga9IIDUNct0zcfhfLXA9qQwAf3VN1pvNY8THdUO1bk4
1ygHSiIWi2i/SUKneVqyVg/B1g9k/EtJUY8Sdza0aXjUTRWuyojpa1u+TpOlwXHPa5ZV+P8oSCud
QCgzYHBvdNKefXSSbbkwa1vOPMAtgkl40zo0wmDq8m6WBHDEVqVxzLKd9b7jVAHxJFGSfEXxz+2m
olPXky/ANbneQZhVTbwPkJtbFwW5QtFxjxSpkPUDJSs4OItlR4biSUIb8JviJCgyLbTGggKyC+lO
H0P0HQlFD1caeVD2YYq/PkjeqULzRY3wUp8ZoFnbWxbx7w032daEt0690eVHWQ6xRfehW+0jLer0
drNWZAZJpFMh8oQUHV8qSrP9+2Hju2pYmjYkD5kGpqvn/Zo28m8jpnBA8gnfzd+O3t8whI+l6hMp
uEYDcaYLsqpDlCUawhDd1AK/icvdGoyJNQfK+wrDlV8WhhtRX400dBQ67HUqXf6a32eeJARUVQ+I
NWYYYM8fEnzhu0Uf734weuYOKqUT7egQIe2eqgHe4GpIWR8dT9+zQjXABzhXoNuaGtx4qB269Ow9
9Y0ELW1S/7c//SfmbLLGmQB2NC94l7QxtvJQ5yGMe38cFiB/84w0C8rfcXdL8IuLYZWJZEPEm5bI
SxuYQ43t9nUpbeWYaZfNpbaqFaj2uNwweGzWPZB95L2RaMtMzfSw1NQpUeQqBt3mPiYzpW0jhgPs
GSClOs2v61v05AcwHagKXdQOAk+Sd+qPjINTgLIlzRm2mAPpAKJxqzen29KXHFEvIZRBuBPQaZib
9SFlM0k9l5r1c6j6M7EbHolOGT1o6sTNRIDEaee7l2mYaLhHk+4wQwunmct83yH0h4l0h8i6c1wn
th1KDylKzVpadyUwcaerXrjhNEHDrTxEiRu/rxPYp+bYbi1xMweP8YL2VaId69iHRDwMzz2PH2ce
WlrgncqpxD3y626v4QsB4z30dNuMYnMQEszykgo/HcLObnKggAR99wsJM778xqB93C6FeKKdZJDg
VFhUBub6u2zDMkaeLrqSgRfAtWQZipW5nnjWarhM2k42HTgiRlftM9OY/iOVrn0KPuO1+4qwSX27
E8AUG7qU7lX+iCihmSKJiRfzoM0kuFVWY9B/46Bku/664sM/IBVPlpngBGvUfvbTTFKdJ+bhkbn8
d0EqfiQkoLFQbD9V8WwVVteexUgmwjU9+JBg44uxs81RU3Hgx149J4+/YwXZz3rJmlKay3Em48U1
hQzYwY9ymqHJvtJuFNw8YQA/2OjC/dlXzRzJK/TZ5j63bGQugUf9N4FY3eegm/N/fJ4r45uYLSFB
ZqVGS9XlmFHRJznkF4jJflwv4vYz4qaWjwzOvKovDFvyJLODGlmO2nE23ZTZ/30CW8Q+kDd2ol8x
WbTvVELOc1+23/MvADEgKrWi3vhZLBuJOyBxzZfRGuCEn4asH6hKUK1SHfLxS5GTqHvbXL9T5Zev
MTIiXrYwLvln8dByWSdFJ7NlQm0AxQepFwCYpW5AEwsO+JJWs0fcV/7sHEFPnEW4ksnUnABe+IGw
i4EhFSplfA0qlazmuReYqz+AkJSfGZ3w+lkaX1EYube3rIDLWiYwiXEVQ4OddzE/UskHA03L4q7s
gtRz+xz9ICvwm/g40XFh5I2s7KC3BnTAVTVZvsc8WMSUSC+FQbozS1RfOKpGTAf3o2tGwiiWKkH+
BjqOgnUOVaeYu460vQYnXPtLPzBaaxWIEH50+zoGTqjLwWr62xKfb8hvzfri05/ku1tKSmeMUBG6
ttI3ruxlBOq2eACvOT1j6c/g0FrvkwSKL6ZHFrSu0Bwvw4SniejNXwV6dIwkYb9pc1EEMifRjfzm
UnMkVQEAR16KfHbPYHt2UKf5WcMtmMQ6vcaUlEIE1N0bQ8BYnYtsPsaMf2LfNJeiCHxFZz28SzSG
Plls0s5qPHn5VuJWa85nciVKhHMkqwn4BpnB3K2TlGD8847GPrjRmqh1lsDJGW+KENDqzEG/pQn0
LbMuuuzZyQOOn8lR8TAB3bzb0vMV6xpyfUpMdRQ6NLnRgmsrGQycms55D5xRm0X8/naiMy+tYfQP
J3wThYKte62DAB/DMo4rQ610cGUcw+QCprtGiyFTcrZUnb2KnZVX42j5cQWYJT+sgayht5Qullul
gAlRBqyG+w+QFZmFqq23rZkm1PV6pCv8tbCeWyH5YjzsEbiTzA5cxCXrYRPxGHc0wq+tSo9QclAF
vPY+eMYHtzjjaQRnDaEWVAI/47D7vqy9api8EVNEshN5PSy+SFbpwS0lFhkofncq1KNMNtqka6fn
8BUh0yLp1TcFTMz75tGe4W1Eg1CyGFU6SCwxN6byDJOeyJBNvO8/kay8G3iLtc7DZ7DubXk2mfcs
kiI5FxmR3lLnRg5FkN1wbBDnc6aAfm5SXJm+Mq5jRMdKLsPSw5NUF7pCAShhpaP0/I7QwzD77z9j
TO2Y3/wAivehNGoEe/skN0VoIpvv8yobQp9a1rUKmK+yceDCdZrcUvWYB2rwDES2O557UNm6MI2d
GDP2dDwzcq52GWAUeHqIPfb8dPH50r42dSHWvzRHs/CdRoFF4IuxcJL9WKcwpO7BndVYPyzb3PkH
gbbBdLcP9Yq2sZvmNNsEMIh3f2390flIEIuGGS/FJDFwZO6scIiakgqrbTwd20gq4yOLByIph5zU
+TfiOBfgHHrWI7PT+Ex0itORfaQSb6ba4loR9LJFLzWQOe6nVIk2tViaAd0OkcvjI5gDpYT0TuL4
ggd2C3vmxo3sXxtSfEXUKgnhotu+3yrV9TwX6icHHhYlZ/grJYr6cTugQsnn8nY2rMlkwgjQoKI7
cJEBQs91n9ceKfIu/EpA3E+gaQuMHy2lIOCsUU/yz4UFTH3a6w/gKFBcqLAVezwE4T5C5bjaCFvS
uSOfgOeAHxEOoLiao0j+xBZeoyqhzdOvI9nUmx5gv0EGYdCO9bjexVkBA/ofbi1ETo+zypaUBqRN
wtjkGuo8ETtXV+Tx41ycH0L0Cs2HLNPptgXhTWJjRKPEJRkqY4JP+xOigbECvZLmjjDztuxCtC0B
HXbU+Oa4iNDWiMuwOgx1tNLBMxFsHHJ0IRJfClNrzhvXPVDQ+QjBpeR/gFhhh/cKGdXjL7hWH3El
PJd6QyrwowqdlHaf8LpM/C0pV3gmF94aV5DjC2I6WweABuTYpznA0PsjlCw1yp8vjdnAkeX+x81h
iDA8Gy67Pl1ez3+3mOPazSxyGnuER7vjRkCUiLPBrTdEARWVc3ex1yG+7x7B3RHKbX8n88b6ezSy
EaizialoDy4RwudRVfrKSdRT/6SWTWHFKEF6OZjTnUY2Gq+6kLG7O0B5Bn/uRm2DoANF6KijvuAp
T6EwVSnDV62ef2j+kWKWDFxoD7IZ6E7Z3brkN0E06VHyOs0OIiN2XNI2yqtZh8/F5o0cmPGyBoHc
eaPAAF7ZXCWa/Fj75m3QSUK/yLpAewXUrmea+9zoaokvu1g63xD7YPyX/No7UjqXLlkh7yshPL7h
CLP1HqBy0fgQ3DgiHMl7hJccyhihnRE5kpRfF7bjeM4J4eni5vrcdASAcMZuqQDXP2c9qjUtUo/S
Gol6wIE6CAR+WcD+X53/5i464A6rGaVUGZmVIemZjGs7wvc+WxHuSLyZ+fWIkmkE9CLIeESFF1de
dhInnwV/xUQuxZv0su+NP8X+tZWSX2KvSQSR7MDf/St9w/m5oJ0tGd1LYfF1bVW/FIcdA53L55Gp
ONkmsdyt8txEcrAGSeztHhkUOTTpBThyVStH4rs+KzzPae6o7CrxqtQn2J2/bAMfGdbX7bDnufwx
R0KlMKEI7vegSkMEF8mUm/bWVs13WiUtTTY1c9Q772x93BbX7AgKtBOnk5w6fkWvQk+B1QC9XQhb
b4UgbP7BALFlvAF6wlXxMUBq493f+tvCRrpvt+FeXY0RyC93gFb/v5KSIB+pIZyYciIlWv+mwqA9
LBdyTLR3tYAcPdQ/BIzxdKKeYSKqpkbqbqMhP9NIQJpqF/qLajYyyHFLwSoxgxMcC0jONOriqOdD
SsbaWh2LTd+EEYSbdgNpKP8+2gybSRSMv8HL+DHRGBpaJSihdWiM4bq0s5KBPqAfjNpriFmIRJNS
kNAgj+ZPk1NDvzEb1J+djvbwCPK60ut6SWSi/vMLmrezW44KpdUfeXda4yzZEjy9bmJIY7FRWsAg
nMVOyzyOXiCMfVvfEaBgfsvmVkoIgUczPIS7rSzQdcm5l2LQ2pcSldAXA1YO+jnP6LS5A3Hrt8w4
LWxi7zaa/8T6nynfMWH3z4V7Fu7ShD6I57ZxdyqE7EVbYgSfKpzcADlWRE/madvXCQtbyUIn1mm1
mbE63ox66o9fm27o9QV8EGHvQQJnQM4dnLg/lotkqWNMf0gJClHSa/Ly7iZocc3dpKYHZ+Ir5d+d
Qfniz/ytS2PHG8WVuYe3hAjnQoqbbRdbkO6ufeMca+3xZqOGWWTidMsq/4kUvtd3osRIE7MqYT87
3iPOWoxI0yMdSqkso+pkjKKA3pX7Rv35Ym4C/DZ9WHsFg8cnUJhvb/nP1GkTYfrFqEhgYZki/xjy
BMDeCUlc34XaWUXJvM6tRI1gCszcvP2B1L6fZZP2qu4UFb6dp27sGKrvogleLMimdaaBZbLBT6du
2d/5yTeRK4pOIha7WjLZ1UBp7k7ZGgVZ1/uGLpMJK1LWY54bZAdgmayx60G3L662fXGIXiIRXMe9
hpJIGpQ7Do2Dn9of7MLvRXru1ME8QIOCJiqweOTligGLagZ1GCmxn9g3z6Il+e1378vi3rNbbn8Q
yl/9KcAgCbX0t/DRNJ/381FQ8O30Ti07emGYUBBjJaIpguXts7WkJxQqXKsH43AHhnEsQvJRePgZ
cf79ZIuu6rvrjudEwdi/myLH1n9eMqOtWqNABcLZ7lbNAuD5Us6fH4/LZTGhZa7p0CypitPkMoNQ
dqm4A5P6a6ShorM8b1qMgvruzS3BzIaxBPRir/ZssLe0SL3PV2eEOcwkXClHsniQUsQXco5c6UWk
iH0uT/M8jTwH45JApTnzCJZGY3vhq0CLonjTI2QO8bFHDB0bdRn6EaEwR5CcsH8ABE62GhkyCpC7
6eZJHCmQycW+lyGXNYnegykViZeUoBdJfC1Nj7jIgtyw3XG++miFUzyxk9AB3gWl+aQQbbawzsKV
R/OKzpmcKykCUJQcPQB6/ersriWDWvJxfAYTZcC1c2hKwQrd2Y0cOvd+cwKkF2I8p+BfJv0POIv7
hibohmeYR91zFpoV8uilCT7gbnnRv33FBjWbjK4n8lqYj4U7jwRUIA92nILZ3Vj6LE7rqI9xXzu9
YNGGUH8g8UH62X8hsmigg2H3/9Gb+PsR4RKXM7IiXpS5KC6Yozw/wGnrpd8n/hrqlpyzaBJ0ZNle
RhTBMlKERhs4ZtHwWjFXTAXCPH1ExZa0XPZf24QMErf6znbFCSRjO7+LhmJrtPB5xItrEc4rXf4E
606BO6dmdUQ74yS5+uNRb3E4/gUTIHeY+8MNaIQBy6nGeGlV2STk8/iwitfZf80ioJZJZe4DNv7P
YqYwXNbWoKrm+AVR43xCFdy5jMr96vT4tYMWAoWoNMNUh1JmmQxtSdpA9R9r+TpuFTNe6jEJ5LMF
gkrawpL/Iy0TbPV20bBDWta3zoAH16zsysArRYOOxWStSxeJLvSwsYhpAzsRsv/XDbQB8/iL4ajQ
Uh/KqFb7dT4gyEVX+2+U8skP1CBQv1NAtdCkbnUReyXrPhgd85giDVf3Y5Q8fcbiAAOIAP61v84a
oBGkGxxkDjp92sO3UHHcEO1oFjsEXWOO2y7K8dLV8kwgMMok5fw8q3Y0q9aZS+40KqtkVj+rmh6X
NFAXKcJYPnXEY6bXhE5XHspW3SmMZYQ8LuusMy38xa8FPylhRZC5ySVDBoabzibUQ5+bh12/VMRF
cTRwm43/5IUKbeEC8nMFgdep23jhxl5NMJYW4dNLnQWMzTk4Q6BE+uMx7JyYea5AiTeOv6RUKeOl
uTegjbXcqXfp8CYaNHjjPw67m5Tbh41wCWfDMspJ84FNTXKGo8bT/Lqn34uA5D/BVH4eHDK8JcGJ
ZBmIcU4VDwaFWZXDvHFe9V10s2+6vI1K9WGVe1PjJ8bM9VZmcDrPYmoxAH9fYTBcC2KRSinucnQW
9F34sTNwfnYabrNJlpINNywd+X/Bdq8Ctxmcf4+rWxu35FqrzFZkFtsCW0cJOkvTtckRpEKVBoiM
Tg6X8Zub+rPDr5e7Zh7EQ47HLO2ouMXJToeoytvVE09FnYpHtRPjawv+8MTYE7gWnGO24w1/kVEK
bHbc2ZUEH76uoN7YNV7k1BwbNxG52D0DnUeGLqhgHlYBYzeiI3DeXBGE0R6Cga7zlIXN4J/LulUh
zti0ePgoM5KtUE5ZHl3jXXusYUCEsmEdskeMoLtlMVUOZ+z34CUgqaGT3zFMrJlL1yXWLRU/GspS
+I0IuaKEPjcLcy1DzNSqiVemcSvsMzOU4vko01VjivRhluDwgVZRuMXcWEY29ZkHaKDsxIYzzXRa
qDV5jukAPHWSjwawGXaLz9SqK77vAgciMJVrlCqm7vk0zgRiEipxL3w+iEwiD1LHUEJRR65BXo9g
ba3gPXozREXM0AAqgcBB2bvW6jP3JfiFU0o5jw04RO15QDGe6/v+3t4uJiuD2GGD10fUr/pBpcdf
pIFT44oOc55e/qwqOydBRx6fm0Od4uPb2EFkDGmF03SmNog5QLH7FNsj3BUaISPYeAe0xlp5hhNj
AGPbFis5bvNrE+VvrijXKqe08C+6XJBwQT4x4HwArR8myT91Fh1hHErBiu10Md9VNJENl4SRWhqk
Oi4TA6BjbNlfNxhPRuqI7WhL0LK5E88OuRSIbZDNS0Y4UhAk9cEiSC+qmNI9nqFTpBV1ppA7BL2J
2gDExJT3ChBg+qcd2Qo3iy/t2jrLD4zSQt2VUOtg4WtRHzVT9Ed8XCHmKJlDoYkkVD4klbl7RiMV
xMmbhipXALn0LyuiT2oA2XSeTpfx8AaXH3zQ17ibZj7aBRKLvOgv2F8njnLxcUc43zZ6g+bg8AuV
aDaHVMJO9ue2gSxgrhVAjvgSAvOuhifxGHoMQtllRm445BfGYq54o2eshTXhvaGG0+cbIeOP74cT
nvWhlVnvBVjNqlFhPbUhGr1wVA9mi/G+J8orVRlntZXp2nvBTwuJcj6aM08fHIYS/8nNoQyhs47e
nLJvlzc6tqUxoNysk8wZ2pctbO3VDdVQPU0lMc8FRXtUuTaZNGEeFugj9+wqXMzPMiORGIkNmmOB
uSiScBg5Tot+UYiAj8H2iHDuhU8UAenty3pSFGvkCehXQOQBUyMVHYRgynb4858MbrpCeXdHzTFi
ArgZCe7hQ4UqSV7Lv5ZGAAFZK5D6NyASznv6KcwSHAM0xk6UM6W0j9BxXuFzMB1FoO2QyGnSKe7e
+yo3QKnip9qbaij/qUKGnG2oF5yx+W445k909Tx4x3uxtx9YUluGvMt1Y47TW6lCPbZC/B5+Z58T
6FfPDEJJaLptnqTUH/oO4pgpvplCKZEpDpe9yeQRJX/h8Ze/jGUOkmDx4HMOtLgtpYqkicIj4CfD
SVFX5sOsrJp5FTc8FwuwR9v1Jx/uQOwws+IuB/hScy8Fg6VU94Gj/R4fAW8HcYAPgPlzFCbnpaPn
xOWXkveY1IshUfZZFSclmOhUpin+REQV7nDEzgcyFLb6IDZUJwLubu1NJD+TU7EkAHFLe2tThdwH
fv6sDNWYQ0OEblnQ4U1jZGGHxKun4QSlnviGeUPKiiiEzHI8Yj7H+0hxIVReT8/RQ4dnEaNTNqsF
BBwOo5eRDajJsCMWqciev5VIRsGD0F1I+RNhyjRTnMMx8JlYrdMpm0vSupjnus7xbNWZfwoTeRbu
iwRQ0Tx+tQ2YjmkQ8soJggoicLmXIknoXnVoBIgoO5j7PFz7NnYGf+OxZUgmrl/ysnRQsCuZyPgn
UytlvaoQ6KBuRuCdtiQ6uFfc3dl6shiPPNDL0bxoBO8FDD1VGAkvL10fkS38llTCsb4lhUN30HBi
hqQEUurKtaQHGW0fF9FHGmkQVXzI0KjO3KRS9sRe3wcZ1frGmtGEJFKZPxvrg4FRrhBv/TZmXVJZ
Gt40EzpAEyhZixQzT2GNK2pTmoDmTC6WfBTmhJSVSwKq98wl0Lox4yeqntXAjh/FgLFMDXtYhS2Y
cIGWBKhVH9Dhd/7LmQ/NikArliC8FLSLbPMM+6EKmtdkPLA0n0V984HQjybUxIGKbGKnKTkD0pJH
TddbVhYYEfa2u66GUXNdjH/4RmoVtzm9ZUS3B+cOIgbC6KFhTqeYQLf/kA+mTiUfpkVb9oEl1KXP
CBjBkZl1Mn1ZcnSYPsKujYn+kT5fd6DSWtAADAvvv2i3EgZh3K2YM6YWN7Xqtl3CA9yY362ApF6g
603FCTdkceb1Yu8dpLAqySxYxRiKsF3v5RvP4C+sSCS+gOC/k32r+gf09Rmx3MHZXMBNZUCDdNHO
/e1sXz6tR2Anx7LhNuGIarmlVI5KK6Y1osK/VzchUf+OZWShkBd4K86taemh/9fGgc0X84Gz8L+1
Z/9uRXtB/M45lH/OcfELBkAoM8JpEuYMJ4rLRpsX9JqNvh5+5BKyCc3HNVAOnaGhgGNPaUJbcoRr
9Uvw7DzEkhmox/U4q3nVvv8qcyIMwuao2/jLHJkzxQM0jiGHWBqmNhAPI9u8FhIqzemXxYMSeZgf
kIsbG2JmehwRQiwLyZWiZiKdfcstDtgTrh2kvNUzwkK/kEKtz7UAlE3ogfFpCo6H7vWqkXa1ZJjm
TQIWZJoyztLcsBn3NxkCy5lUF3nNt5R/1+/1dJwBbmabXH3EZUDMfv0HT2icPfS7LyTk42iJqdyb
p6Qs+fqrrTLdRsTdItichYB908+LV/piBIKE9QGywxaiND4EGNxhQEAzoctJ3jxDdY7lDbmCr0hf
Rcmszjs/D4vvbMBDyNCcG/iQqT+0B9v1ZuOAY7lg6pW1QeJM3SrRf65OrojBAkYtV/YBDv6q7X8a
a6CKUPiorM5zK3oawhlks8g89nj6bUuRBpZFEiYNALRsZrGaKN8FKPHmM/gUNLyonb8DQ/mw5XVD
6sGBXic+8qWJNQpKvUs5QBJNZH4SnMVvtItUav704YsGYQo9B1MTsS0/rDi+N3Alkfpxg8bMSBlM
6wwHVQD91WyMyQPmltkwpQusVv+CL8wPQ4BZxiiql482uTj9okrePhlTta3JDrLmfmz6HNLUi/BM
mj8N6bTdcpzv0V4YROBrdIqhjLJUVyXi4thqvGINk3TZDpncY/sQCt17zegZ2y0CzUpixcZZdNAI
OAaObqmeTNfe1+/gPnlKndf6KoyRQ8nzgztb51P2IRAexOdM7xRgomelIuYPSrbpCQD0UpWgzlTP
6FZpzTUthg8e0SIa1SWbwKHE+Hc0QZRo2lLktp1W8mmm3ytUWaPS4XFTbaUrH+FK/Qjajs7mjE5S
OpCp0Knm6KWPV3y4DHb0ZVnTMA8/ZYdy4SqHar5oupACld6yPlEDFnmqWPQl8jlEHZLjTGoWtA+y
7ayetjo8ttm3sJnvjdnI8ihwa13K4FyQIfbxXkWCpyodPdwhXic+WDQ/v5PQzQEYJ6HoAnA5p4U7
82Yac9UhvDbV4cMPyUGYjsvqU9gueUy7Sqmohc6kc0iY2PpcJxg4COQIMR4vseQDmvK2IFgvQjNp
WakS98/+82jZ0jByds2kt82lZg4pmGCqqGpEotuuIRcrfQAP6BD0pal+eo3mAK3z+VkwCw7eXpI9
Dw5z+g08kw0T/BThoHqnOfVc3rxLjrFtOQumREO0HjLgjicaFivQmovM9tSP+2OIyxVzcmWjQPl9
XTWOSUvrpcl0w6zdixm7YgbflLMn3ehewpn4mUqdh02R/BzpRTwIY81tdQz8rdCLMaB6+StP+isI
mt1gTa32fdMmIesIBXEyR1i/tIK++bVQIctoOYqQVzsB/uehgQcpYGV7cWUmoevQz9mIIkIhX4+p
YOE3FVQca4Yj7NV99/ae0MUfXheJbaGMlYuULseaLOnH0/S2MqZdK8jB3bdBodP+kaKnXPVitwYZ
0REac599kXWpLxtsOBhHOLv0dB49W1nOVhmkYx4dh+AKBLd0V/1AqeiMWneNdj5EWwP3sSO0GE2p
PLPID21jgsALfxK03nI4DhWzsEp3B86LU35NWgwRv1XPJM7XNeysBe/+OoPht1ItJ+RQAQMOJ/k5
tyj7izgvblZq4ZPWSPWowjYdRWkrGVgT826cge0Fi8DmZmo0Q1aQ3n7EcOsKC/Q2SOt2n8ugp8YY
HVA7u2HMufWgQzyPPcpP/0I6HTlSAJtFjT9U/lkADsp7EiWr2mazPUn6kL9z4fgU6ftP0GD5JrPN
YJNsbSv6D8FZkcWhmSfyc1AOoAKTEih2C3V0IyRYzdub4L2jltwZkEI+xfhykY+xNmIbIF2lu28C
vOy7RYNPjlJuMF2eRBGAgt5raZJ5++WVEISpgy3N0jBAkqxZdyza4hfXZtisd0plj3kod4BrFX6E
uzLeKiX/Sn1OSjzvUjDNkR1xFCzMBOl5hnpjf3t2sD19e38ToMfMbz0L4ioQY8XC7MFPHqDmwxcw
I2PJBXxAuHKVFY/nMyxdLCzBumx9pAQTbCaJx42AeH0LDfqc9ZS57saftMNZjmrirKgFbiP2Lvft
legzS8o6C3zBnRvxF7Zufzl1E9L+eJ0PTfcl42bW83A2elxlOirfyrjZSUx295pklE0IsUrUAmgN
ab1KmVque7d/bA64DYcLHPbY6extc7g5CXpSp4KZxhYKFyPXlZO0AJMHePWyOSfH0VfYmRuBEJu5
pmlinJ5tiL723BpWOx4y4QKTdIoo1i9diaYm+w6gWTJJf+jLjMTJjASEzRZYwQJLYOVuDCNzRtlC
+FFThPV3RB7yZrQUT75cNz8qU2tT5CKYz7aqTCjbk121TutpnL7R604uRfGef3piS9uGQwbazf5L
r0VTcOolfv7LfvAqvHrSRDyxi9hNy7HyXxHOdsjA7GESL07yH/J/E2qb6NkTcp6QuSv0klfg01bg
E6xGI1yNOj2dYHBUsVtHKE1PV9E3MEAgOtPRz9wkxDXAx67y2BYFdD0vG/FvTiKCrozReDche4Dj
BKnWWLPP/9HHkoEeAGChwZCmGOkvmfo6d64mRmp1Fp/UZBZncymesfveUumIdVPMI358KWQDxABT
nVQArQ7x2TivcZYD2wM/G6eeY3v7kb1jkV0LmEMLlSvblPL3IHh2jKobiAFAtIrtHOd8ca6wITSV
TpKXNeugd8wt+cNhl6h9aWCsjR8cHO62kLcZk7tOHI/huQIsw5/RJv7LDIWFMJAUgMpUzA8ODJ7H
WeTQO6JZ7X2w7vq1ir/k3sfZjAq+aPHmxCR9T5X+oI7iQ6Z+XPhucdjIfHNlBs6MM+s3GiSE5EV8
hVBL07nGCU1npPDnvlQf56pai2j5GK9sD2mLuPdez0N24b5otzNUHicdrPt3rS3Bz6vDbVjDgzhI
wVS6KmFtw9DgPXY6CcFY52x7D5l2DYPdu0ceQUva7OY+2vawUjJs3ovTzlL30oWxj2mPqxe/L9rZ
//55KarEe5uzWwKMIvf5BB+no5ejxf2CBp6VyLIOAAxEzF5qQPZ5yYLZW/sbYzGUzqJYUqRDepvM
ehi4QulVNfO7MvSi2tVEUJJDMmCPpSlfHh/i8BjoKU4NOd01GPtbOu5BEt5fbllGRWjvTIu/IJxi
jviUmsxq7AmYY4g2/Te7t6ea+A7A6dQFzI8QFUckKwD9FoNu0VbCQmySsVwk1Um8nByo95tNva/v
V0804bjInT1daxSVxTPbWxd8MnKN6eZ6z4gKK4d+FBBmNruboN/Em6I8jK+xSJnHs1z5e0d1hl0m
nT11E5gv/gGteZntqJk/fn+NjJH0MA+aTuWbikMTwKaH64u+h8J6Y0cY/WG1YHc8Cz49fsd9tOS6
C8RPc6lIeAgmmNrgzphDlhMnMGnxKQ9ciPcDwQs1KY9ZXgKSFNNv9JErBahejDSKXDRqKgaNSiH7
QTDHbY3xOI4o1+yPawOKJTMQ/v3AaXIBtnsDbkkdx5N/6Y9HKZdhfnPANqR+GVje6Aje2R/ubTuh
oQgzfoqDiJ4hMEtHiH1bLCZJ69q7iHcvvkEQuooZAA7FIk7UdSVGfP5FSYDAYxChfQfIPySzRKof
xZRov6lOT7TwkhtCMqAns2ohBkBeeapp6KAp/gaTeWwttUdi2IzU18FzaxqKrJrn0K6PGdZSjx9S
7y0Hv3x2rO3kjuPAsoowV5ukYpcz/qCOUTsFMZ1cr20arWgr+FTFVLesWY1W3G+Xk3xHvbOnSiGz
a1r4dctLehN7anPpmt6EuAsrn5gySksAS3ZeM+OI4fbOVChT7qS+Mc2PCcD5+NrLwu0pxetxRxu9
CqHukG0NQ217YclbdKbt/BGv7DHBs4XaRuItlZ0IIYZlRTj3yNYy5Blj5GvtYUpxZ/CWYtLfWv7c
jbO9F5nqZhPCHhP+o6Sjj5TolhrqOkznYbkHNjPi8VJ4++aDnV5ttM3iQfscjS3/rsuBmBMnjCeh
KBOLvTzaF1uiB4vaDTx9Np1ocZOEFnYj//QtuDn+Obci8eF66l0ntJf1cZMW9zTpZgcBheLiYUoW
LClyBaXDnI4huyPtLaic/UTdEH6IPIdokuxBXkm2/kLD9yCIUtFQjIIE8Ch1eUKKXHE0EWfh7mBJ
EpliHceRCER0ZW2R6piaDziO7YIp/3w50QFBhvZkmdZRltXQ09dVqlnf7fneKIZ6KWB2qiWjJqax
YmQTwN97k8+4k2c7Lh/Rc2IIkf0x/ExZxfTQcneJXJo8QL/9RVQUxmH91b+m5prLo8azKS3/GHU3
BaY033LLuZDkCsAc8Av/g+5kLcYIRfdvKThcxPMrzhSISRzsxK/Vr128He5Bbgpdi9OS9mXkWlpr
vrrozKqIQuwFMK8NJvg8v7UbiNw6liFCBo+9qEfHJDdhcvU+MfShWHjjqyDXqfO4QRnZMKfOB6DI
o9B3XeGExt1/T9MgW8nk4qWCd6YNM3bRxHKk7bxM+TQJirLmpzapUdtrytbHJeOpdQmbRyvzvpZG
3Nt5hc7s+Y/38RaJmMuq4hdrDaGmVhDXFibluzzH2aAaJE+O2UVXOyFXzmkSkfiA+HdacXcVt7fJ
f8Krlx5KJBmfd81l7p/PclPLV0i3Ux/lBT/E7D1sasKJei7LUBMtzQ8vmdVHgYmlnrpfzykAEGhS
MjXvdH9YG1yckPs50jElnENm7G1a+tFUvgCdac0f+NMoUW+ftnnMWATv2QPsCCjgNyYia7M7q35c
YkpraisEtf0mXIooI1lrYZoItNduqbPWAu9UQtA/9OvRYk3UMUi98kgFoJwEYAs9HUSXfkO4VV04
6GkgtAO3qgjWi5U56LJ/nYqDspxzSBJhnlqm8gEXDk/QTUKdiA0du/S5RQf94q3gqVvjMxeFyQWr
0osvoFhL519IeZHNt/Y9bNPqjDKWaTtKwGDhyyZP3pR3vo7GD43i/hhynNacJJwQx30m9XHyz3tR
yaXq+Lo23hAMzOo28LEuLUAedOo0GuekJ05JTtMmQav8GI7Ld8v9K4QgrPkex534+ImAcbCERDT9
W0G04Oij0ka4MFKCBnMhMVxXZZjPt5wXPBTN7/Mk78TzkYO1GG46E90yPuCicHWK5hjG2oB8xlGD
IRZAGz+7S3GHXJGWOnxrPZednfv8kLN8sve84CEsYd4TkX+OD8c8FpFTGx6sPJyOeA5tRFG2FmXD
CbDqwCydGaqeqM2IFNLIc0W9Ei7tQC7XNHZdRiE2MKnBcVNYnZC/49x7argy5nz6zNZCo1FxDcQN
qM0EbwaVAlFW8YaVpJHhbD4kwELe40Nx1PUlyGvLYTIG4QfRxskXxBGidDBiYoi3g8brGiSNEPVy
DDpVHCSqYF5FFfLP20xYbuDW96YZCT/pRHKNz89O93FKQabqUlnDaemp6TkZ/EK1883LOxBh86Ev
IUB0jRdp/26Fl8k8udeupLWCdqAD4E/jXD36ymvWty35ob4Ef4fexPz7sb7rnhaNv47iLF5uYcIJ
xk/pUQz9tSVXsWgSt+xpNgInHvXEf7+soYgFfHtp3LhFpXPE7C0gmW4vxM+eWclqtsAXELcGHCXh
YBXimUtpyTi2EF+GKKIAanDzi0F3pPbqiMreICtS3BerPb/qDRXpyzAj0zehyFTcf8VHRwZvSJgd
nsNbBj6v8FeBdZ2b87cOUs1y34xMONR6KfJ2T4u4V8sarJzIRPSfo80CBEVJRuWee4oaRZL1cPek
KwokSSz0DDbyB1DI45/BmSBrLLGjunCNxzuLRVSvEu5SGD9BBRRaE7EUBfqJQYtrjUdNpEND0IWW
KxH+eGBoU840Q5e+JDHCEk894HLha4JFF2lbgS3yWgGr2qB1ZGRM0PFownqd2wx+JMuR4e7dh4fX
zuGJrI5WU2CHaCmk4SRn1d248S3YHw/r1TzghqMJ9zmGoUzgzbLUrpiWd27Kt6/IHCkdjFxZq/PG
KM8rtYw6L+aB+iy47AuDnmrD5jBYNxTX/x0NG1ECaIRLX3sYv2T3n4bgrWU+rWSPUE2eyXo8ZyNu
uOE8fWxh0KXjz73zX9KgLf2ZOaYsrEb+lOu19wY9gweObsjMmQcx92R1vniwVVTuIs6eHceTTuZj
MF7T8l+PLSk+XjJd+V0/95d4O00x5FNuQuKyZI18mswRkFZ6GTV9FAYH3MPPza3gw0XahJf19gdG
RffHYZg9FZOF4/xbDhTYW2MdPdA1Z9WOWrSaF+e0CjZJaDgqyB4Q2OVVXYQ4epkdqkLxuT2m71WW
RGb0M1vCKFsmUAZHv9ZgZo973pn+mC04wRkkDcjL3MfJwqXk0ZfubE9v9knTPUNlBUemIDenilJv
ll3y3qld/PctGN32Lrcz5ApXhsEW5IWug69nsJx6w1TQ5e2tV8rBVHYM2fu3LUIR/MmEFJTWNjNW
x5jUrvaIJSADUYTAu5EiwWq1qbSF4p9x5AAfCJU03WiY5EBw2Rw96hAWBK8KvTr6HiS7RIj4SU1T
MCU1Wx9HrglmnNHXPqNrpw4TP8/R9iTTCpQ4hZcI2MGlRbjs9UUBT+zR0f2i5K6EwJU9VZ2wEoBS
Dd2RapEcZZy5Zr0Al1e74EhcLsMDy6CIsJVqfqej2ppHT6q4cQA13mRAkAF3stRBX5kWcnzgIcqX
0YzMZcBC9U+w6nFvkRCdwqTXPVpC64sPaHYo9CwVKmjF/eliBoSGUcL0pj+t5TaG6oza+b3mN+/1
GiPf1Jbu4l0P1nJCsLoiWQbYi1EbBkJenhLUY4wJ2s4fEXFBoZoQyjKPidNuqHwGpW5EoPOMd4n7
/6N0r5ohRnvL1YnR6ERIGkZasq1/YDRlolbCThlXdQwMBfB6zgol3zVwqYHHJGhwU5Zn1j8YMLGR
UgBRRyNYGdoJs/ss9SibmtMFoMNxrkCBSAyJMEzjZOIt3GryI52NeEEc/d2r0iZ1dg7uEhODn4hO
Mw3hsWD7xPxUrcsWCNKEJsSB0dChOBm6Th16MEzYaUqV74uDJvdSHgH3YNYfutvvzdc3zleayGaa
aX1c5ygUyuhk00HPGFxeSZFtnIHXUYCJTsI3V3reZax/NE2Y2bXOYlxU8ZsR4i3bnz0XQtT4msGX
IHmv/CeQbXMQ+z9OIrtzblRkzj7LZrbjs0FlsIlaggF4s88Uz9AgrD50CFeErnom5kMleD58Dzlw
/+Izs5ATJo1jBImGEx6iNBy66nF9oLQTexEY2SzLnI8J03GCrRYZb7AsTKSgvolWYszvNaz5zigI
ahxk2oro8zsydmb5f1bdYDi7Kck2TFiqxv40qkOY8uoYWSR6cXThsLHQ3Ak69CrwKZIyuSkQM8Bp
pMbLl52Hc1ASbFXUR7M7ArxY2muAc3JgbFwVWre5zpxdnPFGhAgvA4TAGhqb2NMh1w614VakR0pq
9am/mPHGsfbzFhzDrgVyE5PY5sQBMDK7uiWtUu3yKQpU1uU/gzbUZdq3WxUA5CRUFvaA1V3yeIdR
bQd35j57g9SYw4FDyu+gIq179mcXywlYmZmwxhbxmx7m/mFaWijPcLyKRCmO7X/wDBqX6yRJ7pLN
7yCmagF8alMfujpesRR43pW8EmHfzXaCSY/HliqBrsSBVrrTC3YGmfnU9ZhVIYjfAv8nri2aUdx1
NGB5CEqFYLxcxaMh5DWRBJ/PVIrkpeW10YZTrfRjFYlME8V9fLs9peklNeXLkL2+gsh5Uvc5Qw2/
csS6KqxDrb5fTFs2e3NjQQruhAvNDypSO0t36N0DmSLiuBLhldkcsCfM3alcYztkWUmax4UbxxWD
a+oYTkM48c9Q2Gz9fFrVGVyC3cb+NqPX6t7/K+B3Rtkkqxz44IoEnl6V2oWOIBDwEnadmtiwXykx
fc3DgFuiGmyfQ6WjdCWnaxK2wJCMmXYe5vTzab1/xH9jO1BJD6zuTCptW6rRvavpXmB0MWC1yvms
75erosT4n+elj14pp00z79rD0UKnky3V6MMguBp0TfcEQ3fNcngYa2LgADE80uTq5hesN3tgmc4M
V0Gw1apn4Xp37eppu55TJm5Op9W6vI5URA3q07fZGtM36thesN5pFDu7jA9iyEUaJVpPiLvIDsfN
/3EayLmMb4sdx3tcTJb76nDitOtmvM8z9Mka5N5lc80hVS+xa7ousW8IvS3T5MIt8cE5Rgbrjt69
5H1gHDBVZ8IGFwAAXV+6xcNQFMLgc8ccHUwguY44ahbMmltdLbqVajbDQsraOlWIBUVZHBM9DWct
KrOY6eGMMnXlPkmcGD5nAAwL09/nETMtV7bhND2MVj7ThN2q/NN5iwlNwacAzF9FPHsT5lQqv/+7
5nOLyIN6UfxD2/+9FvIaikoWJv/WDR77p6qKSGTfg+xE13Vc6StTSt03R9vabBFWbqCMiRVGGumO
xKjz3GRR8LERoFbRtY6SEwgNqy/ZvkI7ggeB0JuuUpoZBaB/H06Hb7hAG9+YdjmYrKbreVpVASrv
c7iSA2Njltc+A+4IvLJyRSCy3sXHUIUjZgerbKV3RymEtInQJ5aPGi3L8y7yReppxDlJAVu3fAsQ
rZRS+nOK07Cp9YBG5KLH+JMzDZgXYp9znbG0iKWcteJuMDVJImg8utk44vYLF73Ul8DIIp1dk7sV
mvid9LVfAHASYfqWTWS6M8HYuNbSMcYO069+kgBX7g4gbM1iIZbPwfVqAP94aWHWfcXcjqCoiFRp
14PlZu/ifQk0xsxeHyokTP6xLKKgINuRnGj3PM4KLN0wU3GVXCaJa61GvktTEXuOhCMSmYHJuq4D
n+vuEohK7kA1HdN8Q7KmLI7ynvBEQbn32jehxaA8qLa2gMyTpua8mOx+05/Mj6St8g5oYtfFVT16
Gk21lgciSXQCFU8t8A0EyLwedvdQ8h38ZJ8I5xFLzfqDxc5HiAL9n8xfNdkoqVKQo4on6lU1t+ei
CgAYrrB70hJIDfI2T9nAqGcUSikEVgelldKeZ4yW2nV8O8qt2Ut8Btoy0qLcZduRPubNrzcRBk1/
XIPlF+gojxmEkWdTQKgP+uiGe0uBudAwmCh1rWD7c4ptTmFn5ygpc9/FXdNQ7T8mBLkQ5WCmV4TV
lnNJZma++7EAueSJywuUTjk8zWaM+iecQ52hRc1sW6y/AsrW/wujjbcxFAcYyMN160JqN2uI3bpi
D4qA+HNTEBll93/Kp6j0gkqn321rErK42rdGwx3aI/PcSZTw6AoUcPPXwj98/ugD1HKNKQeTmVlC
+vnU/BsehosyhRJcBKTPfZKiK/TUBSQzKKTJoa2MC5xsPvbzjgH+v4hIX6f8A1rq6gCrRhAO0HZP
cmyAoojBnFHGwg8w1BZcttRNp/Gm54b2S1GWdoXQWYvT+Fu5KQKPYF1JjdfDdGp6ACV18HXq0CBU
O5aOZOM8NG0029ZhmerowRtnEmEOKkb+fY4NGnbkCFZw+5fBTEQi8LYDLib0nRYpyXpFnx65Cqi9
XzwgXLlrHxGimDOutLeGYEFjvWJLLas9u4MWIkLrmP+RGciJt+ZqyG3nzriUUN57v4dFKhiH67tQ
iOLwe4z6vCtMFGgpTyMovclDRRS4b0+1LF9ivFhqlUUDvxZrgDYEKumaxRDxwfUaEif8AwDh+CvG
5F0qB/FyV0u6GDPru1FLy/Wka+oFhtCry3NZSx+GdWwL+qTcLkXtl8SloqWNFmuRb9g63u/osmox
1PzEb/eCMiw02gf+vFvarTtNr1xfLIcONroDDTEBqS55MY1xKhIwQVkt3+628N6oqh3eV/KhMUlt
ljdFPG31Z57JBFIPy/wXFzCB8kfOQmbUpSAW1YwouZC8ADZh+5KxIJi5Y/jfeznjo2JqF2g0tXUW
uMJmrE4ybgZRSRLHgrLVYwn4upzISwDbod26dzkrwA0S0Lv5MRH7M/SXhog5pRUdKuW/f+raa9Ni
GjjGsuJ1m+3K9c6kKBGm+AjYnzjzijmSOw/cV4tQbR7TlC3Ib7QWX6e2+taUHCCc8U54rCX+8hvc
8qztHxr1/+uNRKKWgo4ldLfnGKzGkfuNnJOR/BEgCQJmPEda2iSbPRXX/j4mfbHOBKONiuYdvVLa
VvgjzwmVDHTn2XO9jjn+gSdYdywz5bbOvgsHnbCpkbHep10McIVt3wiEjLKtz0XF40Edp4GwFKCr
ni0jd1v1eCuTT//YK7+IHKo0Xb7gvL//C7oOY884wNSZIEhdK8ehzUCTkNuJaAoPwpkkCy15bhyw
IU1qHpD9szWFMBD6bhQldlhPxsoZJCezlG5CrqyhBIJNxwlReT2ao1nsLL4CpOSutJdIHLDjgL0T
0yVup8NJiulrV0t/v++Xm+5H8oGZJPOgRz9ClNohszx6k3Oaeag94p72am5e+BXv34Me2tfz3khL
psvrOUzU6uKsIwBTOWllO7EBWFEGARMmbG2vCk1RKuH/aUiTLJ7gvBVdsStInRHBpwnZpb6WiWb9
jx1JwXeZX58TN+M/tWGGpo0xvIM7Pzkk5qhouZeRUaSnzFfO4lFshC+2bwI1i3GjWL/R7eBRR8OK
1C6mneC7ptfiAKel3rk8hYvNNjjP7XKVg/FeisBUJQTesneKjot6WJEiDfjUyJwGT9GJvgsvv+7E
2/VR00N4QQp377pbbn5Y93XTZsG0sR7jQZ7rqX5RiJhTqP84swogG5ruP6jVMTTJZdmWnwS409df
8Af8en4W8u+wMi6vJojlYur+s/4f6FCs9HWkfBKHzr4hmpum8jsXXMBDBTFA+PNz+g7hCohyEArO
GXuxk/3dz5VN1yINEn/PzShGhTGBjYToT2ulBFfC6lC67mwvNF3ABVcnYnNG3IT4jrIAQJFfOc2y
Egj0yCodaNC9XG2xBZFgzkTPj2UuiyTyauPn61HyiIJtCnNQFayFi/AcqdspZ7y8c3WwpepPYdAA
HujuLU7y9mhcN89uSgGgcbJJ3H1ZHbbvBtmwwmftAZSvnrZ+r6fZ47m8N7MezPWkxxWLAxASgrgU
l5OoIjG+yg2EF1KPxNxxGFQ04syrXTOIV7j3750hh+sFdtZjhYmGbSPArnIOWeT76tvXrabgzkQK
iXsuP1hukmn7xZNv8YHdgC849LpRqKE3DySLfRjZEhgD5hRKIxBCIyGsIe/JJ3xxXwRPsYJwXnI4
Y8Y4uekH7OccryDkXbmfsXHe8jIzfgtxrYkmGC+b9BPMXdBgHc3+QY44hvnaq/ze0b0G3C8B0zgL
5krv37eiGblt2RazHVZmvWM09icAdwdLcYwhRJOKAdNqm0RZYdfkD+zdnXg+gAq+aXAdzLXYAMEw
7+5wl/Hu+yn9eSLsdUzgccFuvetyb5B9mLoJhhJa3McA/mJK4zf048MxOrpjPcglZ3MCy/cuP01x
HeE1dCupmmRG9hUQydpyYeAWgEcJWY7F1NiRpYCvT75jekcN2z4jzrvW/tYP4M3dScxtp1qEZCGx
FwQWyYmWUiG46wbrYyGcuQrnnAjD7rmSwpvMzJNnVHvSixf9eOqB5ya4Sqa2cKUevUtmgWeumCmr
TQjfDsSSiovPHwVfEwyerVU7KKPzeDyV0/6QVWlvVBOSyHtybkCLz7UY97i1Otzom3lcjjc/iUec
5234rKraWOQNBc6JJF1ttrelKsVevuf+Cf7tlUiFhKLnjXo7zZAUFBvsWAB4fB2eY2RqtDKDP4U0
EhUUJL/M5yEWQuvECG0MpT+xwEbT8BoCoyT/RQ1mj/zMl1AmtZqg6zqpuie72LIdOl5cKGXDbzRS
L/PJY6VUjx9j3n1mXyfgjgeVD1FBMfx7bbHuljn1z/x9Re4uQAUBGuTgsDFydDjkvr+fDJ2CKVs0
VoLsv33u+iHxRlE2jQF2sLP0XSx/zkZrutf5QUkveIVZTWbL3kRgcIqRv2QoXWm9aSaiDCUI9a27
hzIsfyRjlSd1iswHusHUzBs15jJr3g7pVnjVgd0ArjqXSe9nrothCx06rCm65cOsnDI2uNuTYiRJ
+kQgiVa7O7WAe60Miw1X+pxGZUCM6G6JJklGmjwfV5sNuQ2Ra9EOX86D5AcUE96uknzN37ZWznSH
+PQMCZ27QuMF3TT1eaLPZ+lWgcMn/C1bGdmGpkZMlS1RBzWKAGF3F0YWNg6nMfietmHhAbLlJgOr
W9bU7g45Bkw2OsNUcsf6Z7NcEMp7Aiw4Rp94eEPJ6RjdQBA4zhfSrOwAAU97Hur7JN2VL3A7jOkl
89aGEosMfVNomGcoKa4ibTgGOSd853B5Tlwktm8BrXlhFwkyAEwxxqvV5YqGTTu4NP2BM9hDtBwD
/d7zGdVeqRncm6A2m6Sjb2pQxGN3aqlB6SrM96vLudFDdD8bInlYB7aETAHGv3Oa6sPogcBdZH+b
FZyjZaY5lYtjPa5SzqULJR8ryxAF5ZA1u696HkXx+0wToKdKmhbKLPTjhcYj5oXm7RAgBpsvFs0v
jqiQUYwIolFfCBDxr6+gt2Jw3AgbO1ozfsP+avcSb4nc12csOa6t9xoW8MpW/2f8k1oNeyvx3vD3
4UC1vsvR656qabROUZRaKr2ggQnXqeyfwdpek8yvGf/W4/Ylaa3oXmAuNJfph4C0hJyvQ/WN+k2+
t80yGbeb41c5ezW1ndlnUCoAaA7lYnDewwJPEa4dncQkuLOZwM4p8e9sSisd2RKsZWsyKItSPju0
jy0lQBOALb2E165nhnwhgQhpm63YyE2CPgY2lv2xZUuK6TOvz1S50FHG1QWFbbdM2ZtKa6PJg/FW
kdnxV01dwXFug08VLTrd+uZJEhN8I80tWuC4VW6iZ0ML7lbbDs+MJRQ0ue4I5fXsZPHvxSir5wmI
pSqc4QDMf0qy9EIiRZdFmpBvGDuORh+8Xk9kOQmTnVD9s+7Er0XCj3SCsU27KSg/HnLjIS5xDHrZ
ETmD9UZqxVl2/+BpeHsOYB2ElCxmkJGOB/jTQDNt10snXRA+qXAbXRFsMeylSqtrPkvV0TcLJPbC
4P+vDsVq9JTp7ijvgWqKO4Ht4Ry6d2d1IWNACLsHTK2kVmaJfDspH7mxuR58uTPQTmTa4uqjIs3g
P5ePyFhYTO2xZFwQhFu96hHjZRGBzftb7M47yuWyA6iv7bH8015zeEMdLB00OKqbNDwv8fRxBVaP
jghu/EPw3/YjSgjLyu1Ge9jEIj1uhf8ODcpnPDLputqHuXj6TrKSyZU8In6u6yGs8thC0gd6VGhN
e0U/kFaZNBDmnzDCrxPqAbQVtNKQ1CjqSuebP0Z+j5cOurRVWh+sseIb9tM5yUi6zXYH6dIhKwTZ
V+Evf+F2CdNhU4YmEqdvTJw7GfQuwJUPGe6ag9pAbVavIEVrIYP6sgp6vag4K8KXmxZDZ5E6/Oky
u4qIEYE4emVd0ikqxm6Wt4Tck9onYavGKibwft0bBVQB6kF4Os4CO6pU/5q4uTUR117Mjjcoympb
THp+gVYJhQEHzgwhufPZhSD+ckgklFWhW64putpx6l6OUtB5UhY9WX5DXvgOgd5o/qlJ9fTVS8z9
fk1pYIz7f/mF35AlEyrTOJx9+xbk4DLz3qnO9aMXWjvvbjhQDyJ5XjZ0aNL/MdonEcI0VAirB3fi
z7soTud2F7i1RIPpyZRezDUDusqTpX34649cREYDD+fc10rbI62NRFj04P6ojXq64LYMdgtUp/mC
duVgBfmOANPwIQI2P7xMVn30bKngZ6X+HB8/y9hiXi88glkGMGBhKLCcV+WpHJxTESY6q6RTkSMK
pv6Kk83mtylW90gCBTBtU1j1/44UK2U0nO0IIvFMy8tAOJm/m2s3Wmc8AsRlgUdCAzwZ9UN4tsds
6zDD73IRqdCvHdhgjcecXD6R/eNErDP56QUSo9VXpA7joy6UGkFX7qakQTdLBHRtHaHNoVL3OQB8
pGYgFA6BqQS41isJKV+I/we6glSGHnX1PHSYaLF1/e3e1Z9LgqMgKjHnzkdMe8jRLpca+jUvb7Af
3Hdyh4ndJi1U1YTaTIoF2oUi7m0tMI9oCvTQa2ig1KJYvFlcoBJvAwNgyZWATeATMkzsXly2zRhW
Yol2xSPl+4JspPthCVf7Se1zIifgkNkTrcNK/CrhqStsYaDiNLwnfqTc7qVOI0HpIxwB3XgQI97h
g1WxZx5iWBLVglYtYPbaguXVm9cSVc0Jh2UzyNyUWBG6vDEpbxuDPek7HUcnb0RgCagM8MRTk4JR
uLJIXuUecVJpFCnrg8mjSsXv4rVlIvHbWPAc3ixFfRBKg+UIV0utrhx/+H9N/Qiryyk2Gkt8u3jv
yU+pzXTKg4ZO4zeE825d1odEa0bXXRxqdKHQ5fU68aSNsHEjzfDPVn4RayWVfD1S9zPi0zsqzWVS
8GKvTAibN+4b9QETbURTxkwXCFvV8SLhlP1t8AFJkR/AgQjRuHnN1PnHy3EQHpeW0qANEhMtPcfz
rDT6zvBn41H3N/j47FJPJCM6R85EE3VYbJBN3GYEF3HTZIS+emFjJD98fkVQDUD7f1feCyrCr3dr
OHCowOcnS70NzYkUbCxS7PEcquywmrNMq9d/kT3kuwSnmqsUmo5df4YbtbihXioq3Y3fLX/mliZu
VGD1gd3l6cTvYxbjT41wz6dn4x7v5+MEOZny4s98f4aXMhkOGIqpbadPWhdku8YloBIgMYMkjSLw
db291sheJb2rKfkm7HDsoXo3x3RwVlAlP6EmTr6AALH3+eH8MiwHLS+d5mnA4+XnEQtVC27xIk0Q
2NBYOdo0yYsheiByHiPuWiEsJKXhkNErjac01wcMmiHOQcT0N1tnoxoK8qIJk16VDmdAuOY4iKKZ
lgLFfKIz0LcicXrfoW7jxq2NmzI5EX+Jy/l5+84Ixo6ce2FFrZRByul0BM739C0ZmwaVDm1kkn/+
cnoO7gL+AQkFP1L/ByeCnAXy5SFkNdmpe/0fzRnnHilO5dME3L4Ez/+KpFvdqd6bMXuTCNHSFfIJ
4sRwyBJhIBkyysdSdrvroei8hLXz0IfSYpC3gyxVH0DwYZXnn9gzlhtcUx5p/2UaUkdU5fXqSJAG
8Cd4vM6eoWZOq6uHhF2/7JEyNqaQuhInlunXI/orlLCeRT+zO3ztzm5djATKKKJRnVsXhoTZKuVX
GhGacWyrMNmboUf264Pww/B5dyxVCSqU8KELNcYIiNFILjAosxAnr/ihezOMoRmP2o1OIEG2PdOa
VaT96h/HcU2tApwHRcEoMJJYTeiEZGgQ2Z4dBMNxZD+qBw36d/k86pDKzql0kphIpidCMK3KoLX7
YoRAwRDpM4pWe1OkxirZftUrvUqa2XLT+foEvuYajwl2MBWzmDxfqyEJmV20bI7dpaoxONfSmyKI
HfsTj/ygwaaTNxaNG8UzgAQ5ki3DzvPmudFPe5R4LHEgX07Cn+ucF/+U7KP9GmfV/S/dZzNyFCL9
8msS+LpBBj71ufgrdG9tQbKbZWjJIySa2GYUgG4vnfckGNo6ne5eOTXO/HcwiuHb7QJoCOzYV/Xh
pGPXBD1Baiy46Qmv6ELkXlAmDB8lj2SxnqB8A8GR6fCqKGl4P9/RyBZ2eAAmgbk5Ljy8LgqaVlYW
ZrWCDdXYYjEqwBwjDEFxXPeMeGS/+f96F9qSow685S51ohJxTuQpBB91BhEOkrb4ct9YeQDYfdX3
xqEjnf+KhFGPELhYMy9fdQ+RPdktyJOI1XKNPCPlvR578+Vk399lVCh3aMrylEWSnqqH1G/919Ys
irXQd//csKINi0Q3T/hvkVM2PRMKtBaczlXpIxsSh4ljN8kYC+dxaCFwEgLiP7/8C2nqHO2qdBPG
f4A02z6iyIQz0TECwSKNfkkQ12ZReJImp7mFZsI7iN9eRl87H0FKsAZT9LK2QLna8mN6WklQE/BX
S6Id9IiEbtr8ksC+FS3+kQLAU5DjYHX7/nIxQu/wkRtYrx+WKl5ZdxcOqiPux/iaiQZp6K40Tbe0
gXV/PwpgnFd0LC85ADRL9ocZJMWun2UHlkCOneAJOxYZGp+c7Ni8WTStCLieEvQdZE6mY/eMs2Vq
/T3n+mwryIdmFpNWF8wiAyf5Al2QEQE8TOtE+AodB2lwb66OQXQNDKO/F3hhhTZ8bXt+8hz6Zo4v
/iRoH5qCMRs1qf+2WTRVvTqmfrnALOPs+9EeQKtkOZCQsbDvmWELA7GCCCThitrBctk+QT2Ru4VB
SaPYrC1QoSr07UxDLduUyrySY81slYoLd+opKAlMSffpErYfCpYl3OFnic4tZt0evOnZ0qk/kkl5
BJne0a//YhQYGhq9Dx9KzzmuxZF6ch9Swom6AvsO62JPD+2YI+av0GmCZtOAAl6shSyc/tUX7J2j
/JjTvNve8mQiIJH0NnWCbf//JMHBIyCuEQLOfMpeRRI9o9XPupvrHTR7G/oGsFqgm3DzrtpJhbqP
lm13o+PHaGP8FQClJFkV2q6zRc6i2ya6NXRSaMf0IOVle+38Xd3JmS+7eBaESx2dt23Ok9aBu/B5
/pNSGiqYkQVUarHTVtvaS1eYZ5WmnLTpmQA2Xj1sgQImUq1yw1ZSXx0pvXYYMrg+aoCxtaAwqx0n
CTmsjl8NyjNanKYRF/+lJbbqhdH9RGvDgt5Rgr4T/sF64ldtwqltohjYPh7QeiW6EcbsTqLrUSUR
fE4vZRyBCeXWslGh/L18lKNrwvP7tBdtah1GeQIv0kdSIiSfVhdu9+Yenux6DiWI4tVcsR+Mixnm
DyW95fvwxPz6fyHBHr3j/rXwZpBAo5pjunUS2tPi54gv398ZVBp2EVnxf0Hen5NtVaaC0e14j3pW
2ljLTURtaf/VIe3d0/7Xgg3DJoNxpJBHbxPiylUFu4D1RyPCqWsglcS45MahEKgn73wAaF0jzfg3
xDU33iXork3HNc2o16dV4och4y5tOwAHyryDpSRHZELT79tdlZwKSqL5cNT/U46pilCE95qODcac
xi/KxmJzF/xbkBRxYSlUrZTZnbCoTdBigb/ixuY8phUQdkl241Gqg8Jp3upSv3eq9EQhSgcTpdwt
Re6a+bCfpfrFhqzJjmL5B4hdjLC+RYGOK92McCvKJWkUM/9IIwvxJaQVB28jY2cshjvpMntFyxiu
jjXRiJ8GmCl4iw65eyMdzPESpGxmSNO6tHewZ0ELFYAVxlfibt6prQaIixuyB387oQRlJqgAGZ1S
3T7hN1+V27PWUCbDIg7gIm7oCpve7xsmcmXljQoE++NAmG/UFKcGKKWy2AdiYSXYpVPcwCc2QS3X
3Il1Qh68JqotyuXXVLR5GfU827hw97b0UUym1nm5tVMz3gSK/JgWJw5k+uOU1v/6jxW8sCnYoAPy
LjL9tHhFUrzGFi6qvHKU9i3ncrAlz2MDnsJ0aEzVXLjaKXggf1xS5Zm+GshVuKpAOczb6+Bxi3kG
m1355XKBX9Lxj7AK8exml4Jmm1mk0Y5uspU4Bg5IcBFHdY1ze27v5Bh2IiZe4evnhtdvvAiWmc5X
z0I7t66v26QRFVLyu0rCqlu2PEkHZKbqZryMPDY14krPoxc/GnpDv6Y80yUUtKOyKjK3x7DKz/RV
nT8SGOC1+B3bAmtXXnBb5QX7wwAtgfXyD1RDOeUb60aNnub5+lRxtFRmo9yPtObjLOSW8WlMcia+
sITw7rqbel+056i5Fl6Ps2o91VoshX1A4Rp+Ckjc3zZvCGvl4HLpbnenzEv6h8cYTHsyhjN6ptJ1
zzRTN2nQ99Hk8gypOvZpQVkB0O2t4OZE/86s/eq/2LSUHYWTmTALPzjeu3nMWMalDoegwtG/JqrF
umND5V0QX9VtjO3WX/lSR6nvILuJYakyA6tQTePnT9dErqvf/i1CdgXzYGaNIQBQYcx3dvrnpncD
+81h7bB7KU6xT9PiiOLFvHYu3h4hVDoGdNepxqng6VeW+RJQRhgWE3bxIJCncmYlM0uQAY5YBIRA
oW5BBQj7dtB9PGMu9BwN3yw+r432nrGGZJI5vsopvQJNxlYWKDsLMO8y4Uj4qVtsqvRO+rWta5Ac
iaHw69LTj8uE5ZEOb81uOSVQzJk+H7RjK+SAbEHy+Cr09+F+VDBXjY2VXDfgQtqPNtOBZgUc0dKl
UbAUptvZfveT11breNLHnixGlW3SSk1rDCLZJ+wr8h9es9vENGN2/1bgGetMbZqaTN8BFAYi1WW5
fbs9eoZFM3VdCbb2/F1SGO1rp+k82Q6P76ed+dLC34hLO/p3qCzgM2BvGw/IZB4VXu+s8wiGjAN2
v810cFUDH/peLy3WKn1rOldrKt9LC7PX4tnknSh/1f/xYf9cc05M5PjVi8CnpyGNQD5OP8L8Jjai
+uF/yD4SSaqN0XeBoPDUSlbzfhSv02CIyvxOW56yL89aGvknLxijEC0NiPLfBODqgwu703c31/VK
Jiyfx2NffUwvTS2+E9J4QoVK5+6+rCcML14Clolma+ejbtUKEVL7vyeyfIg+IVC9U05kJzjMhPOl
l3+PLyu81R+LPAlxAjE/msKrQYmWfiuyp9Hehn5MzNzZhbcB0cYQmWvvUt/vDIlMFAxQUH7v3aN4
Tmr+IxuVyWAv2HLSG9zS6bXWlWKHeHx8gSvX316e+DiJmIDHxLrXlwKuT41Ur9QAOVw39OCWpiVR
KhDpBqmC68dSakZdQYDKw1APfyzBUWoihlggtMX7xwvF5qZ0reScferBochbvVpawFmOc33ubKO4
w0TVa6TFLY9HUrTUG4cgM5hEe81hp5fnmx2F/oee8XypyveY2RPH50zfu2JsAyPVAwSmBRxYUm71
Xyix6rxyioP3P8yj1qMudL2FZgxDpp6yyX6ZTWu4+PIEHT/NdtHDbrH5GbkJnm5o4HX1uCYi+Nub
NYVkIyxy7JLeL6SpvSNev55VCJyTULrMd1I/TMA5aDf+/m9Fjs40gQSwfWnJIuspid76h1NNBqTv
7QOd2GsVw6SvWmrhOwcblyozi50c4s2WxgUzVjeI9YioNl4PCjYWzTRNOAAbWVEwBuf+Tckp1jSd
eeZ1YGJ/D6gwjNZeC1F0owzs0KBfThhIPYvuHUB5d7tL55QMA953lHyGOd6TAmfcSwCsBvhtlKbR
A6ixMXdZphCA5JtL4S94VmXVWVas5P2rqiGT7w/HlLqUyq0wOAAloE8N3IwRqrwtBSELMVAQxvM9
4diAqCVqLNG7W6VklscPephW3MClrbwGAojRlVXj0K68FFUsHx+2yeBjyRPp1ACaWLxtZPlVdXWy
BDfLd+JQsJE/e2uk0m01d0RMJ6e/ggKT8XI5dODPhWCtvuHRpxBN793inJ14Vbz3oDuEixbXvMlX
LnG/F6nwwHtwlFZd0l9kp/8/QYsgc83c6hWPFGccvZbGLkeDsghcESP+cD4a2mW3NUbYFv1WCiw1
yptp/lM+k1wPI6PFCsF6XRK1yneh8dLFE+iBfndcu2hqKUUCdUDvrCuHHf/79Gsdyntf6g7YfMAi
jy71HDPdoNytnwUbI/zaHd1OqMV1DaJiblZgFyBEO3ynsvTD+I3opyYZcVC5YcEfBVNsRZrJY+Ai
fJYP+Fez5gmClct/mNiH+UGjtJNTPB4BYs1I+VyPCpaSWFxOtZvBeh9kfBHQCozV30O+m/DI/fK6
NEwP+hSd3sIam9a8kQC/STsSxuwbo7vaqpIjBLdaojfwHfNKHKf/du4KBpIf8zDHJlccPGitW3f6
CTWzewrBWs/UkYUx93r7s7dei/14dT5buKbj4c0YT6yLsYvb0nbkP7CZCIrdRTrQX+3+/ZCDD1lp
daNI+eUOsQa8st3jcV2Et2QbItKE4iTpaAY5CGnWCCAEHqSI9W0UTEJyGdgI6yyJqGx44F4sUfBf
29ADPJP4O9XwIHdk9dNXvVsu7ClcRtrHthdwNtjrWe5v+eUAyg32uWxbx2fRktAnZjtkUNXnPfLu
221vIdeLAFqbNDDPS4uaB4+XYfPIFrqihz/i+JplLJFys//ge+ey3k5fT9mx85QquVDMuikv8tEz
eIogaoi0S3mGd9vaIbDcGsRKCBMQNcNhoUp9B6uxaHADNLWZcc5q8wMJXFCqKtm5ZVju3bpWHWKP
6pvKbzGxBZ/DXLK4FKseRClbwm/9hbm8pIlS28527eLBDi8XbK9iJpTDBOfmr+J8FKmHg8AdQCoh
n/tC3so6iB7kvpCjr2v2A6RJqdqeVMUh8s29ZL4XjOTUKuxrPndkEyjFT3sVQ2r/M35vK4pQ18a3
bh7MMH38CmUKLluR/0xbp12OaxaDqEpKCgtQfBT6HE/XCuikkG61sVUXqBlRTld+qhUlxgsCrlyh
hzteKDFkay+l37sa5CKf1c6vi6x83qgdtEqTPgj2NLGuTy0AiyXn6NVaAukfeB8SXGmtfzmpd4Ts
D3QVg2Cl2QcWhq8lwSnbwRK8UbBgY9844Y6J/q2cYd06QpdQcuhDpHaZhQ6NO8TkLnFlV32v9ZTF
JIULwVrWTa4A1L4FCB//8Dl3Tin8269hCKX8CYZtQKMrBCwkBeY6syN/StaISH2n8Uw6dsN353Cx
pnFxNAj5CXnPJFf0WY5uUdDEQKhOEcMr48JAhw4teErLiU/AtTb3H24T6+rXNoNU26a/IaXrp2ny
aS/jsit/R82bpiwrNrpjTtmBaO9S/nzKgob3VVIfJtN71o7avalpWGr3IXw6AakMeAOl1dfDIEB3
MNbRNSZp1k6FYLcYzrqZu+8UcenJsxytSIDXiB8vpoBSpKrY/x2xH9FFyl56O3lOdudVAGbuIf8r
pCn21DX3pjLtC2IoWv5OYbhXwaVjq5bhy+y/f6tyZbwHh6P8E2U7YFleHrIn6CnVZLObRbmvws51
fVVjOVopf4ZwfjbvY11xhDkGK6RrI39nfhwbOybSaRJy9HZ3ygrangYrndXSNyXXNTJ/ppCrAuOu
H36ICrULbxas4ddL80VwOc1+C/iDHPmsyAKSX1NqaFhQrR4KwcavpTReViQPcsgIrXOFNgzcTCCa
ntvxgC3ZxWwsvWWcFLnIr4JHzi7Pp14B+zbV+oPB24/4b4BewgglOCiReDt0vPB6TJAIlLp4RWrk
gpRPpIR95/S8RSCkoZRgPUM0ijm3w+0DuqJBSwnnS8tT6JHg+z3nNVLNkxR1l/B9QnqCJ/Djgu5I
BtPpaw83HKI9+948uWp8W12YxqUenssJ8YfDC6bVgYUaMf1wpZM0gI7+CyiukUYmB7YpHpnWoOFd
BHk1PFuTult0ixNlv02O7oYOG7MVbotW3kNA8ZmhX3hlwi1XjzdMmJ+Sf+XorTwxRPskr707S+oD
z8M7EFuj4yEnK8VOIQ4Y5MrC+DQMStEpYinhylpHBtS+LnExHoaXbmcIz9IOwT6WGyPscZfTnlBF
xwNir9Ukn1Ann58SskmHtkH7Bcc1OptrbUlwh2s0+VZC28NgVAkgbpQaLZ+8AMGWyBvSC8Ut7AAF
sXk/PxnKjjsJ/fVYRSstNUcv0aad8OXBoanO9F++mL8jIhoAFK7im8j9JVaaFIwMRg3oh57oNeo9
Qb7imusAoI6UIhn368TCzV/R0W7W2F/RsOwJxbNmTSPJeuRm82Nos+3BhcTQQadY1JkIumdkDQ2F
8H/PSpv02Q4GMQcKKC5UpN2VxAkIYBa+yLGyHfa94USYHcpVarg9y0er1Lwa9n7XSgCV47mHP+7v
EQ+kjEmvZDXegPjn345VTnwzX/yjlOjHKcTmyFeqrj5gohvaoMtWbGPWf6wxlfOoNkKVyLlLcqgP
6ZaZz2/jsBjakncNrTVUKFXlsklwblMKq6X+WELd2Ao+dzlbvDxZSiCy3XMn8nWqxEGfOajgnDqM
0MAUuqbvGEvtxDDS629s6dDGwrxhbXzdoBidy2QbTz8ledgMA8NQ3Xkrc78f1zfRd+lNaUJn+s2a
A3PQu3+rveClGn7Ji5DQhS5kkWdlpTTIg5lgXUEuWCrE5FqBow4O+EfzOSIo4pGiwj+LHoyLxr6c
G5EFr8Waf5/bfb4egy8X1FFhw7pR9p9fXAxTOavMJRZ6uzQvnDdiah7/+fP8kTnx4dj1Hr2Nb5wB
V2/+amAoKEkwJn88tIkzzvJLC79+pbmgBLcjb2xqrywhHHzh66xKoTR5Mdr+VDpSMzm7moLDjKp2
SVM9I/63fIh/0KVum4+TRr/JCSiL0pgN5926WKHJB5RZ5cMtpfAivLnW4s1yzJCkjzf4WfT6/puN
QDKMrwkhEc119AEW+TPAEdaXr60S/Z9/YsdoQihEqbuXivhc6NhcGfCMmy54QW99UDsYRwXfpdux
CUNdvZSxctEwVtQgBkIUHdAss6zh+SlMinSqOuIDxqdAQfXXGsR2+NBZjAUSM8uXRwfqHMzyAjeG
zXMVOyYlWLwMCNnCOxvYnyQkuK4h7fRxviMqJps1lSjLF4jF3sjOiZHfNk5OiEmlN9SjTkD6MgmU
aTWzaDJLZQaPF3svyJ31PESJIQRTICkfp2/2iq3+uqn4bmnLHkGcmZmoS9G3fbt5OV+EG4MxKFhp
JRg27+92JjE6Jy7EXUT+UFvVBhawF4kEZ+qP1OHu7LKGXfK5gAu1CghCzg8oVJP7HPsQImAwpLWr
XmhjrcmeRULHx5nwF6Hh8XuALTW46/g4vozrjeA1VPKfBKCXmMUnt+g3GO1C98/c9sjsfg4fbqz5
u6IzaPqCPMQLQBy7jQuo0XjiJZPPycQrBz+CQ/9lTwzrWZdLa4ikl7w9JW7nJ/AaKyFgLX1jQ+X6
3MJDEIiG3nPYPdar3QtgAgYoWUx6HSCT2eaCmi00Om3o3DLj0vUi5eJETOiEDrRjDcPUSnd3U5R2
9M1sq6eHYkPjxkZvNJ9LnP+tPZEFKHPzcwP8NO5wXf5CcgC+B+liUQTUrh3amNEZs9JhI+GCCtem
BODZ7t4THIoNlLRqxkCz3Mz8ArmMAKVWQyeUZvcUc4vUorVYBa4ZKh+lBGNzhYGl6WLt41cCVK+q
B1Sx9wKh3lPLfQVfm5AuI5OABgao+RpCUJg+Smsy5EqDHvxlK6QceB9/L2NxxqpXEZyWhEBK2PFE
pkLDFAdhk8ujAt2y9qcB2hQKKBOZo4pWbu2p+ObnSAYOMC3w8XxTxcD727ty966+zw3FpraYNHO9
VS9y6yGCDfKdVb3V+rcvrc3V9dEKEigNSUxby5Cxe1tpIsAFw7ZZyhlYOGymyJDn5WBiLNqoOEMF
BHx6+KW8wjUwg9EuAGe5vw6/WXM6bav6Q1CsLMJGTbr1Rtw/ayYGE7bkNQN/EVSO2dQIX76d+14E
HKpl4jTZo+YhmNZrleofwOvphmdFyW0TcOCH6FZUM0QjHZGCwyCMJeAwI8SBBrnVWh00Cihe/eOM
Yu0i8Pde0Nb/yNkhgFmnvf5N00uQ/fuZqKVrXc04aTs/bdM2QG0UwKcNy8yi6EwQCZjGyztoQiOg
UsJRAJNPXYoPFrDAWTXhlgUBohcis/Oam5X9+1aaVoNMzD4iTErN67i6joRI1F7tLgIm+SIR8HKD
le3P0dTOoFd0Lose8fxpRvt+goEqpLUw6tDyLEnxUmccI2pSFHnJO2JKwhN5Vvp25uflMA88UXNC
ZsFtVRwb/row5VbHCVL9xO998uLYX8mZperH53g1BO/c/zkO1CAgksjsz4zCPOqMefwpvf1pSMnB
6b0cMqhdRpbpkGQXdTrdR6uSd9LqV25UICAFuo58N/29MoPN97Kjr8nQ2VwGLljN5z5RB1XeObYx
5arCPz74wodNH5SOrS4lnXjJ1Ky88ekApN7xqUSYOLs4UKlqPNA3xeP04mZilEh3J/GsevfYHfH8
pnnH0YNPg/FdN12sZ6TRF1apaGgMhYdXztz+QJNqXkJ+Q2y2+yIXo5wvhv8cQxYEs7WerEz4LNMY
udsXAW0ycA2uHu0513QMZupIAP4ezh7DQV974oU8bVasIG42g4mnT+25O7Lp0J+JLaqUBBt3r2aG
SWHoZ1rE/NTEnJFD2Lbq+wxXsHm9nMddXR9ccRVeRJCrEdJsQhlJRRwj0Y6Mx65Y39DEQwa38dZy
VISO5aXweT4Frqn1bYolx7q2FmG1H/trgInz6ONzkdvnEiVyEvvl6NGU+IYFGaXU/SmqsI9FUanR
vprHyA+uSzDRxpRfAHKcGU21d7TIVA5AYDgn7snbg24Rj7CG5IJY2+ReAeDFI3yRpHThSpjeDM6i
8I8RajDJEpCL5bbEosLI2w1L5lS8eBw7YMsK8/2LUYrBZ5N5FGVBV2BLNW6e4ccQaeAUcoDDnclO
igFgPdH+iBgPUCqJeiFvNnM9XAeBsVC3I6RjJ3e/BdS/yQnG76GkrKm0p3VeT7R6nWpJktTSph+s
jH9Zl5/+vB+1+ANYQfKexXiFgHBR9xqa68+Keg7fqRUIEz49jsunoMiIBk+89g5lF6ohucG7ak+H
gW8AqJlTK3Ib2P4SIRNuCcl3UYry2AbEGvZSLPu35JEVyIGv4OzaztXSYAIV+vQnWKdukikuiGHS
+7K3cjrjtxdoh2aAjU4g/rxliaLtljmRHoH4iuSN9VSJ2lRHuuCoIAPwT6NRRu5fHvFUT28IN1ZK
F9a5XSjSTJXCy+AbLSlV2uQTZo5nARqB04rdiritpveajXIDW1wFhhGWMFMbLlTJDfKsJi0JPMHK
91IeVMrCoTzgbIx35R1U7NKEiNxi27PDoyJRQzgiivfLVQ9EySHP4CeTM3vrqsN9dlq72JEV/Yvr
yG8aL0Symqx7u1Va2YKqLpKaHf9/E0DqF7L4wbdMADY4aOxUUtY2DVcUsYeVfcVYGq1L5jG9KUfI
rrpSEi/tGXRRka3tQfyGKaYQrRbSBj+Sz4msBS+x4EpWbqtMBBzjXy3ZKyexs8PvEjFAK4WwiaC/
o0Uwauc0oimdw1UYiRks19gSru6pGF1VlgTS8OTGnobLUcfU5wYSeK431iI8iU+xvqwfc+ViLqFn
edZ6/8NwT+wZ9amVi8DAawjJzElXu7Np2Y5UNs7nYlzEYldWo/YpUHm9svsIylvoBIai7X7JX0FW
ggaz4Qc9WwXxZRIswbwdXitoa5pox5f9d5CSmkUf7INsrpfkqQXWLHiFoPfH1UQhYuDW9OmP22NT
pfQgVEofAhV+GGxXDrDG5ZO2/r/8BuyYZI31p7VDhh/3SazSxNGC1ufmrNyeYigLm9A3xkllyzia
A2o8RyGBCqXnu+cXU5V0ypoDS7/Xcqn0ROpyaM7EiYpngbDrIeehxcgtr0s+NJxmIMiv+amAobZd
3LkqJ29RmnWwFxp/9yXtzQJKR3X2Y8zNmKCNPNndV0My+xTu+S7Cjc/MHpNoVPRUgUP65z4lI11q
PdsNI+HQol4zGAhRNUas9wPiwWGZOOeX2omCXx1HIZFmDr++lkUE6sPFvNS3m+2s4+L/5zJSQLQ1
FHaYKHrrloru5stnTOZMrXZE5fgIO3v9uGKdxo9n0BqA+rzE0xJOPufwJ52Qz4u0mT0idi71pqUk
XWCPq425P0xIhGeKC30NYXGEJZC32SoD9HAkB762FytgFzuwPfUKPmwlUjYQgMSmw0wROfOE0wsl
GCLrqXA08yoonzrJE2LiAWIycLKX5j+qfw0uAZiZ6Xd0NEewTuWWcg/0XEnHOd/HGzSus5Q3/tey
sXxIqCt2c3gyIGc+K4PPfJf5Ro2MgamMDnZwoW8E140q7dzAh6f6DJ1aSvPGr4mZyNChjDQfJcE1
7ZtfkKVAcoPeLVEMP0a6OucIabkcbC19hCKGSts1Ip3T/TLTUGGjrYXk5ku310ShpTIOy2fAc2ho
0TeA8fNviK9VUuz/hpz7DX+TiTh6d6V4DMHAKtZ0PmO3V/0jJ7MM2vPSxA5Xu7CNx2H78wfuJHLi
GUG10yXYqAFlV4V6Va+ygL5kEigaiBbLHxdzq0hnBKEskXn3S4uXSXYERhR1dnJ68QDeV3g+4WGz
l53MRtZTHvdO5uYVqH5ElEt0anofrtsOcLxrJlSue3AJYtdh6bQUPf/Owpp+7uYY+5pHn7sgjNXp
BlwyyI0kxlWc3cyt/dtMDu+XFADAnazE3qz6SdUqs2ZU525PJUm1Zo02igT8yz8bRVoSxUaEOLg8
Xy0qsmmMjfYLvu7TN9RbX/6tDOVIKy2nhaHn/3IYoo9XKxZRP7Y+pQaW3lmrXKUBTE3zrz5gk2N8
fYpH8BYf0Njz17DKr9uo7tFjXM1LvNavhUSr7DRUIRG/RUjhiVK5NSaR+13u14lylN3mtiRWWD+0
Mi6PkQi6988Ov6CT1Vi/a0x/ugme+Ejuzu/clQTRRpCEvU2oMlEQV2jByyOkjVbgVG1NxHqajeb1
cUBYGIACIr9qRO20Fmb9ieoONrje/575s+2+cF3BBF3pdLk5s1o9DFKCBOelm9Vcl04nJ4/TDMkN
Lmlw+KBBocHn5dRrIzQO3Zla6ErG5WzRzfpIDxYsnf5pqWG+e9QS1ARr7udL/uOZawMi1vEEeCcT
cl41pTzgBMGN1wjfz7ok7xVtu5ra68kgmdy4uVsZ7L4+2j4rHZHZbXB24CxB9dNeSy2AasuwOAtF
O77Ymo64r6lUMJGpogYT7KyUSHwdOthu19pxmaneZ5CdNNccjWNC3RMvjSnIq6t2UXr2ogDJxj3v
04IIgfCyP6U9cSSbn9bjJB5NRRPoi2wj2UzHFoKKIDe1pN3IrgONuGyCEg4mOM1vFJW7gfK6QrG5
QRv/FfqHM2ETDHnqgFncjR04SuCmI7PnpwT30A9XtWgDBqKh46Yv9q71/KZmxV73W7/8+fTDuuwa
XPWRrY4oRX14XoXVe/Qo2lQDved7Ovxx6x/to5NfgtEJUJ66jWJHv1cDSWUHfW4oddQHDgB9470Y
b7MOcoJqAcSvOGw8lSxqhJoIX2Sn+f8WT5Q5B10feid/WVq1pZmKm83u1a6SDadWwoRj88mEzXJA
ZdAJGVJ5f5J/n6FkgnUvC1hxIiRLc5z5YcP+/MGYn+z/IoTZz3NWK6jAFG4fJvXhmAX3QhJYVNnG
FoQQG+MatA8tuuIPbce4UJp6cmo6FoNGzw0btm3uRk0wNC2gfXbR69WHkpsm2vclyahyTdWbJ6Nb
m2GRPLeBRANrrRArcM4pEkhYgu4UETteUkrDZC1YACS+ud1nq+sdoL+LeRAp1x6jXLXPxRaCZtUC
baqD1xeRJbPMamwzm5H+aXrDZQgLTW7z12IfqzVjm9QURLLPsc/MU74jsQkLZuRWlHC/KgaZzMmq
ALaZqg763StyLbxudfbrvOv0QUwGoP2KQbacfsDXhwBxl06mBMgSDDL1U28tdTG3WS1DWASyxHQ/
qHkMgCvE2Qak1tGs6YrEaCmOJBIfcRUYf31j5vvclG0fexTpe8XAV6jTuS+3EvLKtscUi0pVaBEO
cD0k8fIzdY5SslziKIg5fjQ9tGD0I4y+mSUjWRH/8xbYzo6mZC2RT4YzM7sgxccmhh0PRHme7JQc
gOfllhemlaplV+CSSNunIuRe/w9FkAqxxDGgFiboM0EMqNt+uI5V9d8xmPgb1dJpAMXeM8EFytKN
dmoa0nuVsKAWKsWaCMm2lFJPxGjvXj0hhhfuhLTgaLfDpT0bdDGDDZlxkyWtuXG8OHjR5IpPU4vS
rz3wloM9co618HyE9bolUI5ETIYkWt9XEBlD9IU/oCZWFlkEa2UN67pa02wF3HKXunM8279/33EA
KMvnywppI8y/rU3aJkYoaG1Kwfs9Nc4v+GfILgnksf0RKO27O9CsVx/hamCr0PbVFo8NJ3BqVKC7
ZTKNNPm/5Yz0J8k+iDCBjTKuNmZJHutpu/1dPJ91N7x5Ci4mrSxxrmqelUHMS6a/NA+pFmvFTNnH
4Xqui+a6zGg/eW4a8cY5qQB1CM8FVwkazE/LlMPNUfFBzGe8YogX84RmeCEFfhWqw9+CHA8AZXlq
mmh2MFSflvd7VgyGjmv+p8bAOgC++EPK87OD9ltSy0JRsgrPszNJ30rQyxedKSBLNmBusP4JhsqX
mJnxEKSUvPaIwy2T9zY1XAB1f21LcI1Uh+f+ysgZYNdq3YU1/4WjwvVH7gOuScATLNSqCDLigfrC
WuqAm4BiEdYAEdrzUK2wzOb9fBIjNd8fktmw7hpEgbz9I4S8BN6rhuhB/i7/mW0y0eFu3dfVwirg
0yF1IITVSQeeUGEGsFNoJLZqkycyOarJYP1qcdd60m8wz/BvI9u1vsw1gwKtBwHCYvo4V0QxSrky
5PnpBclYnH3XhP4exAo3K86Fn7H5Ot0jR9J3eDXtrM7LyL9DFo8FHCC8LRSZJisOFvnvo7P6IirX
/338OHGYYrkVZgH+686JiQyMKh8KTBhacjc610euszEwZWveEd2FfTBCkL3VHWEx3OZKdx2ZWG8m
XfXEAEt1F5IavFo/inZdbfP1utZKkpv8ntBQniNcLg8fLOiFA6K2StmuZ/JcoaXu1mOxmS0P+F8C
Y363i2KaYkOip7/bt3h8gzyojf+4I+3FuIHbwwYIu7MZ6UYOfP4WZAzUAylxLgDUT8TKHSTFeJAx
JJo+aL9/Rd9ITaQb3t8BVEHHsOjQK8Q0dtJOw2AkKLfYdXQCizH3b8ezRH8xNMG17doHhu01kAuY
5y55w+xnfFvxSXTgN8xhu7ModiMd/MZNpntvgXY0V6LFIQjfAkbovtj4LZnRDyptsYO3eU0clj1A
NEuujUzEJDG5jrpu4twUTpV/y+5TeC0SXJMfIvFirv29XNYW54BTw5WJe9HgnQvtZdbSPIg2QIep
1KLfZHgqRvVLbKHFehaKWvky2WezSr7fyJ7w04Rtz8sYG22ZJcj7qGsemB6q/Of2CAvuXfA58mft
xigji1n38Er2be81ct/0Q+TV8MkODQa+CJZJ8AZw3pr6K76S3K4ZsJmybN9hM7X5vyv2MmfePJ6E
v+gCW3JYNa/XAWj51mz6c6zHtIlTOlZnyn8MupOsjWNZGHX7KYIUY0SWHpVe8pbYxTx+jMdSMP1y
MDsJjFZ8AXTCgh04RRhed6QajBcFvzMf/dQ4p2mn76ZpGJ5Ml4b8Q89SAieX3MqtOXDZcoUKKMO4
b5LCu3n3z1yv94PfCn4dqSaLipKORtYj+ewkgshJEXydYJ6zOgfzy3TIAh18ER8fVfPBx87hhk/X
QgdzFTllOWKUGwi0semuIFCbIxyOAgm4Jx6qPM66FNri7dbAj7djssPqUptqSzk6nThYuCxj0SQo
MNq+hC3HzP/fhBm8QpdzDpRa6+U0JBb8Wzzpl4YZpZ5l3CBAeIsW4R8w0w4On7zb0FHhdvaWcATe
xYVBa4EhHGV1D+rmeK32vfF8m2J4NQwZuJssTU6VU8gSas//20FioaUJtTCxvZEEc9N/nQHI/lS5
AnjmPvZxb8JAro1jPy4dkobsqV6jvA4MQ6vy5IJB7ctTLMmell4b2A3HVAUYIz+VLLA/AGx9pmVl
PrI3CjfKuWeZ7rS/I4ylOG0goUraEnLWXkkMKX/qMJ7qtcRKse0W5jlPgpR+gffkFE4sOOsPoBx+
CK8AsDEAnny5DqHRX+8hbuUsb3eXoXUi8jFF/3SRjHGIzHhLTI92FT3XjNSgCipdPNNaqwwriDpc
wf1JcKFKTZOZWbofKHZodOKYGcixLh8ve51BwUQcUrlLou9uM4pJrmKbazcs5FPPs/elsxxc6S3h
dWjESm9vbUA3Jckd+lA6FNmrqLInDhLhr4C7vXI+ySG6AreKSdj+Px/6f07Govu0Ri5eK0419Bzq
sA3iI6Zrkd03P0EOLiZ+SRycikxaQe9iRMjSDwsRjdcwhqX/sKKW0XKEH3BlAV6ZN09uTrqOk3Vi
70AbBawB0+4tV6De2uFhg5u6u+vSy/FoJTaalfx+GcAiAipwi8Llx7lNC35NZL6JCrleTrLrm0IL
4t/ieMAIl/ZJ/G/R6byN+bYUzx4pTFwQPd/+CCGx91wZFBz3Z6HXTuX0L5Zqv/0JvFCeByfEaKov
ek7Am0qH05DaCupWUsQyp5O0tOekGdgeW+2Iou26xobg3Tuj9xzO+GwKSaLw+qw22YrEXgNEweAF
Jyov7jVlcX0WnT23+9LWQNH/l6XUsjGw9R9IJzcPN5yeWwoJMdBkHGnvyDrf1m9NQWwyjINn7Z6D
HxwO4DN91u2tC2iy6CGJKaDDjB/JQM2I/36xp65JW7vGKmb/QulYTe8EVtNPFYUVLZvEln5a9CJF
KbxYeV54wEhx72XDKl2PfVJC9TSXVlwZJ7rWI13Vhw8M1FVrqjN54sqoa+90o0ARdCiNjVkHNwU1
2fwSg2PKIc79BpaGu36Ov4U53pt9t//0ujQyguifw8pyE1TR3+s8rthGy17GQi6uJj47RGcciRSi
6uuSCpSKLEJBEiR/lR8fGE9mFROe3DsfLeRLXEK6iHCOia1gpUlg05rKy1UXfW10zJn0tm5MIqwa
9oBNhj8Hvjng4cMk73EVZN9FMBLpFPP9pfk69+01m+4/FsAJrFdeH32dBPzWOrH8BS0ihAEDhHMD
99xWCTh8qvUrpiEgak6BIFbqweH4fOXXHZe2jZRl0n8fDXxY9Js2rdpbm4rHoLug4Wc2l/t5KLv5
ucKvinhFUXZDfaSijEG9imnqdktVzBOUfY90qf8x6IW3fdxjF+paiXH3R0fShm0P7nd2kteHmRgk
INHN3iUmAdyZLvH992ouzrCC0RSJiFqr1nL/ruvUdjjJUrAYkVfsiRes1wfPl2nW6ynDgRQ2MY5Z
aE4HIARjhb753+2ilQb7I3/Ozhzstjvcyie98V3IAUxiVTTbYhs1gR7jkWwJa9WQc9bY/cSxZg6X
VP0fGeefc/eD9fTB75hMdmh6ZeE4bn7yuw7IRf9b49msNN0By+elQqRGaQZ0/p0NxtZpLSK8Qlza
peNBtvm9RfWR3odMqSQ3MCT3UDXzfxOxECROw1wLt7aGfKaX5tkllMwNo/2TP5YnvQSdMPA90gcT
J/h7OvStRlTzmDyeIFdYFkjkUaLyUkzXdz37HMa3W2Iwaxg+7o1wSEmmCDNHl1FF0LFyx/Y3APgd
ylldgW3tEiCLm9fACUA2vbyN0sojSzjp0VPjIKCiC2wjEGTUxeLSB7HvgJ/a59RrKtNKOUrniuat
JrrlB4QAo3zyNKDKCClYoVSK7h4RS/CwyvrzerrriHOQNmH1cH7ZJrvmQerJsDniBrYreOuizKBm
CnwYStnxsSxM68Kbr6RfR2npAwAx2AmjormVqmhwumAZycXPnjqwowRaZGvIUN68ZE3OdnGS0wTt
Z1JUmomQ1upF0td79W0maAgAfvSFWCmTkslWy6XaNfO7fL80Jm29aB8XkS5iNZpWXLEHxdA19LlP
0JihCGwaFB+P3Si7BW6c1iOXx5hKtdP+7BQKsleus1VXl29gVGobs0p/yGgMQ0XGjw/UnfKHIzQK
GT3KhqpnHVFkBHI1pxSRLqDGZQf1Y0jKVkdpZfpJd2eH2Y2tB/rTsW06T3Uhqii4lccZKQcL025x
X1r1cIv0Um+mavCKzB2ps8wEUQZa/H1LIJHyXLCdFRHSATvxB6gnXHLigZsXkTjwboSauxmZdIkG
63aGkloS9QRjga+GlmJlettDA37OS55CKlW5Ngeplbw+Xh0y67IPL5tr+cmIhHzh1Zbsr1HKHILe
cz7NgQl3oJo/gMBskO6W91kmN8bhsipbmF2vJvNMZ2W5BnEq2RcnL6dVExIf2nNePMycwZwiF/RV
J+xk1nw2Nd4PocFsxAJ4ixRr0hTOLkR8h65OPqathp5/hUF+pcdjWN8Ll6GE+t7Z75Fv5So2ZoC4
SqeakA8dqY5neKPbvxqFj4O6h/N29HhHzV6If/MTkNqVlFo0WIob54D33VnmP+nEkrlTFwPTDz3d
CKlOcbNzFuz8rHNi+RRtg4TZsgq8uRj42fIoN0ZZ8xcPUIVQvPkA28oCZMOGbLX5yxO2D325e8bA
mqfl+DSFKkwUjR8g7TlMXZiezUJG1duhAytGJO0VkzEpBClQtn/8dAnpeCUCu71pFX93xy34ICl+
F10DullqwEBqmbIx0q5/AaoMh3IvsUU7SRCJlcrlJabxGqUqRrr5LvCUacpu0QLacYVD7m89BCaw
C4QS2mxqZGLuAHM5Xe2yA9aAyg4tKBylpTpDdE5G1WUCwlmSLCbU+BunSfJWozaXsvgvCO1trwWT
zD3JAFAml0xoFwRPNI74z/MxihetYcR2zJV1duDposuDjcTsQan2xB0FQJyjpgV9J83He2IwKQ7C
1kyvi98oX1XCD1LMs5scftiWVBLobPQkBvofI/xkfY90Jhib4z6c5eNcbqIZ91L5uEfPIVW6+iH8
bPmceWpgD4O6oBqcPcUBRpW9jbW1Vq1aByGAFJ4g87X5sCOUSvv9jerjhI2nyrEhmk1Ts1vT3rQe
c1a65iKkvUp3gm28zTvOOnAGyQPREQnPERJKR4Ws1HBzKdi2T0W3TnGLJF/yGMll9fpgMaWunPaa
c/xnDnPG3noHs5Y7BVs+8jGkJ8uByN19AYOrv5iuh/72dOLCXJwLXEJhxQOumOcDQvoBGLzJFXes
BGVqFP3aO1uCNb2KnRXbrx3dJS13WTgxVm474vfZjTMDgQ3TLo2awD5u3mFHV5UhMrgRqoz6iW8d
XnMzyjZ0qWFtpi7TjYPt/EUeUL0eiKx9GpZz/nmfOIWRVgkME08PnTGRZ4wc3pLx3D/QBdOnMv/U
JjtdY5CZLTO4FuZNoYY6XW6iA1ocPHaaGXUAigZGna1VlIWuipIGZ61txxB3ZtyjHgsaNGnVYTkD
WHJSf6KdY154GGxdxGyUBquDC8GlHtV5XUPbS1ikoU4B2dFw13B9VJwovrFFlXckABwCz50+/mro
4YZUCIIR2FM/rhXd9gMruRAndJpT52VKJRqFzu8XkEG6AKjFI5CCeOwnFMvFroBN9SOP5nwWTJFk
hSHaT4Ihj+dv4I1EJlgUV92pHsnd5tFQA88u4PljEglC99iulcKoVzoCyR7CSntKobOUC1304pT0
C57tPAP7jGDWSlifBZ0j9Z17M2DCa3lEwdTNmkSytj9+4BbE2a6X8qNFsHrObgw4f3ssP9J9xyab
sTs1TN5hbavidZuKGvEqIMbDyLSBZCzu21ULH9qbAn+tQFVcl6/3JTTXIMntlopXvx2xKx8ExxTy
5tWufx3VWN1yYMPbW48/HSy4EKGbbFPwzAoPP6RIfYTjkRxst87RdH+72wyIzI2nP4eFB4pH8JmP
9s/AC/bHZXuHCRAOI6hcE4c6idniW2eEzUmKtGOusUz+CrSO4GErDkMww0SJi9/bl0D1z1Cso1Hl
i/jzGlCIoQoVWJN+wQ/FSzU0zEFomxMRg/5fms0k/JRlQKkHv3KEkcqUntQylSdhz1HgV2ybZxSm
T86EsjM/95HtKzjC9h05RggWeEzDbDjqpriaNQDsDPxK5rrCLK0zvRbEXJsA2mldeo1DZm+4VDPr
JZKbsFdh/bvdrHkmFnDiqxBocsiTsoc8yT21MzHTTz5AJ6xL4WaBCCZscRPFf54B6cLj5TSF9oFV
e1MTRRocf5Y5BZYm26QL0hpoEVVj0Qdmvt24rOhKNWgWkeRNKV+Xn0WikNXlS9RpaFyY60xlBuT8
8RLaaG1BOpqUq9Ro8wTDk3swMlx0QgViB2IyhPVK48CC+S+dKHyAkY+nFPKMdQg2yIqpmBSXNMqP
0SwpYuNLwSnViW3wKW9R2vr1HpkrUO/2xet95/z2cv52uaBRAVV0HbMkbMOc8HVM6YgGnw7C4Ol2
XkWm74NmBCAjCXyyvOXDPqLjkM86XvAHm9HFvGVLHgU+/i7UDLFtFSdeFCdLdOlicXPmh0eqIxor
qgZeUeYkq6yjqRuTBn8YTzHrBj8Hf8Tf2lKPAuYwc+YiVLJNhFFd60dKbFGTG5uaDM/iodcpy1PI
tz3WRiOs88VNVaqQN29epDxvHdLbf4kdRTZcXKRaC3DNvNiFQXk3tKeYzrHBZuwtp1F3dDozg7e7
LbfHsai2nS7FA9Y97CS5uyOg2b9iTm3tC4p9R0MsDSt/ADR8rqJNfiy5qHLcXWzqX2pdVsnENdxT
WgSyFmCuIyBDbzVvmiouyzqIqI+Acs6e988bxD1wO5RsP1KFi9NnetPJNlIBh+Pa3HZ1h6PCvAxZ
Nb1GwhzRZ/vDobUdgDqDcNiDK0idbMzc/OiKpivRDZ57ZjYN051dBS/Mv/w0ExdthIfbBEEvaxhH
vSaSzQIv58pOw4d85njZOW3jTyi7xlXx9fY4hdK2AGhJlRxCiojWsMaZkZLNjvSXvMrkmQ61OE4n
0wVb+xCdki5IXh19rjOl2qdIG/LO2DXOcCDobVPKdEjArcD7vu2MR4j0pqUWEt+WhbJkWJhW5Pr8
XWPI6fdb61qlhokG2gLnv2sSUsB1NFLYj3UYyyKJWuXSaYzhBlg8DGPD9Ld5ujhrs9gbMD365S9O
tgt6f4Xw4hhzSjPeaAXbk55aBIa6s17tCiOtxsD4Gwci7PUBoIwDQvOQvQuk0K+DAZ/p+6+aWnWp
/G5yz8Hf4fuEgvKMCEnBGDzSyr5aTbKbvqKYtv/EeSXT/fQpMXKTAyusRDIj/VhI+ATaBO3o4lRO
1hZsaiRoRf4OItmWmhBYBPnSsJKjc8AYFsphT0mH2B/kPCgveh1mu28fjMluqlClebhV/UpAUhVN
xGA0hjYaEx0jBeR8zeU9iCFI7MUtbd2AWWA9K7zofH4yTzQEAYPfUwsO4rAxImkGlUs+2FWS2mnD
l5z0UzveFQSovQ8o2jOQL/OpurPNFeFHUoKGku0VyXQAw/eshX8aRMzFJs9NUao2EpjU2rd6dEhn
yN8UHyvbd29oP6bPdvnkCEybEXX8w0fPZg4PVTjopayxRHDoB7pMjLqReU7WkigDeO5nSg1u35IM
eRtT3muYxXi3GAsqk8PdF0WtI4w8MTPPG1qDsoDSNPUlYUpHw9GlIz0qH1ma21cPNJN0NfrJ3oPo
DIqQzKJ1xwnxuwixgqkWw3PdiQBUVKVtBwm3kQjIzPqj5sC8Oq7fcm66jFDu2JZbSd0qFWyPtz/t
HHEwnfxDF4K+zCGj3RRkYNlTCVn68VqNkHakqtO845T8bLj6XAgNetu/HPMA3LzQSRfp/jCNSdkR
c3LD2LG9mRULJx7INT+zk9hi6ZEiTc+EziNx/U4TKOC7xDzp6+IOUXnE7tdmJDsdADTUoD24IPOc
sHURtnl9TzIiXxWmAbDqpuOVqqdW3/HbL/bYPGegomOHQaLJymKeqv5zMem3m3pX/mp0vxRH8mp3
SAjBISF2szg5IOpxk61uOXozDM2pO6OR3Dp5oKPhFKTlso8BWQ3k8xUm1uJLBgxJTYFwLGkm6I7m
AGENR5EmORhk3W8Jdieebv9nrQPGCVZWkZx65DWAPVYLhEu4vwIse/qDmqAUmzwuQIwmjAGu9GlM
OZhyDEZuM2T/X8nllw6ptPZwVBTsnIyG7oxAPa6br/OY4GgR0otEueqPBIpYkJ4jbL0Ccjs97qaC
jrjSzgFADqtZTD1LQ6M2JUn55jJNL5Qyz8mclVyqQH/sd2Fl723F4B65dk7HFjC/YTeiBYcg5yCQ
7mBZ2QnNs3NOAfrjo3m5gCHHAE1jTOf15qh1iQ5W8EuoB9Z9DLX1RqQCyfh4uSQC7gj7ChopplLI
PJyG0l6UXwdeWxV/GYkYZtpJ7jA7k4megfA5nkGiO3RWrhdHmJ2ZPTSUOZTYJ7kq1DXHIJKy14Kx
QumzV5Nc15Z693OZaw9QP06pEZZrAfeyVxmG/xDtxsxw8kPnHwEmVkf2sKnmMtF0dNPiC9imYMKp
bC0/91917RiJwic+VvzCKSI+23PIi2nzGqtuMTBmJCKkyzpWADugdIHsBmB9pVIiVLJXazya4FF6
X7kcrfFjEkxIBEnTM8W6aPaNynfyawms3ljy6/E1l+insLq6aWaVJHfeqZs3UuEvoKpfDY51DtOW
z/8Noxt40QBe3WnrsQE3nuzTPg//3coQatBbafewAvhGlIp6qTTGs7ZtdxIfcsHnhdvybDQQWhJP
er7KlZX3Ms+eYoj4W31PDsU4IjQjTdaRKeGHGfrgWm+z22BgC+6A+uso1vvr8ykfreF7RDne6EBJ
3WPhFMjNBDSpBp5NQ06PzWNeQV4PUWcbpvlmFjcF3/EQleR0C8kpsf4WIbk7Grrzg+o/KhYYMN++
gmtRAO/3Q1Vjz5OfCtFkCJ8AKMxX35uKQPwPVEKtdqMowAPIBbWQYjEHE/PUXq2uiN0pn4Sj6Xcu
TTOQgU830d0dNe/wJnZkysqc8shAxhbaq1uUZ/42ryklOuIy4T+elCERae2+rJeWeKC2zl7RDOOh
hCsbMPVrX/bItJX6DQPxd0CGAlkziBDS4yF5S458/Jmhu1z+vY1M+JJ5LPmkDdSK0gakRIWasy+c
w/3uIAsW2rZjcP7spoWXK8shBpCi4zumzuDN3dopDkCv0n0igKVBNJYeBGPjdPHEYRSURVnF+OSW
qJ9hi/ub+TSvW1uGxlWOgdw/Jhe4va2dwj0k0renuZHIlErsbKlOAMk2QJZJPoJuh249JezLFzqc
euPAwBx+HEkaRK6Nz23gE2MupeCkI/G/uKEW7nKjnn7/eKPVo8QP4A/cjIHszZ49mcfG3fz4ZeXE
jKJ98Uir0gdU8peup+Uu2U0RVBR4EHaRemTVR2vPjcW3HKfymJvJzxuW0TDQBDNA6v9tJt7mISrM
pthZGDdT7ZEGNnU15dMSjS1dEQHekatnIfYmGN8F5QC+53HYkIvxXrq4EfueloeBjazRs+ui0M3u
93CAc0+2kVsh/9aeWyyY0hMLg5kdHCAhfkBigJ+ai8Hgx7FyWX6t01isj77PbFl6u48ZciUZpiOi
yQohCiTRN88GSld2Hm1sZl7c16f46DqU2QBaDsmdqUFWQpp670P/N4wbk+tP+DiQFr6GDwRpNTRk
1/kq89lNtPv6z/jZJLL4xGBRwZ3NvlI8ZQuSwYkHwJkOVTfJ7YUL9RXq/OP0lI2NZ25U4dOwR/i1
qFroTpfV1h00WWiPAz1Z5draoR7EV4NDpG0vD3mMKteS0qjQWNCzMXp5u2ixwYhxCGKhjNMHtXoi
DXYQojqv1n+5RU32WZ6zYCZ+Ld2ymj1nt8tPZ00Y2GiVnoH1zMCOIiWH3yJryVxmVuM8nzLKgmtC
7u+5Vo58zI8x5phjrkqFtGiTDIGgmUI0QVRrq7DoWygfQYh6PSK4b0BTKa4zNpvRg64PsCoGr87I
MHrfLDBLOIXoS83iKJxH85FOqO1UyMU/X2JOaUCMgLLhP4mU0dE+AoALxpkoaycacF+3JmOEAc+f
ArOq4XZro1ihpfh50Owwt5sBF5dnXGay424jfd4LOOYWmoKxVldVva6KnCLIretHcTB/Tu3sHXj3
0dZ86q9aPyW3roHHM9n3Jybh4aD6PqF4G96U8sqvjIT8rzmq1JSpcCSRWuoT2Yl/ZmyaEszTnbBx
imi2NgskILBA4RiGpYFW0edJjEfb2AFFzAfpBFhPSRtdTmKcPnprwgUzlTh+o4M0CCcwFnL9R+ky
biOnTz7+wq5GhWrQZ5yhGPTk6eySNES355pnDD+zzQDGCNIX0dd181WqGZkN+Dp0oLgeXX4L/Lf4
1ysAAhexYP2Nv5J+edgZwWmCbe51Q2qzN+AhQwkTFdoyrCi4E7GEs5fOBa0g1XPxR938UP81GP/X
VB7fvrGsqlqKUqvMwyEgXLgXIAHBE9ImgvXrfRjzE8Hpt4PNfHvNcMKTQuiXrKHqTnQlJUfcUOyB
mTeLoxKRXKH5KzA6UBnP9Z45vYk6cpfIGzLbtDnEKMcNM/flM4bKyyGcRheDmu04sysb5thzaKe/
jdqzMbOtzrwV0bDC/x7ezm7CZkI44WF400QMxw9KHzVRUamAx0VsRNtvfcOiKEwqiFd7hfmNLvBl
3OVSA8N2zP0MEy8I5S6Bn55bV9LQ20KmHausiDFn0KTUWS8rqhJSr1kn6Zkw+UTS3z5oTEzAanRs
rmVXmHLMR5ydxn4kBy0+DITtni0Arr+0GE25rJCGrowy3Xgngc7Wt4qVWtSEBL+M8aQkGIetqR1c
rPESAajCxiX81OV6xq4VRIjjAlmZ1uLFQW2jqQdboacegqd9h34b28zYzVYiA4YoEO31OXA4I5/C
uizjf2zOE5q228vloF811nBVGskzOQcN+qXTgtcaQ+EFj3XkMuDzVNCOJbnHQolFPzz53HURg93U
YTPeng0nGWHAtjXwFn4QQ8VeNzcQrgo55Q8H/RKn1sPzDzZOvcIsnS4xDugLqGDweyrb0HTyvgbc
65AD6vJz2kqBy4Tvd5/fks8iCmKtbhwT51jnB3jnYakFDRXvyTUTAf+GTqekrCdQIbdp5GvLGRv7
3wCa84MUDReq7piAoDGyCcfU8iBn6DWSzi5u94jkfnaZOFpPXCAovm9MOR2F9+6w4jYaH3FE5PKx
JjdzYCmdTgFRqTj0k6xcEAChlffiE6b0BwXD1LU/nPAVY1SdDYNgEyK/OJO7xUKICUF60MkAZaXy
ttrIJpTYChWeiM6nPV+1xPLxvnAPtv4+52FAwvV6q9X5EnE+CzLZX8F4gC6pEuwUg/k2RdS6DU7h
zRDOFMGZMz0dRgM4N8t+iye5VXfv4vAC8a/q5lvQHKImPjPAyscjKlUjnJjM3tZ20AJJhHPfzdC5
/z1Ywc+Vudx+gHC0JHYsMPq92tgTf71OZSkl6Avs9iXeULf2kjuWRwSnkpo2OAJdYIjYdd/GiDcy
NA/2L+AED+Q4c8U4tNQ4qTKGXGn8IFyAwA7InqazbyiBedOOuozYdSHpe/6kdFcCpsMQ85q7mIes
v/FBtUQYMWmZVqgJxI+tnpDKCDVm6T+wkHHandDHsBNrhlhRR5Q1cHMoaXuOgnNOc4bcYuMlELVd
IB/A7DZ72tsoUrENEw5Qm8mcFhKAPkPIFe/oCT+v/TAz0WV7/msmw9OuYAvSmmLIGP/ZSt7OMBDu
4PibL0uXXemQE1K6W4pxHivXQoaEErDqN+vURl411/c/F8VQlGTXRKx1oAJ/MEQEL0jcJI40O+Hl
8ElPrGtrZJz534IuYorcWZS8rNAZoE279ieyoYVf4nyhSmQgbhB9+HZPDVbN/DReR6z357gSJmhc
K6otWeUejENKDtC3T8ltCmEY2/mHTFJ08qtlVYYXyX7K1IXoJBvJtOE6ZHP2joN0oFTMRGWqmkWq
+x8eChyRoNC7NBxhf4pmGsiLlnr2F07fjyPbYdO+EmnkJgZImtxQUbZcM3redjmIxEjHzVY5uZ+q
v5QyFLSx/KOsgSv9IAzZTUo0wfAnRpJVr2dwyLDRxwABnypMALDC76zGAuPCzCCTiHtxbWMoQCPQ
jTFN+mwTLDLXsnXPVBc44Y+TvHm8pqECcNssZffaqZx9d7fXbjIL83UFImrPRQHfXQbDYe1L4eeo
X+ZNQtpdXcYUWGk+/wh7R70JkIRIZX5qBFgu5I9d9oyhkGFKATwz4swva928KwI/eIv0E5A8WZ7d
w+mQtSD7g+PSrxsDiK6lzrVhGxqbhFTbH4eqyG7AhTpxdCsIqY/JxWTGbtibFpusQZcCjOcN8stq
bmFL+FwMIbXWosWhe5DsGBP/6VR6jqJAlUraWBD4NCj6XgQJt29fNQhPrQgvUKITuLquJGnJ2cjl
e8HMhT0Gdj0VJJSUZjBx9C53yIwFybXl/KcI8l8BiLWYySXRZcBmv6D3Nlg1C8YNtf56iwyLDHJE
bwDOGsgmfVI4LGNEBGCm3n7COB6eJ/Be3WjgOFB7aCb/uA4aV9WNCf15iMdOqa0LA4vC+wCR28rT
Eg+SNGTJQJ7weedx/GiBTVWJ8352vcjhXJO9T5z7EctYQ7u8g/m+LdUnddqLifyOyMcIo17XUPVN
0t5dyXkhGcXq3sXJjYquuDI7ugn9URP4lpixLoF4/Dx0N3KHoQMLseNdtIND42C2+eZrDiUSihJB
1sNrFyUBZfMAX+SJW3RF+TAW/Tjdpp2gorZ2q2NpUAHbCSEhAJE54U90rPQA0aLnZfjSQQvlkQav
S/c2zWPAAF2Ngwe2stjLNrRpDOTW47mC8U3ao+1ndeZ55G+AXRfb76W2kgdUIsaFf3bKESXWvqko
kqQl1fmx3bwGuzNjCMO1s1I7JQKxKWcTRJwSn3Amc2sOokTI9Y7XP/mWygpxoEyEJdN+Udlh/Xg/
bg0CDuzv1JcuRiw9F3grBW8PU1fZ0KOLoRdgsxwH2EZg14zxCaJD086TCMlD3NaTDnhbE82eNya2
8JBDbnQohVacsScOtS3Nj0fd6UBoTlDGYikn+NkbdTg3p0py2AZ7YZegBads3hqjHaB44TamN5sd
CL2UIarhHpk1OYPfPxTPeeLjw/EmnnxzWhTyZ1728ABrDMQ08NvyGnCAT5JrJegizKbWM4tvbsGh
XNzqqUmddfvyiSJ56Xd2/tM2GVBq9gbp71MzBX09QRDzoSSxGVta/KZqiKxf90G3xaAsLoIrejcU
rIwlNVvXmIldwszYP2e1aR81pjN84blIi7vfiAu5A7TUqGcpJsnrgZJvs9rn6zCSSPMF/8SWGite
f5nvhoHZP2+G5fAX5kCtBAnE/rM7Rk6mNOHwtI1lkTTaRM5DESA6QvHOA94EFPHpS6GXiFqxhS97
Ye6dY8FZ+VoUUi0ekpxRPvecUqh2qdV/lYybgQ1rNq+ygbdg1ATTM+kaDOH9c1faYMoAw5n0gkUY
WKwH6/sSgmfWyw58Huuoxe7zTXBzsd7bsIj7LizemnW75dllDXcUA0MiT20dWg9LHXs+979efOA8
N3Ae74wlu+xd7szY4MXWakxwCVjQpnu5pBCjnuOl0+/PoOZKnc5QJgTv8DCGaymeAcpNAK1PJmKG
s6nHrmn7do7K0mgAezMn1sa/Yor0sHe/qd6tI4VvATLjyYzXeq5/vIVA9n6v1oooiIeFKJDxf5A9
b84f6x2n66WUcpFroFBiS0ZfZjDEwDw93rGe3hryAocntW7USnqxjsx469cTfXuuSd+86ebZtWbS
wXi7UKRG+VDy16zevfT3N2Y5OSI2jSO3/wmleuWNjMkn5rdrOf76LpI4V2Fcb9brY6eV/VXGHWhl
4HZH9dGkA7os+2euvT+Z3BTMUfK1rFuk2DOmf/lc9FV/IswdUCciKy8g2UxwXW9+8Rp5LCH4xNAd
9g1dkdQx06jj1Pb+GL1uvdguY+fPzAGrA2QRtmcO9qkXHM39tvERi2C5Sxa3sFHuW6qmZAH02sds
WQthbyKJCAhzx7YbUFLgomPRUPEKS51ugt/P625t3wMBmrrQQIHsZ+wCGmGhop3QowmAZZfZlAis
+RMFMVq8bgOqFWZhKCs+sW57k+AzOKVzXBmhCmvyQl6lPlqblWD1pwP2BWrL1dpTpXUvnPv79Q5t
aYYWHuHfsd2nokkPthhIqc8G9cw8tTMIOxh5VxsT1CbVfl/FJb37ovS4O99am0sBTvcKM/EhNmvk
XjcGlqr8WSCcHtuiMilFZSwrspIUt5Md5lHKgZxt1IeGNU3WVHZTNOO10jYvr6IpHZJYHpnmyALz
BULhimQxEYHb77xUCMPEYucauDeAdCvmWnvfKF5GXEwe63dAN1iLvU4xW1ZEBJyOcHrC8KPFcRF+
PkKIlUVomIcINj7yvVhSNdNDDfzjvb4ESRV68/+WRxi9nVvKrvBqYXe8HvOrk81jyPke2wFCMdft
jmF+qeIZ5XQuruOW9DsO+MQ8+B0e/V9TWwmvlJMv29UgKryDuJ+SEMPzbJ3Csv5l7twfEbhh3a7S
Ty5llZkieCrgOYhHbhJzADjq9bH+2l5Kc1w6RrBKLXZMPWLXdyMY4XsFawxyzR1dR0GM/HY2F8lC
NhIqtI26p7P2mUtvKrOnqRxW5xJMtDf5KhzhHvObjIgJ83mgcOFSk3ncVmsCWcW1Mr64dBBMCzf5
Oi7BCxp4H+j1h1Du6DJCvsdECMQd90dE1gEFja7318rXeNO82xMXRQJbmZA+zx/Y4zaRiLWC7vW8
f3iZoBctatiOsOeZRBZUHbr16KEjquUBpzq05XtNiNGlD5+XJNVQ5mdtRBNXZ5fh/uPsX9dd5xAa
AaAEa0iCM7V3Qo5ogzJyrVI0W4+rA4Drz5kRaX69ZyMC2OHJmebxyyV2KAUoJVjjRSfFXzQp1VRO
fBEgK4dom2RhOAT0Gx6a3jXpNX1lBlkqFQl8+nDS9EjLv5IgpeWwnyl2sKdxqPABwhhQxGUyNAZZ
KYiZ5DFogwULMI3C5sfxCYFOiQbGKCBN1T2t/WI4odQy0mre+3ABgqPUac9yqoU97BvSOEeP7niy
4bqYM4JeXXZW74VKjiSSd439vAHyMmuLKzj1LKNB7QfQasEZxac3VfzYBN1e5Kc7hY6Idyj4x1M8
aOO9Zf1uYwmG/X4lQlf2XqfuXQGJ75Z3n+zdMlaeWNwvAvkuiU1KHb7ZY21KQ1Gai2xSpzgCmYXZ
XuqeD4v14e1zH0ib0kGrofwm1TXLl7ZWsBWjRsHO8sKfbA3femq57UCgZUKlLAADCjRgNabg02Tz
BjU4ghZg/O/Kjw/umyNRRQ84FkD59X/kRd0uoSlO3f4wE9UfBHrpEq6pNq/ED3tMNpk5X+MvvYBx
CUwdPodfTR5HfIFPuCzfXS7B9QSmVuf9dxm//M1RnJM2/y9ieF2/BTrVLbCb/BEiAmxHvuNQgGU4
c2XtqH18J1H/o0kJRF/o+4VecdEL6KKI5XZNtcZ2WWf4sDygCmYOv2wgtJNv0WuPLF6grRwul9OT
PGi9Gm3GS3KxA67yd5nGTgDPdXXLd1tNFnU/A3noK860sWYSyf667yUVhlP9ojxsBnr1Qmmqca8u
hy85d8LShOw8gQhi8EQ8tyCyuAxpywMV3dr/ZclTIGc2hKyAnqSdXzv4XF6pUrr+MLndkFUFHbO+
Dba0efshWnH1XavlwzjqkbbJoWjw38eknHcmDxX9wY5xBSRuCfMhzyCruAdQZqu8v1EuyCJaTBTO
rIj3KJDk6Fsb/Y+IYXt4sPxqyAH3zCnghlE5ML5SH70HZtooqGUUhEu6EKZObuvQQvrrfjumGC77
klGdxxLz+uOVF09JkqDscwTDqI4wKQICs/wc4E+m3raXuTlMPQN48iuB0gGX6WAX5iyPfK27Sia1
+Avale8kHgkNj4DUjq7ttdqNTojEmo+6kURqiSj3e3joaWLs1nnn3iVOZoFy0PccmdPZ9xmbgStG
NuXF16mpcG7oG/0nu1UAMVz+A8b7S0vUqkCiyg/sqadZEhJxGa5nBj+z1co3XMips5awfk8COD5J
1Ynw6lVZlKOsgPTHuDxmv3pqU4ejOK3HmUgaGoMQbCU9BH4tE6eE2mmsXGEgP0GhQ83jHf5t7OpM
Kw3rEsIZOR/p/90ctodjWK1ooiRGJCWYvNkOXLW0xr8H1tY1NgHjPB2fLpCiFuLIyYEaHMp2jo9n
xhsUfaz27eWYcEkMAYPqYRiivHUAlHqwBq7mFOy4sNhpl8tGOlO5A2nEREgZLBOMN/5dKZ3/0Ew5
ky1XsQ2gMg0FmUMsEmWbHC7zicfgO0JHcxLGRSUFeWCGCDefz24MYEmHWCktDjvS6BzGroRmmBPS
rvAYw5Woeu0w+STQivjW7uqaymlM8jqTO3APfYigUOYunsiHbPGeJE9iW3Ggq2wytCTXNNr1E1Ou
4YjPF3v7FcE9dGYbRMy4+IrHBnkTdDm8iipOMCTOYsRk40cVly50GqpkrHHZF5W0m4GBoe0+vlOr
etb6uyFhuWNQaXTZ/WcW0GHEfKGGnRMygls9ZbicggzCaWOy8u4iriyrzZqM8W0qeT+hdr/Pi/KA
pku+XaGs4jT6i0karCXtewZcvEUSWYq9ZfMS+t+/dDIPvOa8SNnE62l/h4DBJId/7dOgNAihqAeo
SfY8j/8y/ipK1fUvfQ990ST6xrY6vWPEUA1jnML3MpDV5kUFjcXPWkprMWIDwZXMVgUT/yBncJnL
sTdHZOlqjeRk4Jlr2hLekGR3I5I/cTScUNrywHWQOKP9JgpI9CLoYYQXk7VcX4EdfwmpA+wgA2yb
pQYeflpkixBG8xQJtHbs6D+oRgeameQYPg9nUzpAvG0NYGHytjVfdJ1aec8pd95utYo3Jz4o7Xmx
DiHcb+8GbW4SIc8UwHL5T63PUnkAkqKf2EzgADHfG7ESSJ8MzsiQOQnaEsOJsT267t6Kh/DzbHzH
X5IAyTZveYWpI+QghCDUrldglOjJ2dCQymwpYI7cYe+I2oEyhdNM5C3koOWcDdHfalyvwOy6HYEM
96XuvjA2ce5+hVlxBq/LoSvCTlx8Ok5u40LZdjBjZLOmZgyoz2ANnalDaZCjfqzY8TY5RFMKDXu7
QZorw8SnMNo5ePeTqBWOqiiaMnf5ucFRrdIp40NPEJboWk2gT3T93gNTAcsTz56HO7U3F3U6Xeu6
UB74d3Gydjn9clVXtrT1mvyxkNhv0FJaVzpHrsf0oUhBROvfHm6LbRPjU9/oNpI+JyKHsZf60CVX
x25LTJ0cyFIA4WPt30Pq28+cY+xAEjt3OQVzeUTFtmcMEI1pTGk9SyrKWBgHcVGQnG9xYYM9xj/A
njZJpgvmbZtyxLHmwV7r/XJNbgioLVHIvapyKa2MmDgk14uYwe1HUXfDBNE3zbwbgCNBcFqAGrkJ
eZUEdXRp7LX/zDcPf7HeNB/g+hWup+yoy5lGh4icV8a7vplO+E2IkLPFzvYl4uJkNrkJsvY2DV8f
XTqYVkHpZBQrk5OxOaYskJ0K2PlSGaESYXY8m6z+pQmS8/6OvVTbnT24UmIczhGnCs+efiWjr8fM
FJXdd0A3duuarc0T7NpxHQh5No1CJW4/EDqRYe1WgFwLqX6hd6GA9UnU6DHu6AtX8wVAB2ieUBjI
yY1SLPL6/4iffM7IukfTQYIajPyN9p16CLHHERdNm30k2BVMm+ZyK6NFBxs/6JimeBna/GTk8EDX
oKnDanEQ4nF+TBgltzI+50sStSHo6wH3DDpPQt7TEsqsrNSw+4SIeEsV6H92g8YfO2kl6SmRNgD5
fSdtWxzqy7NIAAlr/bxmEFrjGKqg3BF/Py3GvN7QzSKEuDFXUvL1MuL7uBJHkBLUAY3l07aVjji6
XMDhWk9e+qInXFa4pvkDlhxtsGT9JtNhKigD9GRcA8kCH9ZrXzMaPN+++SWkWCTySkRbSQqmRctF
6mOmfUzLSKkUyfeBu6nGEo+RaFyoitotOg4MV8TK6e/4pMP5VtGkaOSwYDthxL/o6pU2d7txBeYb
QhMPjIpesZyV5i9HO/wlI9TvyQPcdJ+vbtb5N/+0cAm6aw8RJ+CF6l4eFVb42DHvyhxzyiaD2cjV
8K9nTXlS2o9rY1SCJI6jKqOtWUa4tnfa3iu50Z4l8lk1TEydRj2LCeFwlXxuoF+gLvqK560QNLzd
O4b1LfjS+MvuFpFP3lLsZN5DwKzUGJPcW/IvYIJaxj9ELihFGl1YigXJ5F43E8zZ5GXhqYrRnX88
nh2U3GJfQq/urq2pwO7NttN1chzmsw2P4qHeTt3P0wG1zqcxATU27CJGHGsfQdqRQDCUTTXk1+PE
gkHfVe8rUWUoy6o0MHRaZseSJqT+WVo8EYkUgk7/K6lpr48hc5jCtkilG1j7LE6IYzmDHlVu0kSp
CVTMwrfbU5n4zS5YuJB9rtc+t0xG1k/ljsJPsFuINtsLz4B+NOtLxvuYgS5pORHIH7P6pgJzXr+2
JgHGCPxIEWaOB987qRNYiZxvWx87DwhGVh6M8s1+7/GkC+Bdc/MeNXrJUUzEdOz7rtRYjCc7i8J8
kMLwMWOTEv12QolN5yDiwxSS7HaL27a3lCLTMUMJQNhkXq17z2bQc0p5PyLbuC0a072avfYB/dnC
VHGrtjCGh+jB4WjIJcn1NITOKSJbloGcmFR5k7vYx0ELQoSjZKPa30IN93u0f0RVMWqbeBX6Mipi
A1OYBqGYCOuGXZh8/QuuoTx/ENtdMtiZM1qaUQu6YtxhAW/gEUS7Yfco36hedjyYc5x9J8nzEMjJ
/yUpS28OHFpsuExrUUfMnYVjdyrZNngZ+mMDgk6pvmPr8P/9Ie1q+49MqCUyOI8P4xR1PKUH+BMI
6o9PQCJlwvhtHkheI21I1+YvaPV0RsT6pFOEdDTVEVGZRaXnZV9tY9p1fb2GAP8UrYbcnCd4Gqft
pfPDYt0BjL950cCo2aeo1L1yeK/jsDS7mSrLfWLxRenqreAoxHjji3jwSkicz8cCMhw/ukS5wCYP
ZdrCC5WBjp5eEBE0dvJ82VVeYDG9hJ3Lz7WcktWfywsiDToRIXwgfxXEV6O5CTUrMd4Qmg5uI9w/
yoPOol3yZJJrbex/ppLwR8ukQ1avo5iydIxgqhj+HosJPOEGaW6ua+95t0jzBr4WyDz/qhNEOUED
gvtbEL7B8DwljJ9N4E+bHSrf3TYFyXSaYWSZLMLjMsRWx28wu1i2oSP6JcxS/J5zjLPYv6zJfIOg
z34JRyxDc6FQbbxfooC69V4gp9kN0nmqzOp9lQMetQLZM850metj7RCciTbIRoJuWwlBiWwHdfSu
+8q0XEF6Ipr3VUkml0mvmHjG7iqPUK8rh1pam4j/B4qiNaIZhE7gHgRzPfFWKWfukImXunAzIOW4
VdWcU6DBBfr4oOcLYMSg+X8G28xZEFa1MqV9T4yhuWXEm1zPC+XgE+Wc04wz7tFZ+lb3Z6xKRmGm
vgqEVEhZU9iWAqqMpWA8BWjzC8d+unJ5ZOQulxS1vVk/XEO/lsGzbolTnck8ay/GtKe4gnnmIuyA
CHm4eo/CchtVJge++P0PDnI4bJqcrHAcEz35IDDNPou7Id2+WEj+M4f1Xr+btANgVVjSpDVuMumT
ALSoAinzICCWMxbNdY1I6SIi+hRryHpNYBIbQ+nvOidLFZ5Q85KFCEWDrUMnCOnKcFmBBdSwa5yl
+gvgGuiu6AIpauSxCnd0NEH7vEyPe47fSJMkATD8jOANgk+hdyXz0XFJ/Zzjx/mgi+twB6M7XntK
++Lje7QSr8Oyi4H9/3IM0VvPF33bMRQAO7IE8DJBVBuSISgg41hUJVFgUSjXiifhl/fQ1rNZHbI1
DWPTxn9wHj/S8+bFRS1ZySZfJurPYi4uNLWi79/dMzTVhSJSZp3/s2OgDhctnq/e3uEOwR2D4rRX
fiMt5BF+MnW9Nn45jA6n3QE2xDKo61CUyhl+1frbVKCcnypjw8wdnirmwrAq/YjYGXBefeDsO5vf
Xxs3hW3QaKsJmui8Hs18+e6avnU84Zzr1qqJhoEozk+oheYsDBinoapIM94qWQoAc6LeSsMkrXS0
mKY+VuSYj5/J18aeAVEqRMYm+ieonzJvDr6noFg6RBnTELNFblUahttEWi4PWjzYDfLnyrREXFrr
ll3g208JULVfiPu2qauC1BcSbJOK45R3vcFxH79lANokD8QsdsYVDjQ8B0Qw4t+RUmjBZjxJRgu8
noitHL3n/yzIAisgbnDOB1IdxyWtC8NxEpj4YNE49jskNFwHMXAOGLWBUXoXb9zy1jQurdDgo1S+
p6HV11t76UamxhmPTKsMjgoLUCwS4A16BOZLlApbjzizxTsP9oi9E2rp/1vC2gJIarQGfduwN/dp
k+oKTeeYniiv7Re9V1nG3j3wrXmzlDrYDgFHXE7ZlbhIHFutfNorMKFuDWj7gCfQYEp6OCUMq/6g
iOxucft4fmGSZPX+DdtiMj719LdTRGqn9qK4ajFwj0vU5etkvCJlEa0fwwsmrrKu/U04+HnW5Qhb
SZXdl3qnx+MQb6hKolPtcH9RiHs8piNPQa8eCQMfw3quKLfN269BkfTc2NAXzFualW+FvQJroaOs
9z7bOoR6/poxUf3qmAqvbrqIfa/S8WjS79TLYyzXBkQmlsJOvmOR9qHUv5birt49CiJWJUMw+Num
wXvuP56FrFz6zdNLiMaqe0WdS67+1zH4JWkfPczf6UF12g85x/Kxb7DyOwHpl3fHJSgO52m7soua
DOMehyvAb9UgZOCGMgLyFnqhkWGhBXoIP4EcvmflIio4j4jN+XObNOkviTPSZ3SwxVZd7KM1LEog
fwdx5/Z3ykuAhTGirbX06h5mp0oPTKn6SampX+xPlHUYnTPOOsrp7umoaqz0oA9jfSH9WqVX+BR1
eGZzi/AFG5oVUqPaSKD/Am1b7Ew5TCarvCh4S6FelTmca/xv1vU5aYs9vp1S4gIolIEkKOSzv+nu
romsdmbFhptfsWs57chvnN4nViaPmx7F8VoJT2lYTT60pXgl6tvrRdCYcHb6tJoSdDn5kcM1pCkb
5rrETZUUKial3DUsfGq2Pcd0MlmNmFYe9KxczzwxgnU8EKVipABiwvAarWb/XSrBmOxP/ZfY++qG
hpsq3/eWjuV7xQkXCtsGV2g8LcR93nAdMvpdCSL5BdEA67Qg+7HI4TpY5D+ih83ShxAUmJ4Ap06b
HQ8hLOEyYiFPBwUcQqLUxH5gfM2fcX6TChdwPXnKv4d01BnGJxKEwz2mdcsiAqaPbcI/BZvXTZtf
EZda/lsQa10oxD3SCj5oYmOqA+vIZW9YwcbcDU4kW/18tEH8o6epSYZljkpjhdjVGtklGQTfK0FO
3qTb4BSUoqe3dTR9vgDXrO+ZJ33ML0/294yboCmkdlF61ZhN/fvdDeMbeoOoArkhWsMzPbFmYUFN
xbMw37EnsjUzAs3TqZygdBX40Rfvzx/z1yJFvH0BaM7ERNJPTalIjIvxQZwh4OyRTKhRX+fGqe6L
EStKK5+U+BJ1jr/UiJD4n7sdMFaEsxV5sAXarD5Ym2tsHtfRamW2Wz8qgH+NwOZaLQFdQtf4G7eJ
vqeBskQktrawCAWaj05w3yxAZhcTVSK6JlOcX61yb/FGLSUO3dnhPGVD09CX5uyk1w70hMdSEpPM
lAyFkBZHqM1DBUeOm1ftC+f9jkjPc6n1OOyhtHoRZzVMenq3fpevralPbJ3A30q2t9GECqHfM7SM
x00hcODJCtA/C10qdHpzlCBAu2/sXE1rd07c0yrLRQFQqaob2DVbCxd7ZVotGPe9bIb1BKO8raZr
c9Ag0LggzfpVJdHF9GNVG2XIZDfOQycMmEiy6DkWlrlkpEU1WAOLkfxfi/PDMNztzJdMHNj1SXuB
35GXIt/dG0uDeOAgu7ca/N+IQKUqQnWQi2LCWD2l3xqJ/BITrCV/oKFifrFfuAPsR5g+5aruIVdJ
JqYW/3v+KVmpjifvHC4Yv6DepS93i97Yq6VV+9vlKFQ3Hw7qFypEGagnYzBcjfzKlJYgqOM4vH7B
G+e6k3jOHBAofY1CsoVH3c8J/zXzGopdKV/GngDM/60np59BTGUptaqrxGmLs29eo2olttJgAJkN
qwShaGZgzfxyqW8cIqq/vJOcJsuP0ui6xSjtQgNqAfwlkv53ficzUAP9LmpkMcqWQ+ubxlzuOfvl
f4De9vLbKgBPN7dndGr8ZqMoixl7npWGg/HayxGz+NTHWEwEHCjvoEwln4YIG81HTmpi/VajNK0L
ZmQ12LyL6iQ7iDa2msaoxUf4gX4Vhv8oJJzVaEBLLXJMRq/crlNwlf9BolvjIj+IxkNVdrfKQOmF
J78HkzY3CUv/CDuw9DS1zLjYpZ+7ck8CRQagANKcWPVVL6QkfnoW7M1zr9B6QuTcylpX9dhzn976
m7b0j0h3zki99Psw7YYSEA8TnN+l5jJ/foobuL8BpkVDQK33N+F6S59dHFXm+kxtpTF14e5FMQRq
Vvap+IogrnkLCnmuzOUsf7hYevQofm+dULf0lrNpTqUwjh328RQnnTJegyD886j50b/pIDiw+kpZ
AIIzP/6YVJA9R8kPzUScAkhTnyYToiSK2vgnTPR4xuC0IRtoG9gghcC+FzTYZ5wSS85HK1JfVIG8
n7js1WfI0oHWhhoudcaestesxx93y0tYuO80weAcuL7zNQUNM0wkRLPV8NdC2AIyu3jLWOr2mBnf
ws6TzBv49n7IG3cU6y2+b0ygFpdPava2ZyKIwoaCqhpfW/E1Tr45u4wPm+dNKEzZe1KJrfPzjn9V
WcW2QOM/cX6VrHknmPAaJ2qsakfF6zJaGVoWlM9nvZ7FfeQ4JMW/unwtdK6bMJ3O6X0QniPlkj7d
xtb0s7ZKH8KpuPwdZoLaejI4rhOt9c54gqS6sIjcFka0Y/Bc8fbbpOvzc2nTqhSL2lhno3lWkJlE
9HteuZzeA50R2TF5c3T7m+Gxn3A/Tq9T1ieltVddtRGht8ADkoMGbr9VmOX9wgZO66BZYKbQidfz
cottknnKswO9fTm6QJkTO/leh9R9HlgipuBBQqzJSZd6W3crcasw4WWGAGo5Ytjkonknl1kNPzO7
WMmpmEB4klIs/h6nxAbLHqB4R/xD3iH1cK5snFMp2RWeORp0t82Srg4duELXbc61Gr2Rcd5yW2+/
oDTDKJYkeIwfo1EVQ6xLc83RO7/fnb9maIP6KoODB+3TL9Xpnbi6KrxMIJ0eTwSK34BSqfC6pZkX
GMzP6H9wJOTIZJXtCOLMjZocwEte5IwEtGG2JvvfPehh7AuWLBu9L6d0co2fH/sf0G42/2r1RAEc
zlzj9A7hFNJ8yGeCksTYQTeyKmgklLvP9tCjpE/iaEk/ZIPnV4/KZBQglByw0v8rwSK7FfOmWwgF
QIngZg936m2uUACkVTZGYzUrNzrkamaOSXVo2fXAxvTfCnCwpgcunOyq9HGf3ZPneldS69k7FV45
6peEu+7DJiAo63vI4iE+sMn1LaWyEq7Q8mwmxgG+haGzXD0hoUVreAdyD12iX0LrFhtsE1rum3rk
CsYdCRepUNLo+54ywNTnW0Q8TFEaMVVai6jUjrpKDrvXhOTL92i3gLquhCVuKMeraaRq04ZiNNY0
8AFKnCzoXN8el+QfvtbuDhe2X3mI3B/Ct6KnogV8B4Bs4R/R3DZHelHGf0v2NzO+Zp/p+7SELJ0o
ea0TowwzV9HeIFwcGFf8Pq1t+jJHsP+WijMUchGhGmz2A705nmJWF8ockwNd7jQvJV/4+/U9d9SM
SS3Pq3UawGcJ57lAk3uOLFFNCUO90OlI3h+dilAs4QkYeSjLn7yxjXTIkVoe1lTu/O1n6/KaDDAW
XwQnCcPPbtpvSF4baWnFMm1DzveYKgjs8O2IX1s8KCthBOrMxiamNgqAeDlQgmSiZ1H8NVn0RIBV
Fp+Qd+Wh5vFTqWrdcYeY6cBHwgMb+WKf/+i2CxSzEGXFp/zfHHwAzA9uwScZzndK5Phb6/P2b3mI
8JvZm87frUiS+YkxrCu9CK3xrvv+85iGA5kgK+feH3CR+PYdIwB0WRyqvTCKhmAGuQEUEW6OMg+i
cZ5rV4qI2Htc2szRTq+56lVyP57liOlL4zwIj5ZitaKvtmzogpM345muYTVWbSdH6bwM+Ms48vPx
LPliNNmP4nET2y/vmXfmVHftZfgfKPM7ZQNG/kU9enKXpFAGwmVN9F6NlHpXFDKE9RN68w3/9y6X
VE4ldAsqx4/9DlsyYQHVBgeJxsKSPdaJQATtUdPAM4l2Z5xx1LQOuA85Y+nb3K90AVOqXX8PnONR
3ZxKfMrRqxs1nmtWIRU5fugtO+5vs4JzzWYbFuL3KamTBkNRez9DJo3Va68e1RWwWHf2NJWHVa01
WSvreujDyuByHqgapVdWPRienL2iyJVhRzYJSly41aHW2qKFrsEG+EM+R2K3z3Yqa+WOnJ+27Xmg
W7+Y/+HB5z9GOIeTqO3RTzRWtMkoH92Nox+nARGZCibuOxcICGi7fV3yhVRr0wWmZ4hd3s/jFHry
8u9R0QyAUFLuwrQDquiugujkIca0OyrLa65jiDOW6/1mHabjudcYGVau4t4aMXUI2baTtGMk/1du
NiJDPz3F/gpWBFDdRrF5xpl5OrwTzEprsH2dfrDejz2oAcTj4EUpPAiPs7yvyYCpTK3In/U6nfGL
KCwilCq/FwuifBSIrEQNjsTRC5PKTrpRxa2laEgw2aBkLJimh6Te51+atWz0457AeMYiSbRcjcjy
/bdNSyPI6s4CIWejhpYg8Rzi0owEBP678N05pFMiWVzqccEt39tzY0wSSKMIhvyg8Qze/blx2NfV
ylXAl7C+5XzKJL0pMc6fk0hEksmi/Q1pOMAw6B9RYUHAGg9seO4UClg0pmd9VPCIHrmcyd4Es6Nl
n3EsDW8Vh2Dt8Z3hQ/syh9EzZunPBfpXWUhbJ9W2VeTM/ZAbPQdFS+twaxJDxKXC07Rvbsv3CBTD
wPKAPPAIgLjAr9lX8EoInDyGE6qGV+Wclu9jiAP8KevZGwLml67NLdoVSSVNOVTbafS++ZEQ4X/6
wBePolpnug7nar+DdhYCQz13KVOjNa2BFEP/NBWgTescDxi8fEHVpfeVL4IS2jOw1Lg2Fv81679B
2lzVxtJlZBHrHQfa8rsLxsUc2hH2DKQ5qB/7dYdP6S7H1/JPAtzhUKdDLoH8vNRBskGD4pdmt61D
YAooFaazEXRMzk7t7bRMeM7Ojw7zstnOUPyGY0Df9EzBFdEDtnE40nEAjtSEMR4yxSKt7Bv/zqmg
7OC3Y1FcAagUVH8GGD2YUp4Yik7hh29P7JeJy+xSECzlOb1grmIrXlY4wMYY/7YGwqJrFuNfSI5u
ROFfTScI/VXZSpsEilvXGFz9ggFsw5afWS0AkP1L4BpRv1V5N0OgURPvmzvV+pSuEmRxHU4PS+Ol
9s6Wp8cKL0O3HkCJA33ok6EwLHNgHsYVEypSCJTu40cmOjW3c1+SVsrZydANZvIlxHoP1zIeYXLz
BW1W962rtyWSUPF8zvrOPLxy12iKK6xqhEet8oY0jTKJ/D+PmWooHyszqdMriEGBu2ZXoaAbOb/8
MrLlf+zUadSv2ayl625XnEBLSUicp+bv9oMJGO5K2qKu2XX6xW0OshqG13EovV7GHI25yUxg1oh7
Rbi9Uwoq84WLOANDtdFckkyYvS3XvIiF7e1p0Hetvj+SWRHoi6vtJvf3oQWJwUZE0kjb6Jba/QjG
KJ5uJ16+MjX2J5pkyJEBUs5D1Qm+8EptMG5m/9xZzA9OX8O+01ITve3pTtrjBWnEnjVDWgwjh/ra
n+dJDdgWRK6qeoXZZyiy/qtiRsmNNVX46g+vxH8ofNy/aEC+6+dPdxtJuswjvALs+XeSX3jQRK0U
c02F3cBGp/JgdVfrKAW5UwUyBkkeYpUMR/sozreAZEYaDsecIo1cZGgNRTze+yKklKVTw7BOnOyw
Q0ioBnwK9ghrqiL3MqSHjdWvbAIZ2FmF4r7bBUN7AD2mXYL9Yj+MJ/UNN77BGXFJ5Gy9WXUMSDHq
cWc0URjFygSISDuM35g6YEF3qXZyL6HHQ2EfGIma1xNJAilXGdJLNw4jyehWwYxs4NnmP1LTfZDo
zx6uzcZK6K9amK+vjBfYir9i3Z6EWHiCqBRl0L7TvdPAzmaJ8zxsQcHPuzJrMRrJpvQmGkDk/Axj
t2739iPphk1xOQqzjXzW+tWjLvoLPGPWfwu6iIjB/MFJiQg0Y9G8N/tI1Wkj9VFxK9iWQiHnh2dS
P87DjJMPFy66i3Y5MnGUaYZaSgC+wu5fqY9YwQuOrsoVo2lK3Ayekxp5il0YxF+nJNTF3vBzQlIW
qnbffXPAvY0lsY4mc19CJ49jdcanUYkmA6RWXW2vYYwYIegoOUJr9hElvWiKrHTLwV9qG5MQe8d+
mM4DDY/0dRjVMEf8MClr+LjGz9joRcEHAPWjK238PwzJYn0e0a5wOmaPaRsEQacsMtVpxWEEdpqR
bCEzY7Vy+dNIjxfJ7+mTiutxwTrRloUMQDFGJtf9Kz6XH4uawiCwrmaUR8Fw8I2TZg13sNum+PQs
o8xAQIIYS+5K/GmOoW2PJfh406jTDbmrQdXxf9ERMzxB9mTicreyHDUB2s6mp693SvdyjeR3KyIp
WrcjDRHMQ4CIF3rIaZ7yjaqjLqCsummYuCYx23Z+QKCTBnhSCdKbHiTlp/SnSKgt2jOVfaJEmv5v
roF6yMDJu7F5x4gSl0gKiqBfETSCCwv92r+KUwa1pOxRbGK9VTyXi5U563jLypro1zodc0DUo+EJ
J3dRbBDzPGvqPzqQkAxyrr6JyYutUWkLSAt9wIfToyTVCQP9+ppPo6GOu2UBK6YsqWq2xLFzd1UV
/zeYeHsYJ558Dbl/ue4ym7KUhXjy9XMinwqW0oAS5l57Ki4VJ4pntuqpo63A3CyEdNBCWS8m9bl6
Za+uJjzgjkZzx4JGd9j4BLzRQ0OctptaoZJJB1NArPQN9W0K2vUR06x5vqSomHerOWukFJhCABpM
hiP2ES0WneQVPqeK61fHUNKeei05ky0lH2LOptGdr6dp819JHtG17jN8XAyoPnA8jCSQJwySSGYj
wF/IpPFQrXtUjP7IyGUlBvXo7CsasWLadcnnAoaHETCqQo3ZWQumMMy0Zy6HzDdxi6JtXbWYw4S1
E6A22vNaR41beUXpCxtC2c8BuGCzvHUBmIBeRdqszYFEzcxxj/Yw7iWa7rTa0Cj0JtdW4+J5xKlw
gRvTs1bTTsZxZCtFmLa3SFkSRgF6XObEFM2CzaDv5EXf51NSkgzUrrqSPJbPhSKuxWgnOSdbhggo
wWftVZZd6hu/auTom1cskxVcQDkCFmL17dF8fvIUiwWdLj6/cNgzF4RQ8AtLBNqD6aefvl5uL4Kw
vejOlhyRPskzxosSMSGhbGa/rxFyTW0gS4d3SBRVunety2aPbF+FgOcSNtCpyPFqg5NL2rWfdGUK
aINmhoLcN7vG53XWZISHtzfQyflGUWyHxLTuCsCvFFgbfJzyTCE8NARSI+7qCAdlgN8tAkwJ36Mk
0MPDUxd40AvzjM2bf4ncV+4BVP/sC0nR+bxy/b0LCRD6QAL4PxdBUkWqE3yrsUHHNaT6jhlWHFpS
8QzNvXji1urX4CcynSe1gfVQCyUF/WEh0QRhbB8todNrckdWkbtM3QLDJ+46k0Kynu7Y19kPk0a2
RC6UzWrwbjo+a0ACGGGL/Nf9LKq7k/eBZIQQnKb6eXsdvjr+xZRY6KJa4ZL4Nzn2pshH8g2FleCj
46YwlWZ3qWZS+sTYuf+Le71I93BRqYdEw82aaF0uazzwJ3vINFlRqZXxVeD/PF9RShHhzXq1L+Rn
ceoSIpZdznjlwVzeLvVp8UW3JQMH0FBJWZ+wNcz+w/OTqAuzHlb3kO58p/PJoXhiLA6cU1J0v6I7
GhrMhG0CU9manGZKESLFUClu4ACOj5dvhOPXieNgKMkRcigtRkIw9bU3LIBK19ZxqX+buw46wC3G
QQdOcW388mjZd7Ttn893Yne4neCpmi74x/k6o26z/YxQw3Q5XteZKxdlBeFASevibv43vIxqD7Pi
BKyScsl6/b6IwcqLwjcQEdLg81wsQIJh8Guc5iG8GlcFQyzLW4D9cDYGOODLmGhJofxha6M0rncz
Kjcch2rKuyblgSjbOxT1UfsE8qwdaidqhR67e0UjFX8IPrUCzISdx8aoC+V09oDrz9YyUbxWyFxH
rS67t3j9qtkf7Lj6aoSt1GbvHVsBL72N3nAUcIf08Qa6ozf7aHwcpiN6FHQbh14MJVWwB0MgojkU
3udsXEG6JV9kg3rNQ8l2L49jjI5ERTJZRN8SVnmQgddV+F4yYRFtRKGPMDOOX7Q30IIIMcRuFvKo
jaCfbr3ZfneUZQkdUjxOl2HguC3GCL6PJAURy3aR+LJCYTdPeA3WJItVXAlYhCL0Nua752RK3zRo
R223raXa/pEe7kqZog9CmWdFX8iXaTPLk8kfESGqjGjqLd/oRw38E4uJfI9yIAmsXKeUHQXhWAia
GS2ZoiYwEGNCAQWkarXFnpU5d3POh2ArDZd8JEEP0+T9giFZdSVFGVLrHl7Z+4nDDlS2A6/kLzzN
qTz6cdE5epAKXTFVIOSGSoRJCIypJRYJzZHIkGCgTgLNN8Ee4HG06odYsu/zQF2rJu72lo6pjJAw
tKFfP1pIpfyZ/cAUOZVEXqaOxSjACHc8Qqgm8YMk6eXD4yUKy3+9u91qkW7PjwmbnnbJsKPpkzNr
DAv+rkXiKPEgV2oJatE92UFlGj7peIjiZL3+PvXBfKBtcB/wrsLl4EW/F5w6y8qd2wswXGElkkvN
KVtYIbWQXE9B7eGEoWYmXY5ICAfBmBkqMktUaGr53aecSDBppyqZu7PdHvUS5oLSOnPercy/IO4U
EZlVS7K/DEEtN8h0Ko8GzjXVGL+KzulFigxIdPtGKQgCU7Hg4qKyLRZOLkuCSJMNSq2m4q9DjDeN
pJRyKSKUG+QHG4BZx3TvvhhBW/DWwfPr++sbXryD2aiNzIpySFAbxga3IexYrXgrlfYAAbMUi8bD
C7+QBLtByydTPwmKGYfMofLI87Ne/R4clFcKc8L+xrBAUpz7fULx2MP6KeEOirSFz03LNgIcZn3e
Asp8ZxjF1epHbIybUYmxAesZu5H6MoqcdHiyfCTvgqM1+Vy9GQpZRLDFfy3WvHrs4nW0rzk3StxP
+gVoxGeLEOO93JyrhVIjZFI720qUUwMs0YN5XlLh4wRvTHWEXp0z6CfH4olo6ZMZoRh/OetLTX57
Td1cgE/Avp7SxjF9qrc3zbJ1uCgwn/zxqrTcqtnu+RULtoO8rubLuOn9xo3cgaTxd9bZ/8060ut4
0r1GYQnx93CxarKAf9Wwf4f/hTPMX113HsraNwcX31WMsH4lUVvCOmVmXQhCo4IHRzaNJT8CPmgb
BcLZxcssp9YZpBBJfC1SxrhQuTIDujt83W575mZ17bCDQ5DMzd/RErCIevo3hGxRMUUCvLbWU0FJ
jIeZ9JD5eTnudEu6I6W1lWCVGMCI0TO1JyGz9CiXKg40z41uzfEIAXbcrNU35uvZ8Aj9ye6Ao7zF
ahPf070FWMABimDav87djeAGiNGTeRpA0ilo2Ky9y3rM+pjR/PLbfF5Q2ZJ3UmYpJsi6MIZCDPXF
OAJBh5LS7jijxlJM+FsYYVJYfPGZNNiMIqOv7N3b4+tCVLO1Y82vqAn6W1ibgSVTW3qLoJsX1tz7
kxE12rzNrtWj+P23PtkrK/vlpkRpip8MY6XHo3jz564ZqkML33QYC4yWutV34sdTNDfskorn4Qd1
IwivB8VwIAUuawFYjqElluiihRuOFcSIruRwhp92cpPz/2UAuN9YeWHNv1EJP1/QRmrLgIZs2N44
hsuaEvOouOi0qqP6MUydTVmD6Ht41iq1wkQeWyjBnEbqLJroaQyh9Ed4jkzy5LpZKGSYQHcsLzxe
2P7w8q1wxf2YLLfdeFvRAaQ7kN7LzmOAGCFdEm5K2qFYdTsvfauXEFqiSpDu8nAH1Rq3XTrczdS+
nPRMZdGSnWh2X5DGu2imED6kxRC1kGg/vrvJUjEdJtOxaIFaPgPfrzr7cMEtgGiJthPjjzrdTq+f
CdJV9BzZLfdbn5eF72NDDrZKpqR2ahFQXNt7OUT+JZSXaV+JTN99IL/M6lsyJ5r8AcZ4N9D5r2rj
U7XTxdXfTpQYTz6yj0BzOUVaZYgIUmrln7073Md78l6dBNVZSyl8++MaHfLz2xQ7B8LCdCiv3MXK
q16n/gqGTJ7lBWY9+iuzwjKfH2IIw4wt2M19rB71orzxjax1+mbMxXofDreXP3uEcUBlngO0UvJw
shpaGQG7ngRXTDOxZmXsaRuGszt9W9HxN3egjOIsXNKt6KtZRh5IlUGZAcmCEAZSDUqETijLBscc
dtxF+9bjVcEWrPTWFD+VZFm0vuNr4EQgicppfT/D16zk9azvnCgC8nytg1Ey1H2uxWKJuk2D9/jB
Y8Gmn+hKTbLKPFLNcY53s26SlXaN+vI+I1IN0LR7SACSJBSXUj/KCZNB+RiiJucPSvuDs/bPmg18
Lbclw/kCL31JU2FM75U0eQkHw9jB9TTSmGuDnRR2oDcqj4IunAJgYpju/Q1di4/y+RPwvUZOFIKN
o3KnONaUWeOnUUb3Lt6M9xG7Wgyb2n6PPyeYMePzj3dHeg+iZJiWjR2uWAc0az9n+9P2KXbhrwZU
ho8TblRGtSZwuIRv+aLhWXGoZoaeJKGtvnGjoDINPLtPP6u9NKbRJwp+kz1+z8rXKYvLLYjKPmBd
UJYIVARo0gobhFJq1OuEgSQCnrRIwHFORNZzCfuqtLAh3+pL7CV6kStRBeBV637bN5pk0hjV89E2
/2gwdJcoR6MRR1KbqQyohG0ZGn2EXROH8qXjCq23HBipfW/DKntiWlRvgC5MHqQPe81HxcHEFSaI
yCekmEWpntGpXfqfWFujVOsiMoYNzDQ73ZpEWrRtT/UMidA1bsE54y7uekt+BjwtPkVNyDelxIYR
uOOsDVjrqPw8Pkm62kiWsofgYl3EoFFBF5dYt3jeIyvb4ykUUtUaysWmBeYDvJnIBLzn5N3tGufp
7K/ldZgTqxYRz8PqywmjN3FTTrKPQoXMjxdKcunpZfB5SS/OIv6VP/QBu5KbLty8Y3sX4MZKgxZD
H+Jh6JpcY12+nfFPUekvRk5XJmFJ3nxavAsaQWnoiy4PZ6riKOgMEahGjAXBW+MSF+AHWIYhEBEy
N2VWqn6WHHTNWAxvvwmhb+oOVO3WzPSEzMOTv426sWPAlGcgvLo8WRaRpvSfqhc9qHXKQGkBkCQL
/P7RwQwATEcRycTVOahS9AloaVi1x1YTX9gsYFVOois85CUJlTBI4+7Pex4AYpknuqOJ0rya5dQA
mlTgb89Syv1Uv2GVI553t7tFaRcwd9uqBb9B1K4CxMSNYUkM0piake8ybFKgzQkZ60JITs0YfYPJ
aENh6zwrR5wUlvL5DXPclhN4a33LsncOVoIfCfEyfiHKi5M8ItCz0VxFEB7fScFj92FjKeH3/g4X
/VrOUlCwe4ID6WrMdIfFUP61wGpR2VQ6OfjvT2jkr0zZh5EEjAAttGnorQWgpfHRLG3nTpMaV5PW
gzuEw6mPysZUMOgod559dwHFIubMVYvg0UdnFV7lEReEZy8cZX4L9+4epSQo8jym/S9y4gFrYbUX
fYIG7sZQXWNCz1KxAGzLafwS0DmhaGepJJrYlqgXMCKclftvRLPMw295lC8FXdioll0gezKTThez
SES98k/VHNWFDczAWlz1AzVpQsK3VvM3NUjnvpLSfvJF5Vtbd9TLv//np/5US/SOEkS1VmVW1v+H
QkFChPxLgsE/2hZkz7mOA4qs48tuog41PVPr7YYayDvduHICXpt7PL+WCmG6WRIyc3vD+s//71ql
mrPojk8sK2CQUmS+0UmNZ/bjWYCcfQRhY8RG/f8c6gsFRtdD9RDL5dXXP5C5ViWrqM2EM2o3N2Su
k/Hb8q372d6dIr1pb9VQy0CjLqBXNNJT4OTU8pExF4T2iOCHiI8jcGgTtaPRfRFWIWjD3Fh2v0k+
Sw2CLRTxU4Y38mNeUrkuwx83pmNsLIvlqt5rtCxv0flm4svzLR4iE4W5zZ75sCP5To8zpycqrFz5
xWvH+eaNOiCX8kScjZs+eKZYcn/e86Y89Sg1t3KMQIQFZRfdaL8/a8Jdx3uQF8/8lfKn2UvWO0Ox
UesedD6h249C9mP/Nfoa2fB/4hAx1MzEvHVRs0lmVxBZ7txP8l+g4xoxjas0jsDbu9YscFvuXhdX
yL9E51Y2IIpfDgAmlab2NDe1ooBeiL2q/FWektVc+5SHotEtk+IXDGvUS7Twd1hrA0Q3/KlZuAI6
yv4QbBiT8VO7oseaSKqWdF72ymlk7W9z7UvkTJYldB7Y3ZPIN56Bl5eXNbmxWziNh6+u8flAEHZt
pvYLLOZWdXPIvJhNbUCqfwPaXFelivGwoKIJvDjWkdCg0aucmBNhlJIgSlFSpYLQYS2YWxSBaFJ3
R20zDKlIjZRCrgBwu7yg5BINiLG00Ah7DPH1CG02glaCcoifHV3Ee1seUuN6+wBkshwO5UXLEqHq
NVa8iX/fkKkDJP4CRJcNpaJMwjm3WYspjBPnJ/GZR4QVL6+QOPQC2KHChUfYglu1NYxtvb0fWPtH
gDgH7AsMS0ee2WtdX+QbIiq4i5Jpy2DTBCZlo89/1X8bTG52rRa9vGvNV8mQ5vsL/h6bE/VrclUd
1P+eqp9cj949y0HtiiBsbpTF8svXd+AJz1eJFNPsBaNUlK38QMqwAkJvN1EGJuY9keqrMSAAU0mn
S8HRUGZ8RKgtmPTpCLdhWAEc/+foCMIcd4EZFFU6p5NGw44J+p9AhwySR7R2gy2LgUNVC4wCOlHB
dV7uyX5E0LtYGmEcwNg6lSVqkY9pdCD07yO+qoYcsyUBsx15kTD0k4/VlnsrkWQ6QzVJpoL3rOph
CZhg9aFU8upz8wnhXDf+uULMmePu7ZD7mXIffT2KWzfJFUh3FY8SoembDEhwhIgD0uF+pNp46uPK
bj0kLu2qlKK8suGq0JB1MeiJyKMU2qbu9FG2L8AXNGGBFRaxj2poFq12WvGda4hx/VGmUzxyC1+x
eKNMG7pBTb9a2d7KqVhzEuNNaa8U83NnAVOmBHWxOQLGUR0pzf8xwb5RROojN3rxG6L25STphx2f
N1AKr/Go4vSF8NXtm37bdF/dYg5weVFSC9v78Mwq4KKy9B8suCz/7yANlgNpSZ2m9eMjL77Sq7jW
mYtbUyG0fqU8Sz/sizn0mr1U1JUs0gqe2ETX3gU+ZvuryLM1heXIMqwlypKdatI11Zcqe6u0UTDx
P2jwC6CktUaAVGfBsEUYSceb9dQwioXkWTfB+nqP0f85IvBwTNJMlWfoqLH5a1+D80QJ7e2tQJ9J
uqC5IjOQpU9Gyt8/WHk9KeUKnarwZWLJ/SvHYD0pVnJCXbHVKKDkLWut/XPLv2GOfrI1AVzlujG4
W7Z142kd0wQVVwQKEzmYeav86dubCt0AZyWRin4xOjQdeItE3jIiXxxGCHKnavHXrGTmnbqbDiw3
G8EmKaiUiOIYyDgdxZbZs+2gyLyGvPQ1LRMlSTW+7fRRraHNSZRs1wtHXg54pt7+LJ5y9+O7Q1kG
2ePIhlbyIQnyFCYG+kwFVzE0i+XX4yKG5HAd9Vgh0fz6eHb4zydbmcHar4aMvAUSld+/opSxJQL3
M4k1PmxGAMSIhQevSvwWYcCJFQH/qpp4mAd8j6/TrxD31lrJl7WqmrY5MvPJ4mSSK8xTyuumdpLK
pPHvS5SjEAJFhZnx3bHsDX3oisAatJhJoqIdzHghL4FFn22XEP5NkxKJUFMaPtYOxdqpbd/GBvjf
Po1/nCufIrVQR5PPOi2aZk+9GuOBdPWKgk3fWZqzDB9h71+cpKaqA2nGvgm+QC0MErBmPNZK7JoW
4I4t72ok4Ba72/ziFf8sClUB4+vp6QDc7KGZxOjUOL8oj/77jvpycYZxItp9Dcc08tZnDzMl24do
6qq0wQGdVHIw+CMVs/Q0KGbhe9J3JCyaGO2hW088obLmfK3J/NiKpXX+vze0ZJ1XGDKGwSh30zk/
Ixo08de3kB0nefZ+d8vQ6rWZMlNQw4XtWx0brH9Ext1pUylgBqzP6zyWUXRAxp6faDFySZRkQAqW
+1mM+QgyUksX2qVDyuS5z1ix8xExVtAETDJBbyIa+VnA3BBCx/00nnxItOskwogjrtaQzeFrAB0L
a9b/eS4u9eNLNV0d6Q1/d1FmehZ+oq124CgiLpUubGeHylteUJgFatww3IhUkYq6kjdS7hQtpi6v
bCWAnQx6eJPfqCj97tExStznsOdqtvroEyRjsfvUTPjpdv0SLWk8RdwdP3dRjQnORFfciaIKIhJ/
6E3WUcun+Vovbxgrx9ORMN2YnWwn0VLTlYIazsoMLABhKTMuw58pALPkfGBWCOnf41aDy8ZlI4Sy
VyMoW1KRzE67pB3VFV9G1BEC79Y5z7OdHLGgyj2R9ExnKNmNiPT/kmSUF+N+T32FlwW6CmakogAs
dshvraGqruCBiXBg9n0eNDiQfXdcB1UpMnTEQEyUW+unUETPU91nyCPOPG/6JelfswWfqaRD958w
1zT8yOTQutRDDwdG5LN2CnktAghVhmTWZsv3LqfHGB4X/5J5gIdlfNm9w15Lkke5+UZVZO9eBRMr
JgyRZRU7QLx5XDF91kMH7mlMoE4TvoyjBaxHZlkS6+jApKSWgzDOwpjwwrXBqRYicqwsKhFi9eKl
sabqahTUTkJYwl09HQl/2YVAqdfKNg79xD84p0gYtOrUNxVeoN9T4Q1jLWAyfCeZYVewLKkOJx0C
OYTFR6npkj/nukE5WPKWR7MK7leDG1E3znx95SnlN/GBB+0kFlvY1OFUOckqMgYDt89e1K2ml5OM
yxsF+S68lMbwDs0u+VI3DsZZEtUb+m1Y6Rk+vUkarW1k8Gk4NVL/kq60z1xf0O/atd3JoOq3hs7w
SEJGWCJbXcIgEc6wkq/4ZJ+/pVBpppIDvQeDK3sYou+YH1JvHSjeChc3chCUBKWV1a98ZD5k1SX1
7ae33vmY8CgZwzU+Gz++jkF/fnwM6mWtEVY0cbO/MakqEjmn0749SkItlNaJHcjDN8O+GomtSqHq
ziakd/+xPzIvbdLSxZsoD05K26kqEGoqcDywn9vQiyHmzuEkNOpRUHPyMd4jHKiGVx7lUBxnClYO
GCRVVCOxy+tzGVN2MAoACjxx5Hrct6zkRp7Eu0cj7/cuVy32DnsOGgecJk9xCIgufnjsC1qJRwh2
eoSOckLA8tqiwprCnHsZZ/kJRkwgyQq15ktqvti11vXtUbhJr6nUJ/2Fe9BxAM1W55NMUuAzN7aF
EdO8J2T0xSr1EZzX0R3g5UEeqyBLukWxVmJ9twQ4oWRPL2iMU36M/AUF8WszeMr0/5ebdJEtZpyc
1ltowv5U+jmak6ya0uKF5BLoTbrCRcatpYq3eH6piERCkkcoUlhZ1OSvhKqeEP6ePsiFYSb1HYAZ
LEicrPTCaXsgPTdzp6yL07PAIZnryZ/Q7KWXy/7Hm0lVCD5+PabjElA46TRTNDLdFIeSFeEDEhgX
aOs3h8wjcWIGCDGf9Xx5ZyNJbrzP634ac2QdjSe2t3qf7kZ4DCyU0vDrhZdPypiGllfh8WPIQ238
0IbTlSfmiyc8/NXm2U487pkC4pDO3nTfjkTLQkNunY0WbCmJwZISw1UK3tck4k8qlBDsZZRGi6Us
50FTEmc7Vsz9qruuQQ0FybUCUYz4YYiNMcvY840s1KidBGTeazJ/WhlttHGoD2NNlJ5j+kTFNCz6
hagI2OXdGng5I2Tsd+uF5WNOsct83RHTrh6Jh4nJ3rSqIVHfMrqRsUthVeAR7PqbaV2Af4a9WDQj
FyJftXA0F/A1BME6xBkUhsEbKFis8vQ2a40w9KLM+4G/4BibHvtpb2pd0tylwY+J43XnAr9pnZyH
/N91HJMLFFlh3cklY8U/9dOwuVoKQJJIeY6/iwoWusEtoDzQ1GF25xbjoZvcL8tcu7QPmfey9QVp
xWgt8zwbZHm/DPdhg9LvdweD+fmnc1aJ5y5yI1tZrFF/tilXLdTFhYSL8nHQZwEHwReYaczrgqqO
BEt2OTegvYRztkh6CTNxRvs9k9BziavD85zybYBznw3yvJwTr3QJKtUmYXZkhp0R6KUtF2BVx49d
0dam9W8AYEJN/Na4+jK8jsxJgWRvnSJ0Poc/5ATnmldH3gNYstoBbNn6bSgPOXumNjcwyOHia0M9
48pbo6galkN5sNPlLBpdmO/Zmp6fNfJGO/0iJNHsysnjShqvaEOiewXGbNzd5ZbFHXI62rLSfXlI
Oz8evE+wXsFwRHDWFAyNDpBE5b78Tw1Mwro9PauQvNFrmIaeMfOmDcGdBTLGHs2J//L1IvX94J4h
VRnTveZl42NMtxiLBpS/MnQtOKwsPlfUzTF/Q7aF4v2wc8mr6iXdK4HHsZKwfjyUfe4yTuhwyrHC
GQlJfSB0anAzjqHzUJ19EGh+mB74s2AwXE+Wov1zotZpaUcXTwBAkXIG1nUWO21BJC2m5Rjfn3Ky
UHJCR1rJpYCxCj5/vo3TRnUUDf6RTsytfQWya7Sa0a2TCdqG9m4qERv8WnifSacOilfKVJMvZTxH
f+OdG8FAAa1Q532votgvAtFw8sFWC5RnKXlbqmUr689FGvWYkCbmKNndysVCefkWiGNqxqJUkXTV
fRq/Pdqye9q0pqCIXpwV/prdNCDZE6rPcCTmjI99xPxHoH0jFZ8fuaeFYl+Ml3NGetCkxl7fOEhq
qo9K8FeW75mF5Z8YdI1HbPJScdP9frBSZUt0Nqov/3mMDNC8x7A3ScRnG3he7GWKarB+av7ODvfi
t0XG1SFsL8HVjfs0SD7B9rjWKVmIEKON/1fyfoTVTYEGWMnctO2sB8LPgvgZNn9BcyVMjl2HplvX
Y873N4M9/74fBaMIpm6MIYfPysNs2OMdcwgjqwSXkoi1cRQMD7EPRYVXkQTzi84u04Y+fOgf1Uwk
yIAfbQF7obxluklshMN381S//++zHWa9kDeLK4Dtodwb9vALY0iM9AJV2uiZ/VEeeWrEw8N4Uaw1
rIRCukl++WqhmNa1g6NPNg7hIgVXVItraJP9pc2hA4xdTUOIGvWb2zbBkilHoQdWfRM8qnlCHSzG
6MSEorq3Mpr74XXOwc3KtM+eBZI5RW0UyU6kSg3ZZpe15i/yHas9NIg0PDySDp+I5s0qCjn7xjBR
etZtbBFtBSmUE1o9Hu3wobmISVH1pYM5BLQdcWkIYbRK0YBB2L3CZtQZ4goDrngQRXYeodJsK5qO
yhv7hhfuWxOqtbGwmlP+kRQ9r7eivJ96HYQF5/t0SVGOLYlc0jkessBJ7CAA2Jk5LHpeZIYc7Vsk
wl/3c50QyxvEZDRNc5OBDH0hK9xygh6r9TqjYRKnVrI1hwi59AyiYC60fAQ8o67mUl2VRRCoYeG/
PGI+VPy7siSGwFAB3vY6q0a76JyfitFOX2qDHQ8pwfjXKMULPQwbr1kS5JSagl7Yxt4dVl0bheTZ
3Bjai/vuCwg6Qry+jkGkiXAG940xHV5Y1Doh4WQAF/TF8069aaYqg5sc1C3XqU3VWG2oxEYh/Ihr
5I+8RkkMMQk4Z4p3gn/imWuvOLhEtGDIfZA4ovG7Ri+56E0OgAAN34g6aixXPtQPcWKtiMkwZHjB
SceoyrmczHrO+GuhReJfLj+9mYo7w8S6wX+GhbfoT3sqWCfqg2GBvbEoZk7e9ermLWviGbnsJd18
K+KfhVhmea+oLFJh4UU/6elJUnVEwrSuWQ64l8PVvY5w74L383Afl0IVzviQqhh8tV84O2cEMQZJ
8vhFzH5z5gd4dlJWfXfNvpxFAh8ajHwx084EXj9NvF/9P/ov0b8hMDCGFPigQUo5lHh/QBrBe6qo
i0luL35yWYJZCd2RqN8l5iC1Qbgg1A6jJBXHklXUIJ7jO7Oihs4r2dXqyOTDzp1EHM47f9fxDwpD
YTxNYSPqQLYIDsdDagD6WMAn5FXU60C34Z7DJSydupGkT7yWK9FEOGjFSTkgafivLGpw+C5QWqi3
lzhRYca6eWouphwzhYgrLfIL48+lxKrsOBwPy94jnxF2Tj4VdofobDlwKrnbjMze1eIIknbFnpqc
YvYzSdUhsY/gd8ida6F8pC6nDaQFe+KSe7q6KKzJVKwL1Yl75ZRSu+Ybp63Z0eEv0XLdUNk1XvEH
DX7zPWNAFXg8G/WLh/XqLXthuWcw/VTXknkXumxLB7DPPB4Mh9VBIWRY/iPaJ2HlBo/9vqunPbU+
8Wjc1gCwc3VS+jIHdoDokLQWstggHiW/Bt8HLRSvquxcYqhO4pBEtZRPGWLPvEYhpIvuueI0eydL
Dz1rvsBr21/mKLxt8LWIPEavUil1o8+s+Zk7d5LLiDW0yFGpEWKSqYkejyHO3Mtu2AfsysbDYjCR
58fPJcZoNfREiz1hJ5UE8PGVjjDDbumH9hrnCJWWgH8TZjcVs9tjRP8OXrOFgmARo9X/NrRAuYgK
5aC8EFfZvEIICEPJdCcJNPBk6EFErQKPAy97omUlDBmLRwbo6yS9p/OcPK+uw7+mKrPdjaQepaRV
8P2GPXRmq1F5l+DD2nvXe5nMXnCVZxQH5tj14ZIAPi0KmIQpkVFCnzmaT+ZubaoyBZxLln/bhHK+
LZ6hCV3WyCoJxdecosexkKLNu2r6EIULD0jhF0Hmbea2YdY6bAFf96YQ+ubcniEeKbMUIOvjr5YR
XeJ/aqROo8lULgl76XCVyoNFkN3ykzqpGVhhQ27vK2kDis55VVShvNSCRYJA6n1XQQd2XK7RbypD
UYzi+OXxTRNsurJrCbbVuNBv1hzJAvKtX1CoWTGkNaQwf+tPtNHUd5rgyX/SFVc0mdBifdDZTtXX
v6Fgk8Wu+EhFolV3omIhnAi80touXvAzFZo/2u1c5AtG9VHdLBJFnG3ay8ozDKkbT/I0XAPiZUOT
GhI4eQaoN6L0cFZK9JHvaTc1WMID08ErtIhFNvgRoDRKuyZFanv/8aWctjuLuF+klrLrdInhkg67
Gr8LTij+L7deXn06blcgx07KcESgQKfhtKeHVNKpLeUt3q3zdfQ0G9nNQLRlBrr3yd7+akBj7qt7
ydMzzCctB9c7fMBQQX/BahdF0SElo7kTobBwibwpXEEjkgf/LezNXjlaMkNnEMU9IvVbyakHgH4L
x7/8ytcUPEOQPFQJciOPOP53HaZ2AcXiznE7NK1SQyCO0iL4t6sasf/bQjNHCzEUppCR8eMGQz92
46eXdmYFOa3CM9vVemOflDC9joZPvfp+Vt5A9YT+EUA1hqsW6UShOTODqfJvGJkWsz2NNiRMDv49
hj9DAjhfakqViHg7VI1/CyKx1Q4rMlfjk4/1rR5hv1qyG1ooFU2TtDBSiGKXO0eDyjKYO1C/vBHt
KQFsWbwKcaqvq5Y8EhEAyRSIfm6G3U5ET5Oe4iFMTVb8L87bYE7AbwkztpjapZ5+Unq43CliJ+da
mX0l8ih5sn3fs5paxYyef+jvN03u+U73y5YgcMu1W6jOSTa2NrKU33OtGjHCAkJ+V7aI34tD2oND
jp1B/oFRhKkzmAJj35mzDqFlJwqbyCPfdn7PQyPwMugnSG/HKnuWjCxtU2ShQDLGr8S/L3nwoCwT
q5/9l8fxW/mbpGCAMUaLENFo45YJmQqc5AFgPmK8brBqDH7I1XaJTjVF+H1K5OG9yDwn7SFnxhbw
bbLtNOkLSvTdFFNUdiwZSppIiV5PATosE5RzsU0pccqas1+IOrB6WJFCDD3WinmMV6CW5c4QVdpv
oxGWE7zQK6ui6LTvdEbsth+FivNpQOgl096XFZ2LL0qTB+tBjhX5QrYOfvw3I2jZ1Hoj176X78Xw
yWu0i9r6s25xUOncqPu6SvPdTnV1mDuC7w6ggTSDNwUVnDcAadgBuPzLs1xTVrV6IBnRmkYKKwkj
7WzqrbKISAVJdAZpksde5ruoCWPbYffP+G7YkO+nUGdhiYUYraPgbSYA1jaECWm9MJdYBCF3YJDR
mR8EtRz8Gz58KrvhdFkkJbOwX3r5nJUJNQo7AdEsg2/6+GWn+OSOt42vkIW56CU076R8okknZ+lC
o1H9oRjBLYu9j238YbYhrRAXzbXBVDDAnoZ7TCdV94BskHoaSOQUSbSeR+76kmztZpBowCjr69Yk
oLg1Ham48IvLbqRm0v1ZbaXXwIgEcqPRS1NyYOnQPwwl0kZ/XiU9gDuK0Q0a2MOBWvAYBLCtf/Sk
1qhgXRsyMxaUvidWlSl2r8IyPIP+VeFDtRjsBe5D6f3dsl4gI6DKhSg1pYEpY/7eAyndHfuZZGkO
T8W3SdzFkY55DeEtSG7tDBORUAw0BEfZ8tz+tvy+dKgjPVHnmP38ysWxkBhb09aLJq9vh/j+QBTx
nR2uaYQ0PaTBU3Dvbbm3JbQhHSnLplZ5F5+DLK7cEZ+Ry/a0yRKzYq9c5kIVJ5bB03hkvpjL4+D7
4OqCVaN6DvsSrLLM524RmrjUCy/tv4ofi5ul5KQZxWtfQ7LYQAoYQuOW9iYNBR/PjcLVK/ZA0jr6
QkjXc9a0KfzbNQrjXKYDVSjWjlJeQcdjP4dmvfbKK/uP0iuhW2DiFzE52RjWRm8hAQcs/ahB1eGa
x259y0Pf/qxk5u/J8NZtrSoxv8w1t9b+A5TGEfY5aPwmdKHPzwsgSM4IZD7TllAigpLaYWe2rsmE
JZ0biq+CJVJrLhVWHPy3xAqXf3xPIaJFXLrh/0cucCGIFRDUHm6LfeVyNiyNY+Ze4LtAxF1Nkv3x
RwwDBHjLkgW1TfklGHT/dXA81svvn+Ev39S9qcPUDwlXsLuO1k26s4n/q9AdAI8Wz7gczxRrwxoa
3sEH8OI5roKsdvselX2gvK4aiid/sELavOi1N+DMH2HVUbNfTPHorpC8ejcB5VYD4x3OK2J+Zv13
AyNeNtQw7UYWIPuYV6ENK0aDiPBw1lE3gGsc/ocTcwl2J2GkVMKeEuzYB/vZcGFHhSk1OoicEGAt
QyvdnDEe+pv+NZeYd5CQpAYPovm+rEyJaymt9rRokG8DPw/s0MgCxSGPwMLjXg0CrAO+WmbiOGve
6vtIqwk+zahs5HDwzZ3iJWqmiLc4XrUHGItEcvP37agrvBwzZuk0Qd0O4wRg7y6+gooz1jZYoX+m
6RKcy5AGZonsw0qPqdT0/mEydqf7NbmepidpPzXf4ZjqAwmS+9PKHu/pVasqrLZPRIHcoAuZEyzk
iIXQlCNQqQlKJ1D+T/QGJHmnxLk2H1Y0gaYD42dwNDfsBc2vmsZrptrx84+XaSiE3aHo1A44p9lQ
RrciGKAYes5+WPAmw/lWYq2vcMsAKQXDZjIDfuvCxJKeDKn337p4E96V9H1qP1RSZw1+NGqxe+9a
5tpTqyKZfIfUGAP60/Oo2O4FwrxDgVgRN7k4JMyxAqJeVVRaE5jiQW4f28VBSCZ/e4wnwlQQOGSv
aaUmBwMiNqxS3YrClbkdUbrcaUrU3KDubyFMB/1+wBygfKUGyd85FkVfZwGY71KSk/DcWW9vQeEC
Hiq+0Sf6wNHWfILfiQFSyWvS9h+QJvKva5HKXLIZlydtFk/jZGd2mx0AK8k9dAHVGUc3OTYxA6Sn
3TclsuB1LZtr70Pt5Z+/xh2dnd6PVvmRdxlTOf1/Pr2qjixf05d4+Qx9l2vSEv+7qPJQXDP6ruV8
1omp2rXHbzk9rwPXMqrNT2iWGPHoc0u0DI2yHmGxu0l0Tw/jXgY2fn3foA2NMwtUEe+LlLKP1M8b
iOrJcguCfExEMOIj90r/tocgsjKwmgRCGObp9mnycFEWyqiO0T/ARysnQMxq20mBsDInbBk67gXV
/qGntmDaf8PLb0s03laFnTbt5ndhTwqKzz6iNAkvfcL7sONzhDMnW85nq0uYcDvMktxLvNx7MKZN
OkFLJ66OmPTvtRbx3CG5yjbL1z1/nDXSMVTNE0RwV4CzSWNyBurhETOuUEWIw9J4wYWWuPXrPsZ6
2jEmYRBiZOeVTcFXf6OPEs+ncBwVabotw9CzwKKJ2f6GbtflsAJSMWIg7nBXC1v2Ebwk6NwyaMNO
zfSnLvlXgapo6RoUHIBfqNkBbI39ubRijThj+Uqr5mIHyUf6njBqGoxNCS26xPbv1fKyd6SqVo1r
Nb1+ZNDfXsLmQM++ZfloEPiLtVtKfYYKCBKvtWGxFwNGYvIzYp1MB+29bkfstwVteV4cxCdJUUFv
77aunmRftOwMs1LuT7vR2Xk/GzKmulnU82zXApHknjzzuC+bN0vk64Q36LAMk2hNcgbSylu4hiSb
KMLkzbHJGoQi4hEyvhxO5Znn6B0Zkalb2FTk8yheTYhDGrmTWuXmM6A27ZMMW2vxNiscqRJ2l931
KgjWN8fxkjqJ6+95lcms6NzRoSdWqlPwjS65daUhk771cu/b72XoAJYhKmB0mZ43RYmWR/nxqG26
CjXEiBYUBY9mEeDL/NzZNvelXnuKJb3W6VPF2yGTbcJZsLkFdrOSPLyfJqtXRPULjU+5FC14UlIe
E09g1gazpKuFFM00zmMfnmQ8UJyduBTdF9pd2+aIBhWH2Ma9A3U+ACH9FIM3boxz2he0lTeTNAdo
cqdaUmroh+y/lZ4RungZ5sbsfNRT1cu9+KeaJVtQz2REySeXhZWfHzwuFunjAGx3ArsrExlI9//X
bGKC1ckLf+TZMmWK7z4tEZXg+xkqJ8ax//xojz3JIUhO0LtIMfUb4yJqmB1RwFoYElTDktWozBLw
WOeHY3j8bBUTA6bpy2mkY33D+Hg4i9T9wrahkI+f2eLrgq1xv7/3a7uz8MFpRRALP4AaHatOkLdG
+ULiQdwTP8WA8NgXyPe+jk/lfcJbYPdB6XDo/2nCfW6v+gWNq6EVMK2GYHpfPyOb64KmWdhDxqvO
ktHUROKTejby2UHJe8VRUaQ8DD/faXaG9E/QRIaRQWBlKYsVvGVMORlwJNNjb1H4SZXe1DXYhcVj
fM9MUYcM49OjnWNCCM17VVxRQnyOTzDwyN4/swUSA7EEIySdKO1PZOEnhfAUMarbYO9WbSD2laop
kTV3u4RCO2Hw5y2icUPiRhjZ4YeCVMgRaoswgS82aBOpuKdaIIDKtMth8cfCWjRSUlg3OzYHjyg1
JEzW3+evjSpZLAF02k7dz9fxCZE1Kmp2EBoUAs8h/C+VYRO77qcr9/f5AmMmKy1lx69pnw8J49Pa
s2Xs/qSGOf5L6L9vMnDgur+qDb9YG1z9OMy3zlwKUTLNld5Ud0wC8UB7rQgvsN6ptFLWOG6SKGoc
DVIA4BhZlOXYwthI5XGNEwCq3w7aKxikjIPsh5RvYBuzs6o5oGMxij7wVxBmaCgr+exy2BUnj8S+
UZWdeCvLGLsg8RRF3E2C7sf6550URbELI0E2jGM2sf5V0A7f/3npsJ6TiJSL+o3Ge1y+sIP5MDTG
3zwP2ka/cRetBcInb1ybjqIIztxsvDPHFzE7jQmw5l9msvOrz0MVACKjw7cA5R6Qm7sAAxfIMWFz
gxiEMyXQoBDAK5GALAeyOh5ZGPZBJfsIWSAvDZHO2PzdM9MA0fSE4/VyLz5GJMha2R8y7ejhpDMj
e6wWYCWiuFtvcRmeO0AeYf8V7GScR6cOAAqKMbDMooUzn5KgFHlrsCWAO8cIiFGgIA1mwQVqUcLn
WMxYwhY9jtyzRT+gt8g/NG9sTTLdS4AFr0174o70xIbnRXhJuR/uBbrSNgyLeDi0HWS3OdOdzEpm
6mnAdOHG7itDQwfdzYhljnfkSGVPmX1qUuC9P+SdVghPnR20ECBB7KwD+kyT4aYD5lYJWvnh89sf
LDV5H+VuLxEgPRBlHfNkP0pK1M52+N1ycrICz/4jGPtMrGJz/IfH391zFqZTHo0dD2fAuMjldILA
+dcFVk7LzRbkVB+ctGyHVuLrZCz+vdByuLyx0+mt3C8rAxLeL9nHIPOOVb+q/tWAOlr82091EXwH
2Yz8u+QSKrvywqtKISRdSIyqO3BQ/AbsAHHyxTML8zUBH2uk0UhGfv47l9qzbDPXu6jiT2xEehKh
BuHpDY4La/VyuxiV3E7ziiwTjj7YxOWDnVd1piJJ91ooQ7lmhjy91epF0Iei+JtaLd7AVsPjPmYz
iOsy/+4pNu4siLF5l8I41QZ9F7Zeo6vWHC1kPGMs7mHiroFCaZQlpiUYNltSEOXjF4j0idPqjq6F
XpfnvCH5SC0VpyoQKIO4fi4HJmlKfMsJDZHIm8mFEU7dGm1XUyqJRDbM6cnYZoxJZWgjMYiyAOCF
ZL+Omue84Rd1r4w4Ts/q0o9UiyZl3gBV9KCC2m2XQaNYtoy2YPguLfDlc83yEhEVA+dyahFehYpb
Pz+PG6jY5YKsRnraH7wZil5FXNvfNteXN0dsWbvfNNFx+B416LuHoHqZEM1KNHP20f2+G5oZQ7ih
y45Smoiklgy69qVK/UJTfafR+pinDN0UYXcYAm+QMsQvZ9u3UQMV6D2Yfj8J62XY+/x0Vs42cVAq
5cmxKc+/UY8wyeiEb7vs4PcEwxcuxPunyO2gM+FGITtBxO/GtWiru2mqOMMyDf6hsZqbsxjg9s9n
n193jLI76aBPnn/XBS7ujgSAGa1jnoQaGCqSHqXsAqEWcDyVoFAEnv1JTnqzpX2EeT4O9aYB/3vC
43zZh7CMmRoi/vja8du5yXFOv0Aj2Vak6WKbZfWxGbvM/zNymIFOVrLg4a7CtShLrmG0K+QODwDz
PqiSkG5FBoXn3upqdP1ac9anckZouQyEn3Z4ZdBJu1ACsBeUIEOYfrFlqTRNNKvFGodTugFuULp1
JEjQcC93+3TCoX7NniTY/mbPsRzpNl1Cu/pLUVCSZRCVcw39KlJZM1nGN2AU6BYZ0TZgGrxIW82t
iT32ZC1h/ETRrnvLPa4FnV7odD1KrXNo9q3lRCTIi5g/rAzProJDxCcyP7GsEzXgAo97MVktTOXo
PlpzlBh8rXQNqOXhZmv/VI0QaZtxhsViozUFbqzAgQ6fz+yiptEhr1okrLYElVcy71DTd2vEo8L4
26i7iiHjaxi+Koq0l9CIG56uTcIB+0YarAGNHkDuXsRP7g/T+qwKwMNGj4v1tyJmiRzsYh57DMIL
shUXGKKNYynZWZMILE3IhNs3SffSouJiSMuh09hd21Ywm0WSRwvFDaTn4AA8Li7lNYYL1iBP24ti
AFVP0dx1kA40EWAwQPtUGERMIPinxfEOo5oCcyusHAQXOTkcEL/EdqPc5BUdZxn31Le7ip7yh0ou
vUcSFopQJG5d7sDVkFnlDBwds3FgBHxNS9Tw/A0g9Rdp5df8zEuEo73dEatrhRQ7XC6mggRyUN+V
TVoJxBRM3d3pYHmwLkFxPC7tJivPolKhARLuf7qUfR4Oho202LB1KFTQpmHI/C4/Bba/1dTIIWu1
T9oucNDA5IlsDKr/aH8n9+rs9PSFGShuDewDiO5TiUGjZD6Q5iunIXQK2nzq4tYKjcgj5/1s2+S7
uJEQp44SikhPAXAIsPo5qrgMucowXPDN6hX1rBoEvGEuf9qLTRR1CoHPjSJlQK0vYB6v1HkxCCdR
WFNultaWZmEumiofdhRpxCivXtCqYDW4RS7uDG7jYnXg2R795YFN9EkKYT6Dd8XsOd8XgbZ3W0r+
j70jmaimG489rM8Yl327an8Gq6frYACpXYLGwyRsW/hp9Am6aJTlWRYlzd02Lql1jTROqfbZn3IV
mmZ+2RLIlXotAOmCuIYCVC/FysJlHKRHUR4GibjL6mu7kFmpM/K6AM5jrBCRu5sl2a8IFXfZxmV4
i0+Jj9tGxDK1NVvJ7EEho6ygODWBsatxYVWWQrXEEinX64gfMWsRex7umpcuQyDszzFssz2y9uI8
QIZlbH5OrAPD8LLvLg/OAq/zux6tM4Q5unvvza+YzKnAQxgDIY+r9jj7ioMn7/KEmchOrtSVbSpz
z0lQOFo+UIpqnFASOAf5f3Ir9xrYZFI724SAfZxXtbjTfuxhzBnq075eUew7a1HTvzcYTqBk4WM8
pRKv38kJ9P4e/lZNL2dYWhV6CavN5BgcBmjV/zaji3aEbI1osu/ZI+uQ1ZyDVQmMEcVixozgn2B1
RXCLpi85u42IfKjh13TSmxqP3SMBusY/fhBmxAGvC6RPz6MmmJ0YclOFLkO+gQCiUDCeM6cjpCe4
HAG54U0X3nUlY1fhsfwSj4tGjyYvfVY5h+5i2b5Umd0CJRyVKVQX1HRzukyM4MNwXYGLEq2ph9wt
BHpA8MuiQT/eW+4im3F6TJoY8E0cPgNqc9ZygRpbxvzprx1hGvDIyAtHyrMyHmySiZYqUzPOgJCj
Ht4CzTXsFZ6tDj121nl4R9dFUrNWd7lBySC6j5pIY3QPywIws85kOmGBCeoIe+XiskQ4c3p/RWC2
4kMZ7J5821EtxSYv9Cj9WSEGE4dO9Yc9EH11puwLQVSyjj2a2M9pNo+SaGZuMl4xzSb2TB79CWTC
hJQsJONKU6lPNBx2B1n61w+PkWay1B3hRChb/5jaB+Lg4CDybrVh658wrYVH3TGRqs5eXF1iDl/y
/BEZznerYcTHY4FejQiCuC4OLB/dli9ZerJgnLb247wn91cpx7oxlvoLkvI4FdKPiEiXJ3Y2Rccv
cIrmPcLtit3aqU8y9GB3JZpzGpQdd9QkQBk7Rc2rq09t/ZrIkVcfE71Bz8j/EsNm3DFJPly6gKF9
wwLW6Hb+8cXQuaQt+ecSq+4Q9Flzm+yuzYxrCblMGwgEcGx33S4ZTlbRjDSMgCSvP34AnoeIqLJ5
VQkhIl15XnbnebHtpvNwarQd7XfEX4GirURFwOWxJKLkO2HYq+R/QYRZ4H7b8AgC5Um1HW/qckPs
fATQJ0IDO2jcKWGoeBe5CFj8yFoa5rmckpuQrotqoWVBVGjuSzKwiv8PpnG56BwhYMsRmS10jVVq
JtQ/4WRmSXDQIEvHCcrAOZXm8fFjOt1zgzolNVnQH/qe5HekpPYY3XuJYlMdzp0UTaxgxdMtDXG8
Rp9o66+k/t6b0zulxuu6mKsIQHq9wvYyxaudkdKhxd7AsBA4GYDN5dyrt4yqSO6JjohvIqxhxgh2
fdmlQtgeKeX7Dj4jjyxeAaVisrJVVPmijl/8AGEkuzPri41rtNzsO1qfWs/7X5MTGNGz05GvbFd2
DAfv9AwIdSpbApHaYfwfxuH1QKuUCGvVDGxifmq7lxQgkysJmjmmwHFbsJNswvcBREPTI6kLrLSc
roqmYfbodeuMu2mLbBJl46s6Gb2RvkrrUqChPBupacZyHUrptAGOIS20DGNPooMc6ZVzQd6YgUju
r/XE22eF/CvijBW8ykngjs+jBmb2lbGm7RfAoBdz6wKTT6CZnm/4t56rSLr8F/ZdBu1REs+NHSVE
F4i5o8LP6EO0kKhd7puZ67aHumJosi7QHFTi76KU0fGPlRKYKn97OHFcLm8LJHZO8muBOhWSl5tP
NNyn1BhnwJamhlqYt4LZnuOMB3qbbP5Mtmm538EwVyPx1CokyS+AxrpKxBtLuG5Ev5eNVR7HMpVY
8/QN4NHLIabUFTIIGAcH/5pPsWB2Cf0+e72Qlc4yFqs7RE/geBONBwNy+g1UJc864QBkgq6cfQw4
CXoF1J5cOiVdip4gwHEcVlreCEu/GJwo5BjaEmAJ30lfJHqPpH4u7Qe3r9YIk/WgFh+WHIrMPD1N
sMB03xsPCmnXHzm+Z8IuTLAUWggXm4bE+cyeep6YtuBa2F4thpYcEjUpptJf3lJcuu5AYwMbw46g
Isl6ep8CQS+4OZhwRJCxfFcuNGEa/Jp/yMRRD+V1KdsIsmD5OqnIYlrNlUVc7fWHNu92El930eo9
CKPHi/HjWe14wFddpIaUZT/In9jYXXhc3CF0tj+29pYQPPKYIw57SwLzHh2pztHx1zuDpum2jlXo
1lefiwLG87iIDw2HzcSH/89+Z05FpgAbmv5RSaEuo1oaoFPrtQOmevg3QKipq7d1KtIaGZuDKrxz
07klwg8XfdXehu7hcLR9wOcIwkOEY/kBCqk3IRL5fjk3xekwbIgsGT4ZU3609WJHkZVZNvAmq0Gy
pU7pqCsV2+h5dv0MtwzYyV5a86PDd9WYizpBcblEE5PtMbm/hi38iU/mE+5qRGSdNkpNdbSoQ3/M
I8XVXmwmjuWSTY6/t0n49JSJGpa/tidjh7SWhJLBtWa4KkSnAneCjcXk1Qsd1yyoOYhHcBvHz8PS
hW50664zNIPLTwtkPH4ZaKp3wcvdWCQoY3augEdJYYFmOUocM0NgWHizasuNeKt7KWeZ+iXnvO1H
M9PIJTh/312Vh/JW0DBmnCwxjnNmazyFVw6QYdaOMtoaPybqdFqP5QY8d+5ovB0HmjQUxHCDXTx6
BJDCgMEMLLgBBnl63SZharHu0wnUE/Zl246+5we2UdHlNQJynbLvyXrO0WYGhHayL/0Ky2Gdv473
iDXNQwoMnaDNNW4VeFR8baESrG7HjjAjv85T218odA2h5BFXfAEopUnTZGvYtSIC2KDVnSnCEufZ
auJKb6ziKUzAgyQo14SZIpX4YvoGSFlMW6RrsE8CHbx5D5UzEo7FgZBkdWSz/g9aZ++ERH9LuT77
B1th9l8WeFCbTYtjxirHHlPAi/SK6JTbf8YOBhmtUNRLb5HAV01f4rESbaiOXxBMr/zRECaF6sJr
7LLR8j4MFrmasijBLyEkqcTHlvtMJadbLgEUyI2QBz3Cnki6qTPSipeaTumUEpuwlfXT0xG3EqLM
4KNXEOvS3fmv69Dk9buzxciw/dULSNEcXPweF8MgPc+lDsieAloGV1Aiu75Cwri74v69/EYTHen+
cqbOx/6zI7aj+ERG/ciTHvM5ksNTJRl6v+C2uc52tkKnlllYJOl21ywYb0U6I/QPiTzhUGO1t1ny
8OiplRsCbzYp5M38t4WuS/ynf3wc3TfB2bzJCmyQIYNuBgTTsF4bkwdNVv+cONu1/zRQbErSEWYn
crhonfHfjnVJbXOlR+gUTm2DXRt86mtVNXCGCa91aS3mecOun4iJJtCweGtiWBRRmrVWUgAzTCyG
SCa8/n+qpPkM1JeL9XaIdslXeIqyfB8i2cjWyFXzXdXjUX2Z9cZCXCMVQcedCZw/eIbl1CNs6+ux
4OWOekMjvN/4oX8Ts8Isl8X4JtcCWWKJcAvJfZ8LQD87WZ395UM+RtzBCsDmFr1yPiZSipe72T/h
NHNiQzWDcIIl032RXEUPJDk9hfy/314asdNXbZ/WTnUf1FjeZKGsfEAxjhpENGhTQ6lLvX/hN7BD
ZYPYlTC6oYbTUqaGbPuJ3t7LIjMo1YwRD6KF8YAvHn0KIEjjWBqFigUCXivBaeFS45YeYdmJqMas
f5J/+CwRY3hw5fawxVU6hamSIb3wYphw5yhTxvv+8rR6Kl0K9OBpALGf907mJhlc7Ud+cHxZqbo1
BH07BT1oAWM9tNr/4skY/jSadSft1+VD6ramg/QS77kCwSV0c9EQOde0aK9WwxNkHgjNSBDZxeXg
Dl3Ujgul8tR/pQ3KFIQEbustlSapqZG3ixw8PiVi3+AgOMBYND6+dswEbiVVrNuWh07RROSyrdp4
iDU3WKSXh0Hglu8gEiobYzonFIlhj6F4hX8WWIgNIVogS6C0/1+XPkkkwdEQiag15kZlZnvS+YNJ
7I9QW/OXno5SB1Y7aLZAUfzHHgwYxEtL31L6apwfHwREdF8kve4tRhJ+XY6xI/sFpZbUQZ8inFWi
qcf3Jhq2/FhI4fCnO8V609zDnCDAH+4MJHdOxFibsirLQeFdWtulQxwPingTZHiHHUOoLdD36i2S
uBIy0AV2AsIPzytNGcvxA3APhvyPMmtPsPadDAS5k7H5tUoAtjOd/COggf36FYx+QGnJ8s041a7P
D8Yem1LzXtiqqP1wdMBGLnYjDjjQTeN4epbXXWYjHyOrO5Ufijm2cDyA39M4zat380n0Hu42fslz
FnP3QSq4Viv8bt/o1u2drZQMU6ypoX3j7iUXZrA66340JcxgGCVB+uHrspbXkllNMQkvZw9UMcqS
PeYteoVB12iwwH3LLd/32ZCkhcxbNG7usjrk1hzNQ7TfCB9+TtGewa8QQSEyrajcJOQ8D9y2mpG5
CYbTYIKUklTzaq1Qfk/dRxeleFRWoCsj5mYHEasWaBFEDUK46YTBrM2Tr1mnAQ0w8lI5opWl2PJy
4utaLUGc+qXMfdZsGDFZ2nR3LJfEJYCZn7idtQqVkqg/ScnodXDUuMpXJQxFPeaRIl2+dBJAy1Pi
Ge9D8ySKe2LqC/rzGW6gZIpDl9f4icOsIdk4uV8PHfCVIvv4MA/0WBnxDkRCY/meKJwRT66Afkhn
W0vk8djfBYQ8OekAhQeUNegkrHseyVUJ/VUVijfcLovJdF5+Az199YFY+jYHFUftcMh5qHzvR9L3
sJXTvm3B1IAbQbvFK7lKs9ACIidwJDh6rIgnDHe7pDQ1xMyoVUK75lwWMcRtAtusim2y1GPWxFwt
Jp0emjMv5EZIiIbtcm6lANbuBv+UU2acHqUKU5psnT+2YiXdtgQBpPWCfhMzcmXgiiDoEKLMcuGk
SoOEoD7fYkH6KRBCS3CMVjLbHjj5YllgM2qX7K5CI+3UVOb6R8CXG5jjSovLTzf+IoD5CEJL/lSw
tXjL0UbE2mxxqfD3xy/hESfs/c7c3KLBQC5nGcjwynJuM5WaHXWiYfZdaPi2uVb/PHE/Fc/yS0xm
zUkPtXYhVWeyNah4irfdebk7r4tzwb4cVINFkIFSkKwGvrx5tsOwLWsGz24ktaNFaEIoFm4BYaHs
9nyxr8xJNEsLOEhMa98FFfb+q597HjqCjKxR0PPgq+kZyOs7H6Nn2xO4wsqtPq13Lwex0L9M14m4
PDIrFQixRn/R3o/XmAXA/tqq8syRZf8aaCS11O+I+Hu5HHWlL0Wvy9Pe5tTGf6aYI8/O/BQdx7IW
RdL99crGHpyTVziugzCV3i2bUkJawIK0LnhKkTdbpSL0+oX9beshq2xCop4DYPfOPLDvMVvzDP3w
XeTqVVwICStrZGbSVeoBozPTtwCBkEgTDbe6zo6af84AMEvRDf6tWNwU52pHu6yZYhSCdcY8zEhG
yUx3qbA/qBHzH1l2q4KfVjcYa1ysjUuDDWmKt46EHtn34UcaWMyifhBNHBXwYpofA6/CPL1HgsKW
hzV9ZTuEXfxXWgHZ3aJHkyYVG0/PbIMWUKXJrfRlfqUopffeErUa+yYkmCGvTZnn9e1YJQMWUXId
gTskEdmTeuC6T/CwWP7cs3CDemBzZ+W5eRtPkQCvz7rdTVZOpJKFwZU87EDK/ndP2f9Yuacscb/a
rsjM5yT32qwfAWy1HiHPk1UcFwRTQRsCz8wKFRs/iP+2HxXVClupk5+7DbjvdqKUePXTOcZJeuph
LC4QOl0d7OpPaw3XT/rJrkVZ1DVNJxdcC7dFcYX3nNEa7ILzqXAVarua2rnwU9YHCnBB9OUc589e
X/cNUeUPBOiXjZOY25Uw3Mpw46Jvm7cOhPpggdeVUOaDQR7y6JNVmgKO9VZ3dp5n6sqLZO58yGcL
acCTCOFR8TzkLsgBRlVNrDPYgDgick8yYQC2+CKw9EPHavJKLvLWbRs7xDCSFOlZkNw8Zu2Z98gE
+Lc7hscWrbUSXfBwy2QlKoWLGipbn1GQ6M0/h9jOPdvFoM1g0spzf8xlro2xt9on7Tw/zvSS4Ewy
lEp/03uwIEGCsmKGFJUabZge+QerrI12nTU6T2Qnvv7AhABa95C8InaURUDYptRMs/rf/jnvOGbp
9BHE81VsFNKP47W/5KWYgtFYz4NpWvFBvj9o0WbNJc/cg2QrSOKXEg8UkA8UXOUn4x/yISWRut+B
if7gCX06272+83bNsuHT4y5FYyswMZGnzrJbPRBAZRLU3nOyah4UtbSLv4GCAEgPqjZ7rRApO2sR
MxJVRLK5rELIj7VMB5+HUaaL1TL6TwaqvMRacGYZI8V9CeR9UpiKrAaj5lWYVQ6/Imyr6Wind1Ej
bVes8UsKbqTKTremhKjDHzOJ9q691hmSglmUiaQPBjct9hMFOXQ4Y48st587sgRIBW40BI0+nJdM
8cgd/pFPcpLSy1D6qgF3uqqX5XVMcERFXLjahyn0bex5yTB1vOgFBsRydvi0bzu6RBFBcCU25/KB
Kq33FNLapqcuqVgQvfgfVoU15KEl3BnwWx2nbtjeGhS3iCBuYRGsijtUGyo+UwZ/vrPs4gfZWDCR
lBF5lcuu3XTqpbqCswOVi/sqnoAcNy+5mt7H6wbOz9j+FPIw8xv7dlykNlnUDDCZYhHhueYVdTA/
h/n5z3dNoYeyhMPW/KzdLCx2hNgv5rTuRaOmFUxeo0sUcnqPP/gv4BrRIpi/6Q6Tnghn+2Nxm+Uc
xTmkjaK6FwHQfXXfiujK70AtkF+kfS/mIL8So4MKMXi3JIkT4NUNtGBcjDbm0EftYITLAVGRpysZ
DE0hGbeKPOarFyeU6NSnerJA7nwdxnjqj5WDg8BGOOo8f7RSXKlunlBUH/SosXYzvsbblDApej1o
cE+kMAEZ1hZ11r9bz28/zUGrGzAJtHPhqgFHV8MIRSUGtG6Z7o+Ssos9/djG4N8a0ubEUcFbPGyk
DAaNjgtUx1u31g7H87dhK5DmlP0Tmjq75NokZuRCDfQDmquPR5YZ0qy/klhIkKvgj0oJqj1vozZL
eCxsrW5GDAf5OZq6uAJOqnxPNsMr0XDW3f/CJ7htHuVHUQlUFlapxGen7OB6/HYEBx9mx/SROFUm
0CI4cC8NYWGewqKYtUjh4BqQBMv6URPuM5334Yfp2ju8yrrYMN2xD+G1vnrR74KmUxKpildPiDhw
vqoNxhpdY0xsYjikZdYTQPFH+4fg5HVMsUD3Jro9NU7LYyzEuq8PQ1tklAn7bMgZfQmZnTh+hHb6
kYwKYN/bcnhj6aPPJGLWpFAqyzcZgGjbl7zVUQbzLEH+rkcLOjWWjvnpfT/i980SN+LvBwClxCF+
xSWXp+iViOSQWgTNFYlUkFXlBqYRNZ+il5DwspjDJKVTvnL8h8bJ1Vs9zu4d9fKI56w5KCQ4H+tT
8KHzpZwD09HF+SFHwLrbimwBBJrjw/n0nESX+I+QLyBoRgb9P7w9rhc8QY71fqm3j2h397Sj2AST
DthbsLyEUekXJD7Q5YldOG2f2CycAeIq8u4xl4FtcHotFdIRovPg2ha+f2VOFcrD2Rd2imZhloMh
MRwkQJ74RpH4FGaG2FF3PiHLhd9wTTcEX5k494gjW5yc4+a4oKPjNFXtKbEnh1vWSL7L9XD5Ah6b
Ss13+8b4X+P7M0A++zXg9u3RGtEQWvenAWQ6uf0E1T/7n9CWSBfdRc3rRj9xzZiUq4wUgRvjrv9l
NrKM0RmiDuQb54E+3CB8rmTyEvkB4bJJ1JX4f/uQLxC/tBPHEptq4t3IKgTuXhSG2mvaIcmmrQkT
CYL13GhKNBZ8EbyT4oesOask/Nut2blwYdVRjObk3w152XPlpAoHkF6AHFJ5CRih+FPQgoqRuGak
J6e1mPNRoVY1a0kDMwfz6QrXk6IPuyxvOt46BIBfmFwEPWprOExwiz01jicCO9oUWHHjaVv2Hj/R
hJIbfnHwcMMulzdWd3bGtavc2q45LYmWSjfeCp3hwvOdwSXY/oTCHbtHY2/gFWia3tJtDFODjDly
b7r5lMGMeTMdrDeYhbXg2HDXnJv76IV/28aN6kvBWZDtssFhWlsqTqQUrEFvZNZjsAE4///rS5tf
7Kdis3v9y3suDKgwV4cKm0mUohWFS+NxRnVrL/Rd5wDjdgO6YWwP9YfP4XG8pvMMtm/X2XZh6sJz
OJTcU+CDUUsz3BfSXIvtrQg7YF6jVGBsKFFu2AJRh+p6u3pdH7RdjaDYfFtYQd70Ribf2JlogBEC
ay41m1MtLjLk9jN8E3d9TbFSx+d8efBB8UUhh2fKkwVf9y+aXyXvS6SUn2U9WvwjyPwHYq+JC3xP
KFbmoFE5kGpBAHngiz+/3eNLNqRUIXYA/b00X0etdr98ONb0PulM/DpgbaQCBeB8HwzWadQ0hHWM
+NDCmdF/NJLnNesMIZcCCdU5mRGB2W/DWC+e83HRNcNliS+mq+wrvjGqu2A0LTtHx62E/zu48MOq
zmdo75QCIKJQrWVy8ODHg4TOkHnS6uraWZNRy457ZPFIy4vaQs9bucQIwoy1w6zjQ6DvvoZsNg0C
Ld0yyJVOuUDDK6gDhFC0iK0n0BwEgnXJGU1YAgYomJCu5EQMgyceG4Dy0qkkIH6U5S9mrfLEcdgg
D6M52LQ+H4lwWXorHnnunAGr91VkR1vI4yu9mz5Cu5e0G0uOhuhc5AowXFWOwuQn77o5EoWwHoDp
bA6latn3gjfv+F1Uw7GVTIJ0ORCMuEg6W+1I3FU06HgFsLJ38T6FBxf8CJcnXBqQmBTjoMbnQTwF
6M/AwexByVu7STM5886qGBuDJeRvihIktN21kn6tsWmRdZxD6GEIB0HdH7dsC7gsDXt5tcQ2z6ne
gL+b/dQG32gMZVH60lj450JlizF9McVKBKEOHJc3BPlFuCoeZAgQj7+Q6/LpWLs0s0hmUAqe7kwz
BufL5Go8o0hqe9xAt1YGvXcibxgRhMTg9iMP8S/A6LMkSRVF0vjIemwRcWugIIy6f4WH10hheRDQ
0Ipv0r8Whp8w6XxYWDG8FQpsEiyymR4n36SpqnQcKBXZJeEsaoMDm+gOjPWqHKsu4eZoXuAPMaSj
zAXZ0igGlKUbFt4HD9y+mjX+Xk1Yi0rTYv3sEXUpnpNc+QoVcR2cavKscHPo6WfwiUnkhvHl7mce
xxDJhCvGhOxj3o6F2LhIyJYYXFnkZ2OorgUZeFsZzLIYSh8UwZixACVwTBB1OLR/UlzVRLZxIFXl
+XKEy8APfjWIhIH2A0P5yCn92TFK6NnqtZ0fz0THPf86WqfKnyp5uLQhi/a5DT7CHqH2jbf4GdF+
TaIF62Oxr0r5Ah5OBfu675mhW74dzb3lue/8Ny/cKvSv7BN1qbkKplgY09suuoayKu0vg9t992uU
i2BQmrn2/pFWvAU4AqeUmVFO93VxZvJZNekYRcDCS8deb8TrhpOgp3f4cDy+1olpblhKmujLCW2P
1TupXBLS0HIri9YfogSb4wkse1/1T4cEsnqhj590XoDHUEFYf57XNvkVs3EsmC4LiTASvpdK963r
AUpqUE1qRCNjD3XJzQudgvjbxpKPZLIag3TGv4MJEH8PsL6K2gcgvdPDInDsb3hW+ES2yVq+aHFO
u7Epv02s34GFJbnTJLFepsys2/UaXCy4rRzGYXVjP6IJWt8RV2KKsuzkxRZHsnPRW0xhwRwLn7Bd
y/I/w/t+NmIDloqgTc7ZeqaieMl0djRxaCOhIGb7m4PL9jqChEIF+vVtUBaxLCQVLnsioebR5eXZ
cK6NvUv0QE4kvnry0eJVgQsj7HdAMCZv6KL7pNKZ6RJPhmVtWQ4r7x2KsW6Y1Cp4bKhY8lhbJT/S
y4oox9SHygLhrIUw3sKKu5c8RHyh0nHpRFKovPdqoRXliVXvnOTjUVa/rwSOgs6Qc7OlMrhlYa1g
dhPNcs5QMUzstmCUgmO8Tpo+teCA73LRP2vlcYz5VX+vKwk1O+FLwZgX7AGDrgX9LuIeYmlEsjNP
o5F0aJQAFdmvqLU1Qa48YPWTvUPvwA68DGSnPkBjgW6inusnl7bprt8KB1eEu05dtQtkNGQtt4bv
ESUtcVrAY9G99gdsKhiceEU7Ao7WfP+B7lkTD1yI8K5nr+ZPWXIjuqPV5Rr//uZ+s2d10wfDd8NK
LfdBdUVqMmT9VFrLvmUft2JRZ23JXnSWMH+F8EU1Mds96EPo65hKM2Jxh7pPLHxf55IK1a+ac/A6
KR5iXYqO44Ti8dU0oBktG0LIfeYwJANzU/do6RhR/p4NNRIWvk70JQ96a7K+OdJJ/aVaj6TMtNNX
7pTW+TgKvUOam63wocL45DvzVd+rDHOhbwVJIk4oIAzHmqq3UJP/gW0UlZlM7+4i/dZersAN4e7f
0v5jHdsfcqyRmfr5MH/PvCizlxZLnr6QulZgOVSgdoU2sF1sMy63X6G2cgKQBiFTZGkl6/55CkIX
y0UI3Pw1mMptKALlzL+QMhIpa5dAs4e2X+5688PKYL/hO4RqQ5DPSEYwh5pE++0WoI0wLLMmn0ss
sXVWQPmnMVTBW37timtTCW66k5RgW8yk96+9WO7k/u5v9Z+ttx4nMRkbYZDNTfCxauQfmbqeursn
VK9BkbaSed4jkxfZJXpPNyFQpnBzAIHLeRsG1vdzLRogNacZy9kIuNsrqIyq4fUg4jfATXOJi0BO
aDJ1kxKETmnsGhB/RPl7WipnonHlAGzYxivt4bk9kN55Y4aK2fOo91m/9NSAHMH4VZVyabVAk6LA
pJtcMItF583igvRSvkQy66TNMqAeakOw20ymU6FiQbfIzN7USkd4chlCtMQ0NdH2fBjbmBOg75C7
RfmaEl3tHSV44OZNipdKUjT8eREMa9C01zMnyxmuQcwr25IN7UHLvZjr/XrVFaLiH97Bwg/0nvq9
VCGIO6qXGqq5svtUBGVnBVZVN6iRs3RnSf1zyGd3dwwHxfVxMDmua1MQ6AWdPNBVrJWhs7F+GmrP
yuT78S7RBzVwWaKitg1RcL7H1mOkASAu1pEos1jwya/ecYKTnFAVJ8BLcVHtqFtGJzUdLts+jJ4N
fI0Lbkl6XEXIKLPrjQwj/U5uvJkiDheFVj+8qCBu1JZP8xGV43OBdkWV9LaQkAchrotJ84sq07uf
MVJSHhtCe7SEqeRw+Kk862vnVVRYcX90OffPtOMb/gESPdh/lACYXYB5ZHFpC28vvlx1i4YS9E3n
uWVs1zn8lHbfiIYDIM7dNhi/Uw+XcA1019Psz+6KytM8j6sFnnLH5dXRDRucoQrgtT5xAQxeTs3/
gVrKDjixlJrYhfJ2UGTmxFKQPRjpFqGOxNQtIhvQp3DvATLEthYPRdwxkzZ8X0YUny3d2wl1ton2
AdxRsKCD3+YVCQ65a7IkMROBlspa6A43J8+jBnv0BwY+SOZsb6Lh3q5Km0EcOmkuTX8pBmTamZD3
M/nILNl9LPH3YrR2he3kS7IRjupzo9UES1L5FTi6GkZ1LtvdjN32ZIjD7oq0YE5Jf/c1GktdgbT3
r8xlW8abUFNcAuYTFgByzNzpt8BlR8MasnZgKMzzUhs8hUYpkqibGXNmvcq5wd+R+2PbfTRG29fv
ajutSaIQoKJOhDJnVjIvI+acv2LBjBVCoQZ4wv/9+a73EaNzm0c7BBNAoEBewv3h0y0rUNithIK+
zO5WAaUYom8/vgSa9sdLQeAYI9dXkC6ZCGs0rKNiBEGstb9de7UkuBYGcmNur5ZP6D/Ir4qAwpI2
St8rRE5oKKsqntEMF8rxxn4L20cd6lMMrjLtmP3Zq8TrIcFEFfDzpVeqwaW31sSVnVAjjO/UtWUt
OuKoTEWB6CLsyCQ69BbT2O6Typ9Pky5MuJLNojle7ibkDo3QOBKlk9LVvKn74PO7NaIFEFZDjPx7
qZ7FErMqxSIaDGEvlDyfq2t6WJWuRjMV2MIHtVeELRvzbgeufJD0to6PTg1sJCflXAwKhPuxhsUU
zfPPtuUeopfCz3uRbrhRMD5ID0wRWfhNyJ4RXppznHSVDv2Tu5pIoDkAbfuOdstmVsbVr8t+2VCz
TJ6zOrQ3YCRtv6nRkTiKIt0q06LjQKH51pxy1Y9le0dbIfzHTviDanH3+leysGlyWPPq63L11GOD
w4jATtFKlaHaYUR2fqzqBkn0onNIJxDjvkHocMxvMUxE3q51FLQ2vSKU+r70tKphgA6pkSf47jzg
P0zXjKjj9X6l/fZI62jijhcJ/mKwVJ8aT68QNIx044lPnaSJIojYQdkraE+LGl9yCEdNCZlypK6Y
oDkrjtT5Iy04q2qrZzKg7XJUsmTbSC9jUHF2zacQ6Q2iI6AiXr7eqGYNL+xpc9O+h4p7TXbtSg8M
lC90hBiETOi2gGV5/95L/sTKF3qw+dTtj0caLiyU5GHVpny4YyhcdV36yuGdcfS9k22Z7dfmi0Yh
/G436uK45LxQKVu74YowDmmnwrKyzv34+DSaAs/KVoVAB5+FpknepOQPOQHZcM09iC8+QB9UwEm4
Um+ivSHXc5SkpY1O4utLMXfkKJUp9pWyBmnrv78jigNc8CEFeFWzO+//gLk9fgzi7ybu4Gnq7XJ+
T688OblVBYITat50WOIx7jur0ZTrQ0tFPTN+Uyl16NuYHje2C0q1SknHCcZwpcR1wWraOlCB2IX6
Jr9MqJ/vMEF3y3svX9bRE0T0Co37Cgf7WFqaeAZwDZbsiQr8fRiBOPaqHp7hjZkCb4C2aBe7Vqcp
Z4O5stjl2k/y4JTyWnj41D50IqXTduKprpMmx2RcD1SezBBCtH5jd6boX4exiwE0c/4Nw6oo7eb2
MV4Ybp94KFfWnXPY96uP7ucvgBJUxiC9gPzltReJwttLCyOYVM7zzBYQN1oRuit10qZXvYZWD+Y3
VYVBYme+xqQr0YmSVN9URAoGpJ5cwlegwv9VKozfyQugxP5waH80BKto96Or5ABJEayXzFSOiaW+
TbF9CRPSpUJ7foXZOGqAk2eilk9EVJfQ/S6GOOSSZq6XdFfMeTgLG1MO4G+HgJL7t+fPhUtm9cno
MVmy3RMKLNhovZwReoxWtw9XCEO2xEGo8l5PiQWkHa1TxtB7me9slHg0/ei7PYD892/2Sd4/Yixy
eDpkAFUjdTilJyaLmGL6Ts+ejqBte6FEDz8LJSuDpW9RSSVCsOPJS/0nYmZl5S1E9B/RZP409PWA
kfkCKgIfmYNsRyfB8l5/WYLIidPbN8qxjYTw5DRSN+CEJRtcLgKPmOVcGbq4Dadj+Em28cNb9+qB
JiWdwziNWn6W8cs8ljCeT6Zb8anjnpKKDNxJ061WEJPbQPj4sVRHDJ0apkO3lqAKP0luMIomjCnr
vTH9FVX/6ls8ldBr9kqwvrLm5GXCYbeoPN+TfJWN7wjoJEjmn5MUxh/T34XHu+X45FXHt+HcwSLd
hlkZDo+zi8JeL7T8fIiBc39BgNLoh1ZCNTcv4CJlcCC5YhZ54JrVmM9+1w0ggSGs2WglXmNWNdWI
njDlWTifRVmc3t3QqewB+tBzH6o20xdC1zct1zt6myhVjICkA71nwXyhjrqHUF1G7lchpBgCc4Hd
CDiaNPXaaLEWGhlgzFa0FFkFsbmKvZQ1cVjl2dDKfB5pwKfndbWR4X7k0ApHA4LuhexCF6tHb97z
lMmGYwJm9uNpyLyf1sbEK0XpBS7/d4tUSh1eDoJ5rqHYcfDffHgDzMAWj+zK1a7kMqbs4CcO67uo
HVL3qkazt/BxRymJQXOl3tqLsD72C7ExFdhHWpDYEdNfVgDxY6jdJ2xZ3jcM3mQ1mHZgyTVi5EF5
fVsiLQAgqfxWsvaNJBBdUSdj99qrp/g5gjkECYFEsbKcrKeK+JiGx6NzyT2KwSt6YQpSphAQ2xVD
5XOupPaVvTxuMkP0Oy8raBL+XEkK4bK2tiq+WJCAVHhElexLP+bz32SHTM8Kzg3wvk8q6PCTV6g0
+JgbB1KexQQ82A4UXJ5fxpNeSU5US0yu4Jw/KKww+RyRNuGLQB37WoJqE+XSURzWdis+c538/Xar
JuCeKKLWO9Zh5miXvYeZg1Y8ruzdJd5x6LnPyJk4+byzoFZxFeOgGlJm7LPr40D5SkcEU1QxGGds
g7bcF5Qs7XYp+zDlWkkt/+hf+tnBtFuXEekNkIVmZfV/l6YJPrb7C8LUnOCoBKD/KjbNCQ+h/08d
xGzycQIHUW2BocaaWsVPqtWEMtQja3ncO/RqKv6UiAqDVqHnGyCNpuEXmV1plThRmugqAbr/7H+T
6errywrR5ZpROJ1J+mgLn6Yb2+cQ3Fegs5pj5QaEjeNyf9P6EJCxZFtyCbBhm2SifvvHGChTntSG
lZIomyMLaERxPC1yyi9rEQrrP1y4TcCXERzSNMrTAbUmgLkdYCMakKnWeS24EPkvg5W0zBHaHJ8+
Gc03LjKxcaAesDPy5XohnI0z3O9QB1WvjwwcXWbpK2ODGCGIIaCVhEwfs+8UM+7MjdWPtEXdrPLo
9/e+3oPROZiGnLkyXMc6IUePYvHcrvHI69SSfadqhMlVzK0wkrATEvHGspP2z8XHVTntcVw8fZhU
ncwLKzxm8CP/eyuzYzu9WQ52nXdGVzlqmGkkls4/FAh3leZvZeXVeUQIlKWVoRdZsyEVftMD6gX1
ljSqQWud61b1tyZvVEjcwttla3mmPYeJx6Xdos2K9XKRdOoxkXRfh0ogl4wlgmVYUEPr/9+yyM4c
Qh/vf7hMGFTaQNPRxHK1r6oBFWTjjWTuw7/Zt93BtqhRFPNO3ZHkaOu9NcarJ9ZxgI2QGtdSxxt4
Ud5dizcdav7Qb9Tq5rJXUJo76s4q9Im1Eb5PMeQgx7XAsEC5xRQj+oheYrgw0Bm8STPhhVSZ5ov6
tgRvWHBDamhoyAe3o1G250Idgb3owxoCeXDssTIsrWzGNKqQTwA0C1o1vRet8o1j71pFJOdFnxrM
xn8xawXhfcyFzqO3kVmEEm5NLvoGySL0EFepwIFXLdpg0xxIQbaKQbzXXdz5/VIRqusadWTLkUBA
fo+8zaZTWnS8Q03Ab5V6eGEwbgNrbG33zWL/Hbn4Z6U6qZ/852mFLTmACyXSj0gj5TujkYZoNJlc
dqpZPZ5vR8fzcou2YkRC40tg3/XzmgYDWzCOirzi5jjQR9E3O1qG7ZCGeKtN4RWvgSxhphPLQDwE
Xo0Fg/UZu5SXrRm8r9kxNY14Hqp3Rk0S/Y5Ylc2/KoC65yCFqMBwRpbHhcrsHnmkJOhy/uZVOcZp
MnidauiQiNTw/ueRio3C6GX6S0fyVfoxD+CJtNPcC56dapVIUG/5yUGShpdXElMYptk8G0iJxNFb
ao5Mw1/vDj4LRu+tOSSs/bY1GYFYBgpqKKRfkhoPvwWXHQuG0nUGCIgzvJBR135bQlk6DN+ujBvO
u50M4kHZ7VB5Lox8Wowu1OYi07u3C0LBnrMTGI41Ro1D6F4bXk/yrVU6EHmF6oJ5VElyU3y9U1id
WbgE79ObmQtzo+52H2Bb7XRx/LIZvqRAfGHRoVVXhdz569094+Nc2nvkqQJzpVmDALcIhkY2cQ28
taVaYz16QfYM9dn+SUxaK5YbzRim/qwIjsTLETJqcoAckrVZ/TbhGhOR0Bl2gtQGY22LR35vSHm8
wyzTZy6iPqwI9ksCPg26+HxV+9OSw8MyxXK3I2Tphdg8yfzOVdDN0HqugSO8RHbuWsqY0J8zVUsa
F8w5Xmp/YKJX9y6cVXJD6lTPtbO9+z4Uwv+RsMtu3jIGLc/ikMeS1o62UA4R4bJ2HsQAvuac3IRx
VpnR7UlRs1J+ZULtUoyI4z/PnjuDFlly8AxCrQtg3LcPgrvEkrTwLKlKdI32SZpylLjVTybtbqCt
AhwDDIMgNDQ6OHZ3q27GGrBWnXYqHI7KGH5QCmA584HZarvJ6CP0b2xDoN+7hmD+2EYhsnfRc49s
E5dMnzlcFiVQ98+0j/0Yr080aIlNRtdIt4LZHo5K9QeNdoOIpIIQUISA75VbItY+onVyfqtFHyGI
hi7fMS/hLHybNNdITSCXgkKi3nD+MgJvkz3Y3On98+783oMYsXgCkbpAriuQxmyF3IJ0JFfugrj9
kjhKfyzff3VkpI6d/vHjImv8Eavd9Fwmh7qeCm1YV5pqe2ZNT2OR/g04vLuzHiH6YVQskqxASHvx
EuGl+sYRrzxcOr78I4kzt/uSIIjB6q7jD++LuXhYScgo6dC/zONNi9MXsnxLKekZvVBioLzS3U7A
1lyz42joSQEx3eiBPxeGIbJrm3lVErwkxxzPXU2NJdX95grOP/5niDe/ZN/ajPN5lJg5X6M4qia3
Paw+H9+sbw3IZvoBYJ8Sefj+UVcP5GsDMIZgveXax+Q77n9UNz4uotpzspJR3BTn981v8S/qes5w
Rk80WpGhuBobHzL7NsSTJbg29PfqYsTHRGH86PR8eRX5z5EXJlFnQ7AS7Ah3RT/jnHvjfj2iF9Q+
pJCJbIKcy1NRfKMdL3vBj/4TU2vDKrDFMoTR3vn0RzuYt3BQm8zN7xt0XpqRKegOV2oIy6qHbSWx
8HfdtGhkb3F9GVVAreeSpxp0iYZ8kH6HTBD2n3awYyusDlL4iIfko1pbntaVj9LCoTTBqv/mIgQ2
A6j8u7+imOG24mm9VvQVH+j0VdXPZKnDBf4/eLoz9IZjsNnuyjaofvBB8Mfwi28stBI8GvhzsfEg
hlRNgcdFNHJ0+uBm4eXlznb9j7w/FrmrfklffOo1k/sNwYd5Z7cqs2No3ISZr7h6s4WFBvCHcHBI
xxKbh44brnSSF8Li3n9yhHtovjg/zvTVbCaRoxVyhyDyhj6KKyypuacZs/r6PmobxyvV5aTCCNof
fGNRR6HhsOr6ChKiHlLN8JBJBOS0SArcIP73jHKIOrsscj/t/RNn1eD31d8TpOa1Jd+g61OdMpU2
tjAyEk5dfdauFPhNQOQBBv+7r00w5s/5e5w6WqQyOUVmFNRmd9eMk6+uBOABMl2iuLtUYIaAtVG3
4GGdg2GTUprRhCbwmQK5pWirXjD+ZNjJXXWanciRND6bacQoySd0UoywiXVpkS1rkyfvVF90KmYy
p0URbCT8LTRtP0GmqsrA8TSAbhqpsGFqYdWUR/kw4nM+8FN2a//9z2+KPlT/QQt2ICHlQUaJDMoo
4/xr7RNIzovfs8mcyTQFuLfpoYDg+GqO8OerknpHBKye6IkWFijfIzzmqIVezpE9VLaLVXRj/01K
Z1ShqXu2+Ow2rPsG2ZZY+ItNLPUMZAH2U9ylSOnR0TB2sHZSGs2v2q8kMVmVNbLAm4vWGBZIysK2
/uNBlttTikFqGusja6bJM+hKxSby6m8KejgeoM06CASk3ZsxYY+OV3/Wk0pcDIlnjZCskK/hoPKs
Ms2WrA9xw4qpqAwH8MraUR+32K+aEoIUEAumhmUpN1zLdwaSVsNEuA73xO3pWCDLfItQu+bptwQ+
Y4cSu40q3dJiRWDzUY/a/90pgydFmlGEYLE5wNRqm8Psm1i1ZoWrgGY3gEQ3n60bw3krksoSoykx
ymxn+ZhsgSwmoBIZ7AY8vnxjJO//oLrNUnnGxS5gbdFleH5tn4K/NsEKNhdMBqvS02StfVxAvOWi
RXbm+G4+RXPymJL+q3RjLQAt1y7nWSkORJDWx/Ng9KvHa9ze/+wdr6kckBhCDqCcVRw27+Tyw7Hu
fVstHYemOzquPbRWeyGvud4qpQV93lW7fd1MCZbD+mITPMob8aJWuJ75w6l3mgu2WfvaBwFYbG1G
4Yjid/I3zKqRCc9mKrW5YPKvo9JUJnsc3PgK1IVGHgOR57xibmcbLGQlGQo5wEnrts7lijXDrnHi
NZXtcQ88RT6q5pfHsqP+gi01TlNdIW/PNoTOxqvDxDM1izPovPXC5pUVC8cWMyWIbwMxmIsvm9kX
WakqjAqynxwNtuasVvL1PjimbA6+GLDHhX+eVPdmgTg1nrHH7Oh6oFcVysdwFpZShoTW31AbMXfx
f7KQqr8WYelr4MP5XHXC7cgYwPuFxZgNYftcAC4drXkriHr0CrJskfKaWdigVxAYf+8K692CQ4uf
hbiJLMmoY8tf/vV3HCD3txqBAiWoSbG4DGFxEmADz97TKgkWcU3BEvy06xknaQR0EOCIF8hwN4r/
70N+1kkuwHGWRjREu+WQU2WU69Gw5IZVApC0995tJKLl6SUPaSgTUgE3NuJdzriDH2aDpHcQnbDV
S6kSUyIFRK3yc6cac9j0fSVrKG2oYPHed9ZYbaYWpY9CiDkOS4mxTG0ZwCkLPhpnRwOIvASVZPEH
ShTHxzptnCVN5pKS4Jkbna5vOoDhdIF+oyI3iYvfFE8YDWMPEOQDaEEFU9jBqk99bHnrJBDBYwNJ
9FBRhgc//H4CEdDjghj0tzeWlDZVqbuQ/39iTGTckkeytWchE6ppdZdzxVCk5VFbGVjuExrCxx/u
ieLNK8dLOV3BJt41BGXrpuS3W4AUklUDavQuio2t332s+TD3imq+d4y2TbI3baAU8TNKLQ+pyuL8
8inIejnJZOaRSQfbdQdxc07KEH+YsX108FO1tJv5OnwN+tkkPr1Cq6JRHH3GIH5Ta2wcfJ6Dk9hQ
sN/SHE3xyrOqjqSMV/ovaYbYxNcH8KPGRouu0/3GJ7QSYT90iytSrXmS8uCLTsZ5J5IIwizJ00kI
zU6rq2FZSfrdURLvQJuZvH793s8xL0M5CkXVFpnuN/dif71D43ZHTlx5NHe44cJx7cK1IquYET1m
aYOz3ImndRHgv4DDSPMW2cP2kRu3l48z/Cv/HbtInsbleWZ7IJN2xjaVj6v0SKBQN7QGrZNS3hYz
KG0tNodAypgG3GCmkgJfHIXJVG85BAe4fwu9gU4/un1MrtJFTRZJwIk4s423Bi5Gbad6Zc+xmarq
WZ7sNp9OyYEau4h7u6FQ4NCH8rEBQMGeivaGDj/DiNMHu0q9MwkSrUdiwXSwGivmL7vI4N/PSMOB
dsjsrclZN5naQwbNl/CHRU9Ze2yXErg/s6tHhZ8XVtTPysVv4EuO6l8lgBaA5D5nzfpihIdtcY9j
eQ1vodvqj9LFDjAK/oRh8+WpXXkwhQyczLD/gH904X31yE9V/80CteyfXP/urtK8A6x+YcqkvCDz
1Xe6zMT3TYyn5S8/NhKIMeJvqKkaibwk9xWXUXhA6Mcboo/ezNI+nouLgS3refrcS9Sf6QM+hh6H
8snroCsPVwixgJAq538iCNtckGPdOv/H5hsoh8ALmBZU06iivydiOvxw0r7hHOp+6abFpLO8g7V4
9Pj4w2N9wb0aHI2AaT0x/RLiNx3ziEpXTZ8tCVe1+UJ8yhOOEBMO6hwqh1tYidbAdG84OlFdrfx6
3/8eG3G1vPumNpa6/7xCeileXlkBSPyH6MhTMvk/1IDZdd3a+MlsBUq6EcCfxZHmx+CvYLrwgGJ5
0fQKipINwXJQG/GLH+MV6TNJ5gkMd0PKBDpTijWI7H6XCqabb33lDNJvIYQVXl1QmIKgecvct3LX
PEkAWafLQXF8gzw1jy3ps5bFQpSHSwv/lvWYsUgO0h/5emDQqF67t9mLD1UF7t1gr3EefWEmYxSq
Gp7zC0UeSblGB7hlgL8A16wQJcxju2QXWfdLwbOdJStviv4CnBL+EKGvbmS4yHw31dJuqYwCDsr7
eL8J2fkrOy+Ng/o83N4XU+fYKgRtCwZ0NGop9EYPjH0CYOfi9x/0UFgpbyOL3QQa3gL1COBMQyGU
uVr1m2JXECNWfvV/9ogY0gM4yc7wd51o2E7oU2dwfSqDneEdC/yg4N0zzwk3H09hHUr/MWgBiRkS
XBXKFkclkyg3z5YWJpkO1RgwyoPR3DocqfgVNIl+wSmA+nmHl1gDHfXLkCpHGWgxJyuH3jO4gqVr
SHTTpMJ1MOe6xKX3NHmfUya9VcJygcQMusx7pEcETWj6mM6oREvZ3P46uBl5+P0HNiG56phB8Sco
u2Pv2IzvTlYin15WU/9Fpp3OSPMbazTIR2m2Cm/JFsOHMKIGiZJ0wOUu/TNLmWu+kMSpmn3Sxsei
xwnVDByoKB/YOiU6dGY2nPH9w1BtGhTV9YtgZbz8GZ3LZozwKgXQua5l+cTQLA4a8ZDhXx0HpNZl
Jqm6KZDKBxCIF39sdU9WtuYd+3+zBH4UCJpg4Er9k4RRO0t6B/6rGnSNBqWbPjZQpfcqYNWr0KpB
ep6ka1wJDFfpfjMvSoefHU4vKm0xVnbsXxL/9TlBv2reJPW1e0zEKS9G8sCrG5rkkb9P8G8s0qlv
4TnLyvZf5aTw6HlEGFkSSjgMjKGLNL/WwQwbMVtn2rMZby7kuG6ztNDO0b1LeP9RfepOLAZ7wS3X
mzHxCKAgh0px7G57UAXFi/oK4L5JWom8UgKhe3pk48BryMd3lwURibh+U+guCAxJXDhekFNXeNeD
hKo0+MIZgrlbBQaGQ9oHcESyNTMRVaKvg9s56Fn5Y6b7/gYN+h2epfeGfhRW/L4DKgjHZuHKeJ+S
MTTx9ygP1pAlIDNWqfbf/igvVgxgt3tc9sLVisE+Lje3gsm2nLcmk9Uzjp3BOB/608t4BFuvvu3U
Hdb7IqB2C5NBzB/U1GciPChL5hCVLu8ZtgZBH72MhFReMy14BzHL1hXfdvVqZtWaT6hE3+tWHDDX
HiJl8F8jK/P2/ehy5m9py6F7lLRlmYaFNa2+MbEItiNTCruGtfupKM6/csju2B/VoAYORzCc2TVF
+2+S2lwr4ow6lsF8qu7NOXvgZru/BVQSOX1u3Q0BqQpd70hpPBZ9wF98Ic1vypC16bSg3Vx8LriJ
PAqzw03NIigHOVw/mIFYix4uyzPezWoXCoFkBvJwS1k/Omt/OIhaU2CnFNl3A3NiVlxkXYKOIMS5
/9kRN79ptNCgufS/ekNemXOaYWCtnxw1/4b8V4dMyYAR/prmyuEdtNdgxMfQr0c5Lj2wijSFilek
Pe1CPBHsTlrr9F1Q/Sw0+eEVAZpXuT+jeCB3hnNu9+lZEQ9XOix+O+33VCzaLebXCgYwNhSCKuEq
PEiEdPqhFeo4cjB3khqKZvbqRRj5tVPptZyRJFP+YQbnZawg7tnyXPQdPtys5E/PtWJK+BIwfriu
vTF61FKQpWWJ3JvlPEwy1rPB5sPbOEThZVIPVh12MliOuRbJtBnh+QTrdoLMGXRDTbtdsB/9auvE
48e4kDOi6hG3hqgbnUXnD7cS0angNd7F7PoJm1NCEv1TQZZ2/M5bPavhFKX48hd3lGbo8pFeyl4v
b2GINR7pb/ZYwx4GzY+jFvsa2moI2IXo0kJYieXmRQXJVmDsm5i24Pf04dVgwYtA8kzDqVpP1Ey6
4amyCJw4BLQSVllBLCEllbPQvD5Bgi3un1zj+e2PVZ/Xr331zwXFG5MHTX9/oeyG5F/j2el0uHgM
xB8mW6CafKrTj9S0xDCJaezoS5Phabx7BUQr1YimTYAeEhHyfyOrxbK5qMBuwT221OV5ZidVw8pi
ogBEXvuc4wAgzoWW4xE9OYG+ytxOQx5/LwOuroBujXL3Yqnyv3ny9++Cv6c2HWNV/DlG3umVZTJK
xAK86X+5C5Oe9s2RamdeO6kUy/i98GOGibG3g8Chxzi8MiDLEMigkSr0D9uRZYv2uggtcJQuerrO
pAUkQxsAYxJlVbfban8I5vr68U922j9ny14Aq2peLjmUFHi3VMxDerkNWDEgjB/jWdwpmbMsAFj8
Pi9nxCI9FmcCwX6G/Hnp85dCskpO2FcPv3v5K/yx51Oq+QIPHQBQNrYrlkg5wjSivSPViWe31xUu
UAXBCRwLLVt1DVEdAspfEGeuLIr39q8DtTuD4kaT4+AR2TWz6gwBpzX76Jz6Dxn1zHypDQ21Y+Lt
e7P2eV6AiioVwypqCn1xWb2MjWd/UfbsPgIGIBJR60uez0zsCqcCHBkw8PvSTIgrrdSeEneX7aWX
DQn96f73yQouuKmCP8W4kanEoytcAyHpuPffkHNg+rOeoxRi0AmxLHUxHvRhvRCIi2nzNV0nAieC
XEE5yqHZFJN+RpOwFljYYGXVxRHp9JFktmw/8kONsKTvTUC/6bdJaAz3FrwsATrDKq1bsAuPLXwW
qbyvQTYcxhJ+qjO7HK1Rs43UtqSiI8JbNg3KgqU249aj+VkdFlfs5VMIj5EZQ+mubWjIJs5GslV5
/dQwOj9xBUMGv4dpKOmlfQfSEBTGBBIc00Ste2jI2HCgApF3syz8cDq4/4kI1fA/UpwJ+Wh0cFvS
PLXxxBxyBNqH9i9EGv3kODfQLiAHf7aiUct60hizRQ6GLT4FfmNIPoOkv+Ru1OrB3qhLR13yVTS/
Btf2tF9x97NNHQUiNdB7IRuEyio3SXtAcBD0cj/1IRrTewQ4V2PchyaJ1Yfn5ImatIuG5MfzvIK7
v8vRd+giP12KAR9yGaGKQlVRjVfkPsJbCnqHZpve/wj1L7BjDCvUUWzoVQlNHECpG+j2bj/ceNlS
eG7Z0OtASFJllGZwQP1Al8tQamRmo+wa+JrSLRDi5IqmDygksSc4ijSZNIBBzzTgyEDL2w2L0hQL
nbLUEav0ZEgmyu71ip2AIzFGdb15cO7JZeJDzTsPnIjSl4b5uLjIezOXMHsYn1tlFaRiDuPctUci
FzKXnFDjmIMqU37VZvq1/8ibIsU/Rk/6S/vNnMkWGapgqx4Q+4c8Jw57g1p38Xkig7PYO08/2NJt
T1/Va1aWgzhYcyQf12MilxSe+/iohv+qXwQZGcxoxWJKr3UwlTXEqa/YkqiA+qbt4cnWskSrKjbV
QTXzdGTojyDXD1F4GvYHxsCVYHInrgODyHHfYsueIbcotX/82q/M27Dp1SZLQQBx5l1SAA8j+Ez8
SC2ORi7eUU30XN0xRCXGcUuvR5WM5930jvUbPvB7R1LvP80ac+49s4w8e18l9BcsFG/gHmeEI8lb
l49pYpgAMTa1S1Cd3VEymmmBqzcOuZo9ozhtufh9yS0vSyqA2EMX4npvsqOLdS9f5dqytg1jM9LH
zIyVbtaplhPFwziN3QzLoHrLjVjyvwrYcAywhxwbaQ9P3Gbz/B9jL6Cj2kEfFFOymbZJx1IEAWBn
B7ADXO3KdLLqhr59BpJpplN+YiNBLiNyuFB1e/Ki2aAZDkDfjob6ywemgTc4M7MegsIkNxs6NTwv
9SpKIJ/CqgG5vxplxfXZia/pUzLdrJX5+BT5cY5CHZvvKzxnLXcjS1O35mVUiO0Wk2hjgTnUkd/+
5tnjQWKMTD2iiKj41c9rTxhIjW+sTNvImqr74E6tbCKD/I8zZ0hXdDiSyzuaUa9TSP1ujpxWfa3R
pZ/MiruH74tG8/HJqAvvDRg35IMYt8lss85v2obcDJyXMwQ6iGPckVwS3IH03qWNmTortJlxYHXJ
K27ayqrh/ifkEIHPshg6gIB2SqwHKfKnGthRjqWI4P5NSCnpFALpE8aTqfSJVvvYW34PDo5VABD5
s0f5iK543ENgU20prjiG15bCO2dlrhuXUiEcTUJLMSL+xjVNH/gF4Civ45KvO7kseUGr+fYhjLIF
G9vXFcOzXLrHmZiKcbkSkMLrMbA/RVC7qvU05aMG8xQ7aS+kNZgIh49bZJpxc8fQ/jjdZx/ZOoHh
r2hha4vyGvQLkKN0c47YqmExzLUeKf3dCxZZ0zModS8TARE82+GTDdUovDGQOwzKJzWmm6AbrMFZ
4jRu2PusfQUScDAWeetQp7Ax6gyQf82xIsh8aknXTmPHjOuPjaYpvZY7NA4Q9Wlip3IwEysdNF4c
uPFsVT3OUGQYNXH4eylJaDFy9uYgawctF+y1PhcCUYIxl93JN9xf9vkK4axBCzh0Dw06ZrN1VNv0
eFi9Bvp5sRMpI2DdSmdY1BUNEw/f2FWFDPMLG6uY+NVos5fSgChc0g/q86tpE4V/LnuRUht2tQiC
RzoIJwrJwqucyEwAAwsjcH2aAgLLCyfg+YokfPqPATD2B42UuG+Qk2XAV5HDBivtgpK6PB7chSfp
X0lMkPQDYnC8mqQA/jYY1byTRf3yo/moLWZUh/7y4o97rK2o576PEtAjir5+editkFEpVSNtDWIM
/2yM7KwQrNtzIy3p71/FfPNIwJU7v6vNytTf5/gke0B9d1TfDTtHZExeMHTAf3wayuIErZU616aE
M7yQnYp74SGAu3mvR08s+K7DisdJipNpp0I6FcnlclXlqc6hNQnaGv684fvplG+YQvqfAF80NrNH
oczr0ql1NDDEPAag3MoW7rAk7ddoxT3pUflUxP3wckyISu22u8yLGbRo4dH/zR8aj/1jMFKfvKrn
sUiaFmVINNTrbCVv0Tf2e6DK3NpkpIpuhxtIejxv9vU3ztArA4VdQukQBxH51lUFFanbMK6DeZc9
mHbUoi87iqo6NngcNCaHt7slMovK9JMJia1I/V4wYU172xierpu8JEVMW3bVj9TOBHU0NzokMPVn
SBiUQaBb5ChXq7SRb2dYFYxjXa5ysdaNkOxGJq0mPYN9KWoNAOmiV3QAK/vhXvpkerK+LPW4NdMC
+ov14wdzZwRjD/oMnQtsp99mF4OHvfYg/xR1VHswOijfZMr4Ur7TBnCyREGhkeh6HYG5mCiN3B2I
nEvq9pjBNT0TiISgRlId9LovjawEs0ltFL1J4H5Lk+L03zHcjy8ya8Xl/H/YwOasyjtGHta5rlVt
O/Xt9cZdUEX8UFkFSpaPI51n0x04RwR8Z/sybccauVLhplrKpJWWTQWiNaDzTb1OfVJ/dEI78Di6
rAhAgGM2mXmCAHgYsoOVCDrq//ma0C5Rrz3fx68CabyyJ3rCnT7c/SiMoN5UFkWM5z67lf542hUt
3Sw+2s+tGfvAeZwtmbEnxnDccFU8ZtTr2Q288h+gHT7ONBQ61RjwbzifYmnWRFzYxfN8T2ZkwW1c
Npp98v9Hu+JGuamI0QwQTmXtFwE4bJYsAyhucSQGthT02rbRJETkVA28Sq+irSvorxjQw8/PBxTS
psy7rLvzsqT2gOZj0lwxDC/r1AisL2bkuECInewYwmEmGzxy1Bt5FjQWU85ty6Ds2g909tfOArBz
hBpE8KBsz0bHlB7gVymLIFNiJkg1eMeefybWRr+JHEaYEbjB/4M1JKBcmXIGrWdyVsPj0lNZeb/+
9sv4FzHFIzM5X15Szn7x771yWkjtk+1C9QhCfQDs5J8+vEDuNEf05RORjMKGzsblnWsWGYHJCaQV
X2v76fl21FiGpQNPxKRkaotga8F1FqQ29xTQs9L57p9NvmajRL5GTiaQv8HwZ0fwtCfdYL+1600T
hcSABhJoi/0Lic9TJ2pAKSFQCa8LXHieh8aU3HNYKXmKHexQMQ5ki90O5xwFIBeYSMQI7ePcOWom
WDEGmB0gZD5DcBxqg6ybTZ6QWl5jWm/CPvacrGolBy2mDc7oLcJh+yLU1w7G/U/NGRBx2rdNomy4
iM/e8L7kEzCnWkdBRXlOs8iPevL7APOJDsA/Hu0/qsp/BkGOiCG3hnp8xbZKJXOcGiyXv5AH3q41
PIUDDlcTCDi+IGIrsiSGvPQzLiEdRfgOIOf1jThpMy7c10W3A/bVGWIRaCBMMTAganroDC3xEyFy
0zYvH0RpinIIm2GKcc/JZ+3oFeHBkJyaSv6ITkz8Hmx6JfyM6IQHcgp6+71YsWZxD7R/SmX1HOvJ
UdabvfKRnlRu9Ze6Ru75/GCejOeeCaRKXXeTiIOe2FXfX90Ax5wVSVF2NrB9GJ5Rh1tUu3TJJdEn
CxFPwMAByg9c8JiMMwad2s0B13+xJZMI/UaU2K+Wm9o0Ju7AFASgmmfaVs1xhiDYj/cXHbAs2B+g
L5WrdnOFCPx2kYccnFbvtTdJflakYTDXcTgm+qqqenm0ZlXBbEorpJ2SKmZh28SCptKpuS4vcbA8
ZvCY7lbDbRSEXBpLFANdSEd+9UzOYDngd1NeVUyOxcf5a1jzwdJ9nCHp53C93CQyOGvpzxulRGaL
sK38nVisQNNkGnag3Chc5vkeTcfV1Qo8tEEYL+PLGxNUJVvUoLAXbzrr1ohD9GjxEgnCvB9YstQM
l+bPCtXdrIsInrIFKb/GgRnXmLHpcPqC30dDIwaD0JdQ4u3u8JqeVbERaGVDtZVbIy55iVOVpUEz
F6NSe0m9fZPbO2eVdqnAcX27wVv83JXDfZQ8driimCEIP/QxW3xJGmYGGDCiSclHXybThaNKlACd
yt2iJVb3SmPiNoV2qMQGSSYKSm250jLrSxPs06ZRBrU0DRN/yIZB7OYCYgdg3oKN+V/8ckRoMutq
Jg88RaU/ouvKIkfSrHwBSRqRQ85mLqZ+IqVv2Ee9hHpToYistrbAmnLztYhruo/VL71cU/tZwl9v
6fBFqqzdJWQFIOzD/zTBfq84kp61p4PkZVNQo2IqnWIU5nZSZSNNfw83wdJiXIuY1zBD8TZvOeHJ
M6Kr7OagMgJBs3F/ED9GC2lbQKNnFUIVON+8R4/zUpr23aSEm+8OHmTT7YFU5NfzH5uGS4HJy/1g
S0ZKmDfKhxEhYqE04N3nv8ELVupLi47N3vsYQ/oRB03OFyGB5BHk27SpIV61bdHQKsNHTOMgbB3e
QXgYqAivmooZckfA1x6EefNRKDp1/C3mO7VYh5l0KGFoWACFD/YSOLRGscsXKqVpiprFEtvGuPvd
5t+dD1fSMeg951A3T4TSe6ODipybgFQsQM4EzFe3FQJowElQQB155P6Iwx8glDHNjOWhN2vcC7vj
VX+UY93fPShN05TuguU/AO2ZjUsAlKRs2ux+XMTvyTMqBJbx2iMiAcx+XGjddlPvuy2ppeQEZ8KK
Yn8zxsyrbXRdD++0yXmu4UmTVc7BKYfhmGP/9LE9p1c+1iAR/Ryj3UlgO+moYr3aBCkSbxicyIya
nMaGuN0ZHx2/L96F3sx3IjzY648hAmeQ5enXh46agDgaRTp58tMlqpxruFDPeloQmx6T4Kgyp9Y7
6p19KaEqg8zpZAnxPtdYuoZVk+ca+nkJZIT9FcAX3RfBU4JpzYSQu2s4XAGaG/HmVyMvCyasSz5L
ssT/TUcU4Z8gv7PciDXvMBC5QQ1ugWZOvfgUQZrwradjoEQLqO2SiZVMqPLXlBoSrgx/myoMCAUY
2KEzH8633K/wkKxudjjeWPZyW/XbHxFcKzAgp8ExKXLLyu8W2VbPzOin/kslZS35srVK5cNJZXgC
8y7ooyyA0OR4EA9n897ZVYBZ8iJXoXEiDk3D2vRyHlwhCOZEx45ixgWtVlELuPLoIdcpxsiYZiue
46Y8fvi3YV0syGaEdRTYO+rjTGGMJug8lnMqCkIZOYfwyhnh7tUmf+lxotzDllSDxAbuX6LHiGtE
1N0zsBENIqGx9EhjVL+dI6tXmtkUAxiKEsvzuVgbZMkK3V3A0PWb6bnx51IH++I4Rw33AO+6129x
3NQbR7bLeZ3zFcX1GVDAD0hFdjdGrxXI3bVx8lk61p6PwIuDW1H2Er/fW+jsPvia9NIlqvBvAX+e
JtW18OdQsLkvBp61diBpnPafan+4U+XcyTHOQe+EJV35slGT628BbDE5s97C82u8sP4DIUxX9N2Y
ruflFCsQZ4Uz42M+lj1w06O3jHuAyb4BQZQ1o8in3JhoEpCaBk1+EVCbtiCdnzcs9N5Nc7crwBa/
oA15x4CpEUXvHJI6bFSkSoIUpxTZleZsdEqq6W9i/2Jef2b+GEs2chlDcrWPEctgdLvkgS601QIh
yBh41lsaVDIr2TZg2HjtvA0KErtMtQRhYnQWPVhs2fVdyi9oGXChrhPLJC4UIri7IgG39gG9qYBe
VkddHqvE0JtqPk/drmWyP4gAfTRJThB14S9WNejTluRjOVXSes6OsKInx+9QIJbiH3ko5crT9kP1
QIGVgmHj04314aak33MkgW9DjpMwBcV8kvJQNMZo+jxeBdh1NwRvfHND88zH0xk6aWinAXUk84FS
zMk2ekm3jyOCvf1G4BlGrv2KoNk7p+xMWGFl4nI+Rv6M+e6rorl0lx11hmKGgLQzcUB2OPCWa6tS
sJrM/gvcDs2t3/1ZPZdtzJzPe894WQxTSOIOyWJ31RTWeJ+ueiV8sY3P5AYW2X2dx3Jv7TZnyRNA
3eyeBqwyTCm4tL7kFTVOeozw/c6+SFr6999WkRzYOQNPX6XBrdGVz1/AXVXtKe3T0qWmDNunP3kh
OWu3Yv91J3eFRJ7pCMhN8IqsP/E816UZFac8CsJ/wO/3u4nNienOe97mKmzyty6ziZd7MU9/fp6W
HBc7Y8TbwUILzHSWIJay+YAI+UHxqaVpNu8AbS9rYb+ETJ9gq1ukr9OtASV+4i32ZRtn62lZ8xlq
HUPM5S9K3Sc72fevUzt2g/BpK4631M41uMcLPapjSgExQgVUl8wfdvkYsYj+LC+cgaZ/th87gAL3
oEuv5hKT2ViZh1UkqThX/xDQhXRJEaV4qc0SKuZDVhIqiiw3cmRHxrmlytDxuAZRops7QmWq6E91
DUFDO7BPyfvlqIA8SuRvyJzob71libsNQeFUCm2Ow2e1p4sGt4gBej2MLcK7w1HRBNa8RJY9LVnq
3W0Nd+vz0df6wwykzjUmuaNfuEt/CqdWJTOBrQ0eCTJS2Z7IQ7H0WQ1pyVJ5MMGBbLobriBmSvvR
jCdWqN16qG6kGdcmFCn1QX0k7e8mhnvP9a8MuuIIWyyKBv8UfUntdxnu3nftk+/kSLBMQ9uYNKW4
NsLba82kSHkTU+LWWEARpPGjXiEvT0l7qlmLNUfzkqZPnDeZvKR0W4GDNecJdGzMPkhN0dIcTGd+
c5QZRrto6ExGEIY/0qibKosA8paSlry9EZobhMXXyzovPvvPS9QtG4tzcnBLkdqygExOkmm/UkQr
kQUnetGMJQBPTZOpZDZfikywJuU5d97A1GW4FTw9r/p2K8dtHwT36e0cKc7nO5B25++n1pz2FiSP
jMyNtNx5c8wx4Urf3NPAWoNhR7eaIKhdDUvcVRmVSyk8fWx/OUfUtlRO3Udx8/qnPWWEZBZ3okfo
3VzApkopx3xjnVKhQrYlzuTg3HV2oGiG52De3YE78B+mSOWw8tHxQ6f3bX7ZGgXzhgv93up8PC+c
zJxLTDOs1fvUXHF8I02XotjcUJJULpVodIJak1jOulkt1MIB0SaitfYNAUcIiPX5cCGiTx1w3x82
9EiNQVDFpXbwAybfuszbkwYr865CXCsjDeDWVei7OZ9u5ENGYfxJp7WqLBSInQRCudrEC+wPWoWu
aQUc3PsHNwp8GWBv38DCjC9zKnFA4TbQdfoTvO/aD9//u/AUrzTCFam/Oc0p1fwv/ZhRaoZgdDo8
Abx5gi+k0h52ZsjSe6TlqxM16LUxq5pX9C0mVTSyDdK15ptQ6DBOUPzMZ50+qlX7jUAXjETyqKMI
3DAbESOCg3BAMXlqF2dUyO5svimNu3QShItZEWNmAWlsXsBQj0nxnVPKRt+4lfoMw1WC9n34UeZR
u5as+tSunvbSfYy3u3AM8OCB+a2CHiOuY7P07xV4LfhR8huqfce5kTVaiVXhlZljBG1dRrF86dQz
azl7ngQJNniGGqCYr2psVhYkt+cFo/tvYa9FEAuSyuuiHrWnZKCPQoQSCgLyno+CFTtTsM20olCP
l3vw2VrDLYqz70FXSFqdZr7GaZ43fCrrqYbEi1vTM6navI8YxzPJiLxxkHBUXhNDjnhAE4qxkwSp
TPkD9Klifmg86u4EiDdLPuluMEJ4SgTyukJpZvSeOJ4eDZDb7BR+xyOc01nVDurPtCSqdddFBG8J
KgziaXQ0YVYqn3/S2OFUJt2xyDxkaFISRBXWB/P96ND8dZLWEooOB2T3vW8gcSOkjOFZH9NsVgG5
jcrq51IIFnGwU241BMzihm+i+QWqC1Sr4pCNIS9vMmCV1LAQI95JbOiQA23XBlVvCUOeh4ZR414t
tDrs5Y6bChA0L1juQWDG/QbOyPHKMDRTjPCKJQTbTw+5OcXdqmTGRnMGiNwU760j1Mx1ZgI6d0WB
PDebFz+Yv+u/seXPvKmhTCHtxHVSzqfxExM9EMczmNTCTb5VT/2v/WZkPUrRTL/cB8rxqgOcDLZf
0GROHowVF/NEv6kbVWSKXv0e9hze2krZN2fyOXVWBJERNnfGWNdbh8xP8RP2fbkQ9ay+Bvod/Rm7
TRFdNdlwZmwxX0azZ6bJ5RzCnnln+rsPOOhxeFCsP98Qn/jD4s3QnsQpv9JWGf5+UXw6PxahcOIU
XBQdxDf5cScFf1msTuoUCXrVAKaek6o0VbfQ/I2bU4oyyFJvYe9JThCzzJGmiXL88kvrXo96PaAa
6fyTmhxtCCPKrIEEBrDSIMQgApqEfGz2lyNlrZ6FdZQKJkgAZoe+4WIX5l3l0s/e45N77nODM5vh
Ogu2SQnAlG7ZbxQSWCchCNo2QBlAqraGHHhYNkPSqhnDX9DO1O/S9LdtgHjA7iFDqRPFLbODFfSD
Blk/pBmN/s45EiMzapTXG4btAYbPjtRQI36wqnh5auKzmBlIYGyeVQNYOb+/zAJaTu6j8yvtKXEQ
orOoePNx6rzDwrglI4hgqsKcCI/fVKjGBSUqkdv/59Vj/HH7H1uDn/NmasgtGO9lK0m6WJgTzLEF
WcngR55h/tJwT4cQpU8y3rdFTuTE40+6O5KzZ8EaYGJ/tbZXkA7wAQzI95aTBybHMnNNvdo/8WfR
rZl7ctafI3SFbrlYFphU7ggoKw42Fr4IvaYfvUoENYKcJTPeYb1/V+PRbhVPKlnGXk6Mo4IBVF7j
QqnYd6ArjltpPR+HI5+eztMu2B2CqJSOaiqAkd65KIRjVhGcKI3vSMtd/nX0X/tG/M+EjP6qHN/o
LddptjfErCN3t9kyl3PCUvtrzB2hJvel3I7C6Y+K+mAolKfaeLZkO4zWqPdjGhqoS7pnLEuOXP+F
EwcLL1dUnDPRo9hkcdZeH5pMYl8b5UkaCYp79ScczE3A+JjdXjxS5Y+QI9SWDenZ81aTRDZGRxlM
k1LOBHk4L0/M4J/IO9Mjxf3xlHH9rm6fPQPjwi7516GYIanQLVg3pkYdX12aL5P5IdmX1BWWIfyf
cnm7IRgPg2KZopo/R68L+o2hSd4LHneNn/MCJtlS3Sh2ZzcEuNDFUdDuleDapK89JAqlHqEVTW4H
Wi0QJf89HcY9ji1HugNc2Wn/mpLCXgDNhG34sZYxdjXzzf6oMI3ZSgDgW49IOcQ1tN5CcTFWItb+
pphQa74Fbzax1tfACwDT/dalBn6lHAku6nqtt91q/y1sBqavDGXLH+yj5s3qU//ar4PZ7kVJFp6Q
op5JBh/Zn1NbhBHKe7SqgcIzc8r3KVeAU2iIfCsoDhEy+4aVuqN7wJMSQidcLubGdmA8+Pd7ABki
2twILimtKsmYaCgbWGDFgHykxIQUMQRouJnKpJOkDrtyr4KqeQ+wjmnTrGu67zh0siDS2fSYIqXt
9h4AORZTblqZ8oRtiGHkRLdvqnDB5JMwprtQd34FmRg3UkLfHHRhIEk6AfccWHVQZODtwfxs8AfW
/SE8piLOxsXEhhhWhr/xRBRpRGfGiMGkYVidh5WimL750WP5+D04nrn7FfYTZGpQmVw1CvcyKQ3B
7b5YwbT5vZod2p1DqKhNcAfhV0i+wA8TAequU0x/SUsjY/LAw8f4Wrmfhr/IToBqBUpVb0nZUCEr
lSRSbzQpFbEqjJQV/07tHDDDaF02AhMyHyXwWJu43CHPadpzUe86DlOMrscnb3S3RmhYWZAKo/Q1
f8JXd4Hk+60dP/W4FKwIgRcPiTEyyN92JjGVDcUbx0gU0PdcDeGHwb8CndiXKUA36J0+kf34DaH1
sI+TCPvLQA3TWFoUY+iswYM0K8AHOekAkgdpidP3hNX+I0/fafzmi3wulg3Fjpde8P99m3z5d15Q
p0aRdzcd2X4WVDY5UCtJABcW2VEPgwLFgH1dNfVd1IU/OZW9uilwOdhblkBHRof60Oo81If1qo3D
Ik8UeTyvV5uz0GQ5l7/03/qtQ0Ml5/RhiY9OzNt0nKNNit0bYnf8sMaH1igr/9GGRCLiZPYo5UUW
F0A9fiqAECRRG6LQpaQSSa7gaJqGROLRiI0IAIWyp9mSuRy1NwpV2NPPJCEUIwdvJU9x+puN4fjh
QJsxa/w0xkWI+IZBV1j3rI6Pq3KcPHN7U670fx3sM0WU5YQUudIawJTL8BX52E5UXIHS3JeK1M8R
vo28tTNgPp/ECAZM6nM9/RKlKXCnSgDPNvZUGiRZujL1t/GwSP1dHlT82EA/0D88iL3Phf4ndyKg
4CEHICQA7Anihazo5qX+6tIpynF4jYVSv1om0CW0Gpj1jgWnikyMBexYvwdHYi3/t5mSRmLhJcYY
OU8HssC52+yQszAsvCfSYCnKsSGB9QE2sdgr13RmQgXwV1pMA3r+LB1W+mTvjCJanBeSA/8JXcky
BQs4bpRUjbas0fq7UoBAhe7AlM0WJEh3GoyL7fjYVKz9Eg/D03AzrRPlM19beoPiRdJNRz9KsukP
VoxahaFZDeaS3XN/HGNNJj+AE0GzLu/h8hoPFWtRF+1CFsha8O8CN0RWSaP3O2PtSC99hPOPdf0b
Evcw+EZ/a9JXAw3QGu44staWz+PIy+nys4/U5Y+jCFfD5WeWdtoJ4Fyf7DjIdCP9KW9eqP68XBJR
t2/dB/HHWq1e+1rEyorD2TQ6blyCiRezJWlXxKBrS/jCNWvo9e2Ybo57c12pVWcvUxlPORRDO1pz
kJjU+/lFgLPHnp4qtV+FlSOrCsOtKTR+lqo+b5bfyTFLHW/PzvZjNnGL4WMRythdHO9f0FELxRKt
fywTpnd3fFlv6k4UCBU5v9/o6zMzNEfScgA/dVyiN1tJNGoxkFBIf/tlhnEZmtS66+mtlkGD6B20
svXqmO33soiKZDLmwEAevSMZZa+CZpJsae+AtsIRVtepPpMH0wOoM1SmOvAb5m7oGCzTVDfGiPNe
6gTyRvqMstaSlXBzhcj4tSi18wmt1jeWlfLcMABGjqpRLJxaQZP4XnnKgzKqj5T4800Zha36lsrO
SMvimoQS0QFhTMpLwMwHbKUbgoNep17/M/Ns5ng83YCgohk5OqlK1HIcFihd7K3XDskjcVxzdlGu
0Wk4S3MiKxl7gPE5wVYiCNWUqYxuDVFRU5HSddlvWiMDVagsF++ylRLTts+X7bLt4iRU6QwEi/Fp
20T2ZsE0nkYGS3F2b54X0KxCG7ms40FeYxaTd1LWICG+esAXsUP+p3OGDKJJS51J1mTJ01kGnCrx
Z+F19cYEPqWGBNvrmL1eTlDO+ZuBpbEWHF8CvLoprKPd60SWjFrEOrLpsRnlHOQsvqBk3WNNvihM
oH8H0KmOXUsrSgu6ODt2tYv2dCtNjciGRQ10zMBjg1yAcU/Am6kJrfh0dMTgKhBF1WRbBJEKrMhO
av5EAWPJorw+h/7WUojt9jOJDjgfMxhxclSxisSdTRUDJXpgtBeeToQ/SSw+0xujrog/Sodr8w7r
AFRUV6YPftbiCCPPf1BAYCy8PG8LlsoXgkk2uXmc6dmvwiBjO+vh5QqX0QDwx/tYTDo133vKFRzT
ATT/pc419nUnfogLun3K08nL+OQ7sMO8FXSCZ/Z2IL7ZHwTyS1HIQO3NcARSc6mJTP0iojXGgpCp
QcV/J5Hqf72J7klbRVwqvEv7a1zEK5NjUIgCT3suFZqejJADSNxKe/6P//s5b54sZfTHhVfTLrPF
LRJKMUCGd7Lzv2ZHOw6T7dVFWRiO54W10ygWcioH1f9z6R7fxamDtlQHF9l0Doz/wNtpTpNqoN2J
zEJQ6CgymHfxE0g1MnRjDmRPws6rLPGug1PTO6aXtHPBI3yZyZkev3gqETbv0DB98G5sRvPR0PLs
WgeTrsnUuMtrK8aNnweGMM4ZL5ptHo7O6CQ3vKVHOj5WhvlqnJqSDjjU7H/PcONAxYwN7TFcaScF
x9GkNsXG+ZAPwwbyz8pzA2CKlbBfu8GMEOivDsB/+nvpU85ph6mQsWt0AdvuGQxcy3w5MPzk6mIJ
SFRS4JnWCRet5QH/8r8F8WBZ1jY7mMKth0tu72yDc8Czcx7tpqZfPI7ZnbKKCRt+dJcaS6MoMQKr
L1UP3dCgXIZrGsxjkHZrJbDkBmx8nXxDT5VhMgsj4d3uXcIT19ZBekUyzKdByQFztQS2jrss9zom
qOHNNeymxjhWFE16fYNie1XRzuk3WCIylF4sth4nZNkCH7/EqLHJCUP77m33rZeQPCEp0UGlKBUQ
osJt5VxIEI3frdoabY+yuzGue+PKi/DTKCC3qZ7+5ZMZbHeHiNrB4eoLW053xIDnHVMRNzgodUDq
DVBuQbRy4si2K8hyD0WjHon8evxGo6qr1MXnZCJ1P5bVrsm0VTokMCHnPDDG6BBpkekRUeLhrzZo
/K/N1t2FUX26k3rBCI7MvHADYwbMu3VuK8YIC/2Ki2nIksUaCKDHvcxeEeYFJ2RH7OaYU506yvEp
oqIkVX8k9G7R3W7d5sZ2Di9ZNrw7P1ArrsoI5JZKfjjYU2oalTUDwYQ+CjSQyHRKYjZGlS+8KLOD
spTS1JUY2iPdm2/NRmBMSjkkx0YCsPDQVxm/cWLCl+P+llCQ/VaTAZ6TKoH4MqD94YdUOjGJ8ZHU
AXqF2P7tjzv8IW3aFmHmzup30aeFZo3wIMI1jGGcmEVw/32x7lap6wxjvf623pvrHkD8HorYOZEl
ahMIOYaUq/pGh/yMYzxZd/dU2/Lpc6IZqP1+hkpce4qC206m5kowb2Oc/C/yxBZWCHjDSn6058qe
EfLSVNP2oQHac8pJ8+/yYam5hzIHZtO7F8VS6S0udBubOLy/o49L+1MrrMivvMD4G/aD9VGXeZRM
BMomWKttayHzG8eyP5VzVpMQULUYkM5gRhTvPIZUDSWcQee89kDpxaGlk6p0Eg954l8EgDrbEmLD
677+qITFTar4ZBtSsgBGGlVjeMNgrmUQuS5ZuFzrFARxs/lRjnT35W32vkXbVcs+HfHBmdprRnbH
JGxh6I58BgtdaMvR7xDw4TcveJg0kAShYlAy4A+g4tCXIZ+9IFwl5/IS7DKq8TAzXQDXN9/Ml6/g
kgMw+xWBTvC43eXypOQzUbggVN9dSdeXrJlYaGqZkhyBmNkXPNMhuBa2Ho2otSZENCr21AVxvy8M
XbTcruf4C8HJye/QoKw9MBdfb+8vrzwVNkgZR+1390OGcSgWwsH+Lu5wKze4JIt22Uyk5G1pCzyc
ekqR7Xb+AYWe9+c1pce29xNKXqEjygVY1/yp20Zr9YkxZj6NML6m97ECcrkrLMXoqILa2NDNFhpY
LaiJJvLrywpOmyOD5TKpFMpzelsl/XkaXcMgNwsQzoEwJeVi85gBb+CoxQgGGeYwGv9cjOnqznda
E11SUVvzq29Y/EtiFCmgejHHj+Rx1s7YwyOSTlBGlYch6SfLoiDGiLrjm87NJOEkeHtFobs933Yp
uwK4zPK+v0uESZEzWq2xsKieVp7BqjVttOB62mqywt3JLZ5M5DvkDqh83eGWsTtbwpeLRI2CJJak
x9VsNFaaxwRNOLfFi6DDZGppYu1goPtsesvgflr6Zc15KUtyAQ857LdWL4UxJacJCb/RLUlCyjIw
wbSFszVwplluPhhKR5KoKA5x/A6n4nQuQxDQKP8zHks9fqle1j7xU0mKCt5Vk5BR+ghtUJ0AxMh8
lN3dd7sIiwDvxA10Cu90fmbl2o46478wgZS4AKMqwyRqQD5JICcLJMIOFY8mXUrn0rJ3EggUdT05
Hgfzx5dTZj8m0l9M8K/mYGB0VUyW4diAz00rRrxrTEUwewR3Eqw+RBbjzuO2kOPD1yjb28/BWUtC
5p6XCHOD/589Dn4UmmkRLI5M8lF0sxHXjKWZgi1bvnDHaZE1PF5mPlqE9PkzyHu1gDFVBmMhIWgg
0Rl7UDOHGRtrwh3C3tzNYXeKq5z8FOd6T3rOO8U8AllFqmQDmvHSBVPyhP4WzUF4/z47yTY+3TvH
/711zrQ0h1vFoImLl5s4pjK50TyxyTreoiUhqXdEj3p7SDNEjLm9KZr507qf8jgZZpaaP4QxltYs
4Q/rv0SC73+Jru+qlF3XjVSwEE99z0vIcqr4Ekhdj8AuIlucJRFdQIHPy9Y8zdeeNxqGczHUtMo6
XRZiw36fmU1MWFtA7STcgNm1N+9QLE+7i1Mno1Zsx6+UysXPwT5KKdSuf1OySeaBlRU4Qd59uuBX
Ufs1FtEoovzSLVMZ0MMMzfEFBpvzuZe57X0W+Marixa7UAgpCqMMHTwHljGOShxCyZx0HOYifqTE
ErSetlpgXpX6k6WOW/tutens9ZL8B787zUKhRX/jheXIsg70mOhjhASFs14BYmPRdqj9GafY+MBj
Rsxm5ysEpVIfrUqaOCmJKCOz/A/i2scikBWf8HB3GJhEvYt1x8iK4EcWBJZ/NkWh9eL/cFd1YSwn
SMRL0uuwFgt3zA53vnafrR9Kq5eCNOiExYVeweJH0W+86iMBjRJgMTvVZDn4lu6E0w5EcCJflykH
ok8clTJp78oRayJORgyU2muMSnKIepcF4RlhBlNVqsUymM2C+sKMr6SKlqcZBkDHRhx2FyIq7ph5
SVfRQfMgWmin/E2ffv/ItWtL8/5r6yHcsd/Y4eODX/wWxeD32Cd7UgnlP4VgWBVp6rOnGwfiqJcR
zD/2LJ+WXNwyMceuh6+bKdQcNyW7OfmB4W+3Xl+oKSXH66qL86+cuOM9NkhJV9J+dxH13YQv+4Qy
CH61/t1ENhE52+ZdRIsig8MtVojWeW9YGJSAwhbvYrOF8p7/DDUsFCxJCVgyhvCJJoz8pv28MQhg
yEiz85qtdJ0Ct0djQ5gW8vZW729RqpgZU2gWQrk4fvgNKVo+Xq8YulRdTqAyR+Ygp9Huyas3z4lY
cAmBube8jiYAg4VykHadzPUIW33oQnYE1ggW3NnHG9JssoKpOink46ScdT9CurNyDOOSe2y6zKnQ
3eN9fXJhRv8C64ZPO5KV3LFxK/oN9hUOuRuEz5GQfZmTBEC9qbEwtwCA6oTvFuvLtyuoePz/Gey2
B7GAy9PEOZJ+ZHMGhst6mytyS8e0zcjwl/FjAgUdS/3ObiYrA/o1BRt44M0OFlqLaKd2hsR9QQQO
sqLYjE3R8dDy0rskZT2LHWOke2jn0UNsGOmHwkEPHArL+OfjxuoRXw0HlMfw4TJ9oN3eFviAv4wk
8TZcGUmFa0IuIY9E8ifkSkYmyEnOSw21oCQzSyZ7QEq9WfrWp7yT7y06LdHI8Hq6IXXl7m7Mpx/9
MNF1nkoSiaWxr3Ocbi32i6q+k6fVHZ30OjpMALWileHzfhQXJIfeLO9aHSJVK2ihLMtYOMxkeWdU
3DtTrFEFhIU2Q7/HA+AamZuh1CQDdpAcYSbNtZO6nmsDAZXbuJhP9mzMp5dY+MrpBYFugnL7hPFS
s24UlDp0LRhcIFHz1XN/ZdVpj7mntJ3acEDyc0W901EBK3tq0OZhxnWN24gRthYmOk4CNGoci3DB
lqjZNgVvdUbAKtRNSItzn3UBM1oJeVrB3+6fM4i4ImxgFLwSnkKgIkPn4irtf82BYVLOKsrZOxkW
LpW92J5euZ+R1TVG0Pv/GZX/YJLff9maiWxSNXgdz2lMHEO55DF0XrOxmEe9BwyvZyuK+ASWm2Pi
8pRZNSp1wo/IpjBZrgi5cXgf30UAyTtDLcDBkBV/EYM7qtNeEfVtZCv20o44QTMJxMmFjAWnm/ZX
YUK+9PB4bUxW2KbyKapeCNJ3D83GqsTv24WW6022Gd8kTBM6y51F3MbMGQJ8E6chF7RA3iiHICmo
dQJKzIkJ9a539xiKi+i2HkisV6cPLkcM7ZyA6+xn1dbsgs+uf94oFiXg7IYijUgIahmyJpsKrvjQ
bhdDwH+F5DZeK6+B8qqOTMYAFWf9V9CD0ErvJ23eSxZw6wK2HKixWpsQUNxVyyyX+lRvACp7BSDY
D5AzS3vNzqE4TAONti9RWgdBGCrsMMWGY+oODRXerD+W17Xde3fIYaC+dfh8Jaorm5DG9fkINCs9
oUUWvp/gLwF9Yxo4MxtNqAmHBEmlQLWDdIIo9VnkHOtXtCeI2Esz3P2oCjcZs0K0ZIefoZZod/Xb
b7GYWx8KZcnPDuQiyUuvOy9kAPFkvpX347nVu2vrsvS9huWQXdBfP+nhFWPNjOHj2SOa6exO4GiS
HkBGh4LvxeD5+GKXvP+cze+IZdREUTYMml+oE8layDCCkjbhRFMBw6kk5Nhy+pBbbEfVvmtfNP3X
CBKAONhbMNcde6s8id4M2N53rYdSL23uMrzGnZhPVtI7KIu0GGaO5KX3GIPtnQ/W9VX6osij8YdH
+ndZbnsUbJUsxwpIoMu0L18LbiVy0/1ZERE0HeUSl8djEiVenDiQQ13aXafQN8wotCDknlAkwuc2
EQJava+2XbvTNQ9pTxC4oy+ep64N9K+ozqcJBoirXChLtPfOZldytCHIUcKZk5WoXWP//p4yv0pb
+uU9TKE1XKqh9WOHZKhtC70JuwPNoj92d8kTXtXB/UACZwFC5TD5+/sIoJD8WZCtIuT6wTUkF7O4
MnUTz17MVVDcWTUc4G68H1cAPx1/+0k7FRFRc2BuhbJiOeUfulKcmakITuAecpq+sKmZIY59Hy1M
UXm1LAzuGQ8caD9qggw10LA1t7Rrci+rPgvqCVap383N3F3EtqAA4ZlYIC7Fp9S2yiKNUmVMXfkg
HxhQw3JKG1Adie7osll+JCXERK8KWey3yUhI2OjjB4vz0eyHwWAv2cmAvIdLEelhgM7t1w5tcxLo
Bx9SQFtE7hSmBpv3XuEvhcmDEuI/qTV8TAF/EgXzeS+jtBMWmyy3MCumQ4/YbXttDzron6WwEOox
wvA12gGadqqZ/a4mahq+kpUXmtl0Z4wxIDMyugSpa5OpMg7P0BAsReGmEtkz1LB8ZorVun4ywQyI
nfVjM2L+wY+eQh7/DrK5EJzX24mdi70gdsUoWxWorAX/9v5n6Ghwo4p+1hmGOkXrhQF00YAdAZWe
IdCi1HdXG/r/CNkVSm5VuiFcUG1/VhZZsRrgrB/T30UAlyG8w4vev7l4rYkr/LR/a4FWYIUhJUCd
95ZIWPfI1VluJAqcOoqLqLfcshptrL6PtVN6CVgS8SVM2CX05hOjYEEZj/3O4LzWj6JdLSlol1KI
xj7/5x8cvMhwC2bzAATAyE9az1bjScFXkubqod9PeH3fEqwL6+5mITMX/Ab3mIG2gkQPre677wJB
/d6jYEg9zdjgZaFey+6djbvtias9NwrIKcH3gcWpWh4NKjcvuhH0RzX8AItrcw47An9qOZHa9l/z
wy53ZMzG4P6ZoPn7bjKn8grozTdf6295ISUDLNsM/EqoPjxZDALN8gqf6ZrUtaWiWx8fRMMc0nc2
SncSi9Xa5tijiayOn45GF+3/OB7wZXodPAYHV9krRr0mHeHpBpdp3S+RtHs/5JP3X/7bGJeWgP5j
UzrZfmlTrbJfMWYAFuTTbXAdUYticqDviW9e+Cw7chAOjBes9pWOKnODMet7P/V7DzuJ0LoogX9N
5alq7aCSMjizkbFXB9RxQ811ZhQ2Al0l81Bvo1palwYogFJTzk98M7c+aGbowELCeMnaq4901qw3
xEnasb8gvKMzRKquuoMylN/jGAY8Dfznt1CF4vqy88sgreTUsQJODfjau9Mz1E/23iWxK7g9p+SL
1MhFC5EXPPEmHsJxyD3j+UIl7IyGHSL6A04tDh1vx11tyfAGHsmSl6zu/bp99JB3mpu1eK/niNT4
OqMKtcjz5t4x90HbZ8zWOKkkNIXHBddPH8vLAP/y+G8Io3tMmzZc+LEBAbRVOSOndx98dYs/fO1G
P8a8HzBC3wdb+MrlWWnPEgB+Dd3+etD5J+YLoNvb484xWLOGdKvd+j63kBbVpigcE/n+kaM7T3yK
n5oAgiZ3KNpyjQn+DqfLmqZi+mE/2RjOYW9cAnntc4E46Z3HyUkJpV1x+2z3z369z7RCn5j195sn
vyoQ2vKY9GcsynfTbQ9FgxQOVyF2pY+FOsT+0SpGt/AE0QYVnmMJAyEfZgzzBcjV0m7VgPW/8AZj
eavFsvy2l8Ax8PKIAHjBwEmnChhyR632FmiAMrnllkHoeJMFG23jlYjrMSf7AMH5U03E/varbITQ
UVAWwHeYLkpcbYgq/QwtgVbqtaGEr9aAxNpqjhXnl8xqiFtibNXIlFRBfCKjk9L961L9+OR86KHk
2nodDfgDK78sxzHoHmu3waXXWyAivKIly6DhxMpoSMHSdtFsQk0mBtLHxbA6ciwPuBcxFX8ekXBF
Jrlnr8w5Xfd/8g/Gpuq4ShDvbmfLt5IxRPpleXw5PHr+n/r8J3i4n/VShr/z7LOZaDQgBLqLNyMi
SSgGKnmBMqL0VTcmYHLrLZuu+rk0sKvYEs41gNKXXuDJbM5tiEJ7ChFRnkbf+enCX7oUPqqeJx8Y
4ObSLTk4z407g3u0tHwYPMkG3nhn4iItg+wBgnUoofK1k5sAHBpgzGRUab1ITZlDOqM1aW8I0K9P
KolG+wMflDna/x/dRjb8ravp2pxKtHeSwzHSpfcqDyy6r8ulPyg9P1gq51E7Cs4v0xDEDdHrsbaS
AGsq962poj7b/t+9pz2CF0oqv/uhDy76xt9CJui6bOCQgVCXm6jwFAZBbFLLBNVD/L6uNuqPGse3
AlHJKy3MCtipv1uubPjBYilWJHv0+ihHnNMPRMlARkgOkcSowgeNnCnmda70BkmHNITKYOuP2G3/
Um1PZjX/rGYhZCzjBi0o0ZBv942jMPd19i8I4xM7BM9Ubgm4MR75/gge2EX6hdQ1o8x0zhDWX/8G
0lBzujY91M0XFETQ3aa4fU+ciYGhzh8PErPyKeN9GkRR54khXaaRgKlBIEvvnhXxTCKzEI/JCoWC
SwZilg+JikMxBfjJKrJXz3gjB+KqKj7vQSOXw6JIZ5dXDjRU15tTQedPDmn66enZCF2sstHUciJA
aCP7XHHdlLosVSaatKZMJHPMaCUI1IM1Ru71iXQZAXMYDHILiSa+CGk5j5q9GaunUO6l/dGX78TB
X4GwKWGumSeKedOTdQ+9IUtfCwnQqZwsxn6nGrM0phMoiSoqb4V8ZjajZeW1lsH98pNwNI2IbROe
/hhPJsBNG3gnlMLtnj5LkmMqxFUWWZpL0oGVujKlqPfuzwKDPRjVFWOI3MgL53CJkPg2s+mJ93pc
Ho15W7sb474AzXpZwX+dNw8cKr1TomJuKo3BFK6eZJjRB/ef7vCi3mMZZ4DZvlUu1ta1+jaZgfj2
SHGjyu+2JqBokpQEY+xPfvU//kJZAKyVav5wyPSGiTd6g/WtQAXgGFRchPnBC1O7owNf0JFXK++j
RZkmWjP/+LflEUlapqNqzl8A+wwmA3t7f8DGAJ5ISw1NBh8/zAQi7M/Fl4Fw6DWCwy7NRB9ttWos
ZlKCmKxZbLWptAiqgiHaB3C3s+ycm36szp8ltxevhvyoUrlDNdzVweCoUws/UaQjHmnFTB5y4Lz9
2u5lPex2h1xyn1L1ummbdl4UqtccqHE6z+RDinJOr81nR+Xecey2NHY6mTEsbt8xlykgKEW/t/iG
ZV1v0iyNv2+Rf1owLuT5oJNN/B9A+H/Y3MteV43bJGD6F0KjmRYtc8dEg5kYYZqmLKy8ErpwnlqA
n9dvPb1vtwIOUMu/yJ0zLsSQfYAdI86yBmKreumK8Be0wKQaqEfkz1SGWEDr1QqR/DjcgOLqTnjM
dThHxR53Wp3+lCQCHwbPUPY6jBMfc9TUpOfxSr7Q7OAnIWgvFpVdqX/duyASXYF/mMxyt3k549Bv
Z40kCYuLll9LrUMBrXOt6vV4ureOEUODbRBsygcftsia/jBDvHtMGV5SHa1RvI2qCRxIkfPoNeF3
6jHBmnsljdzmTaY1mBTPCmuP4RA/q1BWMLmi9UikdKHf0J6jjEol3FtTnKWbD+IpRAbwPVqisuYR
ZqdadGp0yzpNrlEnO6Xnib9GWMqnpdKCOCSOJX48QORl+dktVW+Xfn502Zlj/KOyNum0ZSDmyrVY
Mj+IajRyFmwLIytLLhu6vapBV/CSys6rZhl4XS1NZh4amzirATc/dY9eFIw5dlN3qtM6LH0hfRe8
ffNYhDumZrBGsk0GfNovtXDnE+4uTihHo9J4OFgBRvA4GGKMZ8PvY1DgFawzUX7DldZHh/jt51Lm
UQfvU9ukdAHz/L6EXKamJ39yaA1YpM22KNC9PsNIXKbGC5dZbIM/GVE10gfRv28nMiJgoolzxMCH
NC509PA44fUHRoS+ZQDqYy5KxqLxcYa7XmLBHGL+nYJQPU1faVoLSHzpqtglnNWKf3FQZznP2kI2
1JidlnbC6BOhBMW9p/0RYy/ogRXQPWUyO49/CCZNIFcTCksMwWeUm+XQrurMmclwK7Igm0NaO/xZ
aI+/9WkrYTc/8y6lOovbl/L9YC0Zrg8bxTY0G6TzoWYKa6z8tBZVcnU2Z5zGqUmOcw0vV3ExX7bk
xXkVZCwklDU7VBKBzlDf2V2wSW1pmY3FQ5BlBleMX+z43TkOShajC5zFB9qgDDdY63S0B/SCNE0W
Ad3Rn+ADQN3xHoxBBPSzAbDY4ZfV1VadO1klYtS0VfQqITJLspa4mHkXVVkNOijIwT6aCsVsy2sD
jNhi9jnsC4deuJXsMo0J+1xNmpxkbYZzuY0B8H4Mmi8aZw26DV9aayhf2R3B8vIKAWMmq9Jw3f+8
sbgG/64MfUvdoSNvv+QjTBSsxUb2uwU3zMv/lcYm1QN1lGQGOC36e5qdkogzZOZCT7g63iki3W+W
lrsocxSKEtiDo54QMdMwtf80zOKJm2BQIaNW0oHo5dd8cO5SsWA620j8XvV3jyhmcAT+kcRJjAzZ
4OajQhcRbiZFRREsDRlORwmH2TaVKnlwBQY38JCGzL11oTDyNiuKCoNT6rP6PRKjNIYXRc7LZIEs
cqQPTix/eNSPhWPsPCvGGCqbnYbsWUOn90E3zKYYhlqdFnTD8YqHbhLlf3CE9EIRiai/BqHDxiZc
JiMVTsN8vE33JTSWwMcKrGWnjkfbZFguvMp1nQrMvi6KDvZQoqg+bR93cZoIV7pgP5R16yJuUIIS
P/AZElCJ8hKBCZngrwwOrqPkJcwFRHs2ResHaagUqlSKpVwNOSP3T9WxToKG6jqMyFvlivXI/7lu
if23RYdDBDq/Kv6GhpS8oN/Altlm+ePenG/I4pNpWpTJK55+hKOaP5d+0aEhYymD6PPbNY9DYj5m
CyMBAofdgvhwwE/FxZyE/jC1+H2tBQ/ESaZMV7JQl7WRVl14dXUNsMJaRbw4InUoaezJ533fTXRS
4dZZUSEKnVmRphN9CquPQaBWALzR/t8kDpVxJatALO0E4Up/ELovoiO9hDHR0GOc7ultrVWTa48J
UDJH3M/cBwKf5onocST6Zz5nEyViIL2GegHOk53kLupZwC54PKzvcmDBsSGT3a8QISbGt+XtsQGM
su/zY1m+LmRZ+eNDoCC/R37PEMtORBTecnPbVZdh8PP2v4HSx6Va6E7RKPARHq7E1ucBZ0gDx6mA
u3ys+hNEK7i9gK85KStstKckQkmD3RAIbJ6GIaH8AZYGVZ5sQsf0m7tJhK0hQ0Ba9qvS3KbsYwAo
KPrgkUB6HI6G7/gxFWHDuh9vQffVy9MVJco7KT+kCis7/dfAEDf2ON3/5pMEYKQV4gZgAzwyGrtV
zWdkZKI859UxmQCXufbp4I61acWEICY9+ZK8YvJQeK7mrQEFS10JXh1Lm7Pbiywf9A9hoeZ0+uOO
7uoEqIIe0sOlMIjtY+Cb97geoLAg2uHQlIIUXjGqYS7aqo+aNTENXbiMPyIQ11OUXnwWK7lcn9dK
fWL6A2bWPljT266ltXkNYA+wH/s8QIVwgCH/6P8Au0X7vhkeEeh0IRail6wmG35RtHcxOwMFiQgj
kB5ZMt/vZETUYckOOfIV5PYxyCMmaCNEP3ok2YDv/wAHi+Dm8Dfo15dtvGHSKM+h4RhJQujxB/KF
Om7zqFLb9kEq1trp7WulHQ/crTrxtI05LBArUaoFQjNCaZ/WlLGbZfV6T0zSq5m2Z4mQh5hgopQx
eD6gxyZegNWviO4O474XJZ2eF3hFYOp7fSBC9HmWLlumHU7T91MSjcS5oWZLOEkQd57aG1F5Xad/
N1rukE1odtJzZqB39lFruSRM3Ypip5eHHghlq53K30nH1jTx7+mUquECSgZvl5lhkGYIhwRmYUc2
+gfGQ0TxsdXy0yl+HF+tUprKUoQVABzgxxCV5cgoBRVHKCHejUdxRKnVtvdbSTCy0qTLYHNlGTV1
7AMkZxhoe7ctUknH78QgryvSDn7GkvPy8d1L4dRA+aKtPk4ssiW6qHXii6mgO+xARGUtSZy+TtFN
+FLVoSXyKhQYeXKD2QzC6UULvsGFDSDv8RQ7RGtSECP0bs7AEZiqWol0Wo9zUd9tCYZQo9YMzSXK
8fULCc6ylicuY9dPPzoz3Jg2cnrsUc0r8gkf6OLHGiwhPtq2wnN4VJENwIM/vgN/Re0Ce7OIv4p/
Hht7lzs7m7CsyGg/uzINT8NVfIwWEEQ/N+nO8p3SRO1TdalsAxwJlJ8sZ4+ZEhAdFwxWUuQk7sNJ
PuPlLuns9JiEyvhafG7T9Ve6z29GPonPCxUZlNyPk5DVTOy4PQISZGcw9F/lnRSWjfS2lQpXMric
LnvyWzXtHCJeJdLj7F7bm2nrmQDE2itFtTXwyRhPTNQeiigFzAeg3nMJcjBjpTO5NuC+8ogz2leW
9KpCF1D1Or3+LEWGxUs95FKrj0hVe/2cWmWx0884kDXSev2DKUmSp4CcxWtXUs54dUTrw+ztwuPb
I8JNDxTFZ+KOIYfW6f63tce49QH4ucEjPQf7x12BFuqq3DuuRXxIEdc0T6el8fLhqkgOSrytFDdf
B30gYY78898f+zswbmcWlAFvpZJ4oc4TufXNERMA94kV5hDC19+xp0I+IBDt3FAzMDV9ndB2jyKo
DtaabmrjUUijTrPfk/ye6vBwPD/94k03zzIluXvoKjwIvK3b4Nm0Mk/go38ydTDRJoMDegYno2CG
QVn1ptbH/Thxm2wL0Ec8QWvZjLTj3FK4HrMPj17JDxHRzChCKTC/eH6pN8cyEVsQ6aJaAhaHXFjH
TBvQLZB1FDjAKtBf/lp0M/dA9l4bYsCQioKa2q1XScdGn/VC0lXVhORTO9V9v4ZXAOzn+TLIQhL0
IPSLbBEgVhRMuDMBbY6ABuysUkvW4mJ9t6LG1GIpniBvkLPYZk8RZ/p7y/YpsuBVcnHn5Ph/9k2w
GkG08UNmk4yNIAtF/lVwaWyTg9GQaLZ+My87RvYayx4O6u7RsHWPlbgmQY8cZcYeLyrHgJGhLDNY
Cvfr+mk33lJnUOq4haYIr4NB5fUi3so1UDIUhHi/VTd+q/VOgAkofz0aklJQgZNSga8oCnYeUW9j
XUngLusPJib2GkdgeZDw2oXq0rABQw/AaH8FUEv22j/hSHMTYzav3cIDzw2Mr3C9n8IjT83+hj+2
XJPUJgsBbTFDv13sM+3fVY+XctowlXgXZlBQsoP0xnrOZolNXRw774Jrc8+8uZJ1+eyKnTcYdMbN
L8AfsJXiPQt8yt741ALgvnJwk83bSN2N1C4OgSmWDG5e6b0bRBE+FDlTURagEFmSR5XR9jNFNydQ
G0XjQZKMh60dPEfSEl2M7MqktA6Xo+PekkA1qcg1jR3Z8pzIlmr5YR0+ale2ff3tjB1N8cDaJ92x
Kb+sz4Lm5Bi5RgIukKpuK7PlRxKs1/R+g7+O+XzGXyxQ86Ouv2nqPJV2gFpWTJNbywwmEfbG+5TF
zrRh1jmwXuri915sOm9GceAFsT5Mqm/oPgJKbF0brfEn1PR3QExlIvYLfosj196LnfLVJXLVzplC
kRmelCDb23EUzsWJkbd3ICNHJLOYsu5dEYX/XsJwGn1Xj0qbhonPgC3St6h1fhHz5onvmr6kt7XO
xT49QACwSd2rGwXa/nEUTeBRa/nGJvOVlANQJp/FMc9zD/tEVu7KENO0XX760+yEaN54boittbtw
jgesVB/U9xujSjNxHIBO0+L0ZoSC79DVdY4ko0NonrW/0A7mMMEv5PSpfqIawrYvh503WMTMrXjH
sE84vvT3LuWQrVd9VWSTUeGbh2oeV7sAt9BGycQOH32Cp1MxofThICS42SEJTIYDI46qg9W8r6G3
r04t6rFG3xWSikZlN2rtRZbxb3CprOlQ6xtJ5Opyp75mMA9XUpAO4Vkq1YSkpdksTOaYE7pZK+He
ENrWTl67w9PyMAsWaMYv8EAZ0aA9qtKNa605Da0xF33ar1D4m9ilHpryYvgVPNuMuDnjYP/asSBN
g531HTDGjsmU+Yhm3asJUSIr9XZ9zQEwPAXKg4DEzcJHmDGfA0fAkAP1SlC5F2xEmMI95xVwXy4D
jja628aax9XbGSeLtHHOcODxT5aeYQPlqvSexD523IjRW6q1vptfr/+cK9Q2SVeM8453RtHVw5iK
K4GAFK6Iis6NDC56hkjheurrNC4sASnufntPek1T0jPEqxs4/CCo08rHgUr5Ow31gf84mO9X/i5f
yBR+Xbt0TFHyKWP1cAnylr2AK3euksR9AG7WHzyuGPZ+dNVvpyg5oOesBUu09zgkpfzsIS3G4f/u
gQo9M2jReWlPRHSvX+ekTdeLhbvKHO2RvzGu3SoZehpXVFQQXhW3oN8/4uvCFk8UEOMcY6JfXmxH
odUlmTxzYMsZnCuGT7xaLe2yt8glCa/2QabK/WIdEtOOr11XkjbbzM/xwa0ruBSgIuoKYZZkDt+D
3dnpHIVVrrnAma1oAgNKMbNI2qdjfyCV1PE5Y+O4bHzPE6vndWXzg/W/ZkahCzeao8VH326UmNNa
am5h63ifNHJkThz/2eQAHXwevpensXYew1q2nOdjOkh5jrfDhnEk+oBitWryawBBwcCGWzTdNLlv
Roglmqkvri/9Lt9ppo7/QSNUekeMuBIscCrOgiP8W8nu6ZmLaJVtnXvbIw0edn5yuR8TZagZhoZZ
LJHo2YYR8/TJ2zyQj4PfmAENudZUMSfWzENvAJ/PjKGhVvLwgtRfEv8gHASBCSn3bLMB8J3tSpMg
QIE/n20djeRZJt5sxGsdAkz1LCHuDyvahQBuygcmm/r3/sOmuZNCuJrB/qgDo5WCg5fN2SKwrcQi
UifEsiU3Psd6Di4qkBnXxzooD2EeTPVMMgvUC5WTochq5sLgLsXk02O2YHF4f8yoAFTjliGzyX41
La3OXIRGMUYmW6yCIXHKEX3mVtg6vV/CQTqc4WewVEVdk0pxyXkSmBv/2ricLuBb5nQFsRRfDPRn
PksekR0v6+SO0ei7hvzie9FpNnp115UQPdgqUs6JBUX6ZiQBr7BSlmqjUwYKU28l7PN8obEugiQF
DPjVRxBHyaaX3EuRkEqpXgQ44EPoViG0Cy/qhps5u4zxzXxwn5bip4d4wW2wce/ywvFm1o++pGH6
GjCMFne94ogY0I2MY1sd9RqAVb8jKSRKqm0phM6juRmXoOTr3p+GG4obUpoTEMde/3RXZqQNFu61
JDhI2iThBnBvSDVqSk/Uu26MDWkwa+jgHwFQJRurROxbWOlFSJcR/91xOfD1xlXONuFasADMj/q4
jZZ5GVGTVHANnedlB7uLRIMKsLoe5PaLlcKJwlsL1rjYWnQZ0WNm/BECCh51Eg+DbvHT8v2UOuC7
ojMmDyog5ujsQG0J/zWaI0MXUOYYLCbm3XFm448xUs1Uht+Dae2YOdtnEy3Zr/HfTw7Lx0qQY6ao
TLtyQqGPrPMHf6Hs8wck1ZRPlaPFfjujxHTcm4Kc155hBRs4m2qoAJdTTIK3Q5l0n9pRAYYV/LQx
sKjZeV5Ex2AzQjyNY5Xmr3+zJOJyJvYRxNCuP33gyQMnmMoNl9ZdgKFzi54TrM4T+7YcO+3YdaRN
VGVrpXyysFiBGgjgnRZwvybmAViUCp+4tJufJ7yjgEcz9UdO25GL0jkbDhxQKn0CnoL/jjxDunbQ
ShnnROuxylmGdYOAn3HvkIkDkC0JR8as5fv43NYegsPkNMHT47wWc64QqCnwVr/XGi1qwt/brKzh
L2g7JNhrBRxpSMfO6E2oI9LytiwPn42XxgTymV1JlzXffKcXuh4OvmYOAIXCtBij7xls23haSrDS
Sk8MCiUM+5woo9ZxwSBMlZzzlKDvjJrI+mEvkpMI7tzxry4S18X0mR+9FTH2WelWnFxA02W7aHLN
75Zfn+Yng+ByKsz2LuO18Ee4ZuXMF7YFF6a2RPfHjFMdQiBWzxDMsqDBqTi/q1etAiKV70YWS8as
A5O5Obhd82np1vZPOMpJLjW8S8mZFqAQv5OTVfclLO9p2uGqTu+d3vJVj5leF7whu++YNxaz9n4+
V3RkuMbQPKzSn5scq9snQ2p9Hbxhgxtmk3IfnYtdDJ32Y3smop3a3SllqGMpIoNnEC9pYK8/c0zS
EDFd4aB4Acw6uLlsUhpJHWDZabULL1pllTvw9XRRKAZ/VbTTVOGWRZU6d3g6pGkdgQ0h8oYqSX2B
qLrzanrToY2EnfGCahsZNpgEiBPg9YleN95EcbZJImlm+KHddjxxss8ebH2FoDErYHNDOp231Ebs
vWn9We3Nr9Ps758KAGoNDgZH9cODQFx0uEBv5lX1gM8LauzvekIte2nY8XcBy3bGtFm2I9hnte5L
bQK7zS0KNc/Ndq6oJQxKnNFv04opjcVvY50Pp2fvQkZmYK4wCqKK4UL1wj32yK0Boskq3MOM5Yq2
EO8/DWYLj+tMERauLnWOUsA9M3U7w7W0L7PjhIcsTUzijqDCtvrPkHC5feU1Scg9eX90Kipa8iVQ
mRSIxxtoOR31I6PY+sqpt1wZStAchop3rlc2lDkav3hkC03qX6ib2LSTZkvkh8ccGQez+R2IpeMW
hw79pPvGqOkD5eVwx2vRX/jAyzWqbfLGfV8poCwj295LBYMsckbJ4fxtOMFh5MCAVugjfD8Azjfp
1zXOW603pJK+9evVG3IoX4tFYIaqqG1ETVv+y1CsKo1VklrnoaG7lYEA/3/fasTXeoYDl6EpAm+Q
7I0VgGuvToT6uun4rjXT/Q9ub73Z/YCoZ2JwToEUP+TtaHMsyeZR/WX5CUCyxSshn16tyKP2FVpp
ivYcevP7Ew+0uYQikgtYRp9z6mkBmL4JtUFal6z24kPKZgSSyAwAH+Htoy6VUJF3SWD6cWkOXIQ5
CFgFXkfrlGiI9EeKe5l2sTylbaVES5bpQZwwapJ70rsUl2aGh/lO5ycTqmmWQMahI8DRpxXP8i9n
nelAuxsfW3MYqqd8RWo2CAI420JNZ03jjWK7wCftpvxdZTyujFcj9EjkSinBCR3A5mH9FH53Ll/T
2HVjAl0N+ANc6/j9/FrTzhQo5bswfNIi0I8w8++f/hLRGNOGjqJHNkkBqeBpK5QwIfPcnAXgSQ59
VSJiNTKn30TvlEFoiICRtDWO2MeWmNyD8XiXjz5eqL5akuFrEZTS7J6pp6KIcDR6VGAidiUYp97I
EK+uiBGT7Q2jIzSlfp6GGhE4+LIgMh+rG2u0jMWqPKGZVRLR31QEB9M91pdn1LXazgvu5HjjTvOs
FiHC+YWops0rd4aTJGTh9nQPtOJevbOZLRMAA8y4AudZcFwG8qAdYCctdKGA/kV+12Aig2T4saO9
S177HcQGMixa3FGDCh/BPapTglK5U/62H0TOTVujiw7ZKr4pZZDsHNSRj495CC05YSfimxB3W7oX
bB7cEaAU2hv6+iBmnZSW+6ySReKHsJw+PFxb2LP0C5H5xXB25izNu0MhwfrUZ4Thi5cF9w1fYA0h
n51x8KXdvus45ekkBxpiUDF70Po+IsP+0qHwvj7bbmOpBp0FTRI4nczD1fMk/WMpXF10F20oLp6F
s5yp/x8RfZspHrSj6R8/YSBh/eV9NOaJU4MhelMvNI9Jayw31LTuePo8lVwwHCwcvwWeh4ECjJTF
XwffR8dQdIyvxioxrb79IBqwgWuE3vtACVJMQhVEKe18WnBjQukKGMnvHtlPwj2Hck7qz4IDIaD5
1Q2kMa6FXtZRlTj4qACReoTynk3tNb/aw6gXPCPTbbQhEWncvcIQvj+7dc8dFJj5pmUY0FtgePpO
aeIZeae4aTSuYPXCVmBB9t04Wm9cDryDORy/L1+sRR8bjuDgJE7NW0/BuirSEuYwahifVEeAbose
5ipxpAnTCXUKdiGIyHks+TmZ15926qafv8DEV35MIbXBfy7MLo/QUdnhiNTA93ReAldmbMyVQchi
4wb0SioWJ1JkgrtAeh0m7EK7wWlmUakIMJfin4e1L75T810852LaVX24UvvNJ5Typ3d31oDA3HGh
j18wYPEQ2BKFED+U4t1GRcbkI0Dc837czKg6FScCbNX/gp13j3Vde6zIGVoEY3ccN7Y9wuypCDHk
641v7hmo0Y0z0yqrfYAwwOrahY3PlSqlMijBF1NUJfguZjLdo/YVyMN/o7oNpmkvj53hQQBVsKUx
RnT4mSrTNMJnHONtmybKpqCKdq0+Yho8Bbgipq2Ckdpppp2GKi8+5jB/S5Qj/ww/jIgKLVIov3zQ
8c68Xx0ZEa+gE6odUO1uSvR0lgY6WjijW91ZD4+dCs1U03oStJcaCZuG6Lf3GIITJgDIXNO8L3v5
/FTcMd+HOaUCJ1imylbEVyI4t1D08oVgS84+B78j5vNS5O/FtnVJs05QQykYrKLKtK5+Qh7zxmI3
xUVN9qVx2oFXGtdNlnyIgnswpOgjraya6fmnvAp5XWZ8n4FnTUyAPDcphl1ecWt/RLWiifbmllCd
hx44kdbhNby3q08EfH82xzwNFCUZhVPTyddUykY9AbCCYghkxqZu3E6WU5goLOsHvgwG2IBWTFx9
S0st3KbxfjXZk908pZ2YyA8FWKbJ2Y+jxbp5BFhvMH1uEZa1zHdxuHvx7AAEFtJB4dB6tKmWbnwG
UHjfGPADLS9IhrjCDOgmpehTEEsyeTTwjjc1ArCqouV4oItkm/Jh9Zv4vSZkqV9V8zKpGgqhlBf1
jhQuBnzi3FhoYVXlKyil/H4vSG7cFdTdugAooEqylzJLcQIXZgLTMZ7ZlSLoLAAqCbdfcIz2o2Vv
leiQSC0kBYEZIJP527l9PNFzuIPSIQjcyF3lJJofz7/szM9Nz7m5H/zeEKD9hfkKjQvxpiWH2kdP
fPjfX9zTRXt3hW6o3OdyxVH4rfFMauvpT0MwLArPo6bOQZBaZhrPv0x7E94r/Hf3Sld/h+03/Thh
0Y46ymSMTflHNZRPQuZM9Bo+n7RazCiQQh4M0coeVgXxzagCoJZJS1w919Hgn7S5oWiVjxkqZSUt
MOh9OvnBHataPTn+XFx7flCDin4VzoAF6gkRfWLcvvatpejqcZ0hWQQTtb3Krd/QeJaA+TrVNLsW
YB+LL1NvSRzb/EtVYaPTLFlH/rFAwZlybAqiybwNxw5vnIsOwHastDH6iPiYyBz0K2mv39SH20l7
XzNz4ksMi7GcGrE8+mCdESvIAfa7eZuRA95gM0zgHG3+AGA88Ca2r7YEMrpigw0JKlPyn0NHKs92
KBgZxyTJtvT1Z2NjK1wpy0rimYx2GPSJF0k+a//AQy1MVBfsKkNJqOj1VIpDHjz1srRIi6rnU1bn
LaDxDOYJzf/RCcHXjZvB6MPR/Rn5HLHSuvVuVHJs9UvRGJvRObAnOVJk5VB+/RFdnlsEMTRf0hyI
5jzRAibZ19/4nkf4faF/MX/FEzobkEniQ+UO65x2fJd+08KfaB5ROgCm5tBSPHsgWloc4/0GdMO9
AESbZtV0D7fBGAd62Unf9lzpeDnw13IDS2SJEDtCgBQYqPQQ/d5xRk90csVdnvRQjpHo0fnNE6dA
ICtvLYG1d/OlvQjXsxNb8Mnwvm0Pb8FELOfGNoWRed320FLGKxhMHLlMz4aEwy0vi8hUBsquHRGg
oP/9bRF08qIat5tpYjvqy1ux3cGxOCJGhoFKcsHpbJRyc417ndPxXib/ipKfTr7G5rG6vo6BDTzW
aAXMv2sTNOVkuUFYcEs6WCnSqCqAbWqO8r7R3cBDcDKhVOB0sIq/3sI4lBeB3FYgeCU62K/2E0Gd
mIqx+/phuM25OsPq0PGl0Q6IAkYEPPI2vY8mhNCMx7MB+I1tFbvM4DHKfqDklzXvfaEGFOp03eSi
0Rz98TMhEL/nClHGByYOcM16/Ao+ZYLIZi2e8vp7AEIL9+Ol2zQbI2osZWV29/KRneOh8n4DbdSm
trHXEGxFato3jep6GMD3WS2RhO3gSh6MPHElEZWGAu3HF4frhV/zNuVk2taWRclPbUSR/0tqSa1M
Dqyt4lLIFR3fRgki/lVa3AHtcimPBxoa1O2VoQbZamF8Efea0YFDt4GM25XUh8gqMnIWpchTWBkj
6jhjI4T3uq9M5MtQPRWnJX0BUgmweXk1RM9EJnau+lXXcouEl+ixkT4QT4ty2QSpsm/3nIKe6pYG
N81Ra91fN6AAPMXtkxIF+HNUK0k3Ue8mwoeGKwD6/FcFp9lKYiQObg4cq/YQn0GitXoioi5hrmGZ
DqednZK41n+c07aTuUeC8Cb9GulAMTUdXeb3YzcSoLoQ+3R/m/npmj+cEp9a00+LM3RGpxejybtI
+goh8r4g/rj+SgzXU//F3WO12PhHltLH7M3o+tOep8J9DTSaPHXpG+cImS8pl3DTOO4Xd0DOkoB/
P3I8VE8cpYpZAuaoN/Qy9JmZ3dKJMSHMVUCgY4O075TOnAogVlm2O0Fg4K1DJ3RYs00Q3T+aOGBu
wUpTMEax9Qj766AV6wyR3LOh/bpXq/f11dL4otbgbK7zuknreowUjx2vPSZlfmfQf6GA0CuwmvxZ
9xD9pGF7FEJLEsvk5gBW6aVZcMQF/2RbNQQP74kXQX+0YeaEK1HTguveEofH3+zhqLd4EqDThZV6
kuqsg/fZRBKYeImSDck3NtWiP0QrY9Kc+oZrmK5ZepLBD9QXRGRIMYWEOBpQpD/srhWH1b4CT3kX
EO2DG/+pnrTAytO9qxb7fLBnwScIjW+w09UxC92TpIgPE2y6WqkA9scAo/oCm11QGHxVEHPDoP3u
rzAEbGzcphpqtHaSk9SJQccTOahG9zCz93h0eEeQaIGsVmK52SFW42zJBVXUdgJzLoiz8nz+GhEQ
g8l8KDcjfqa+jWVeNPakfGf2DocSTjbQnhXvLMbvGR9XFq07bOthSwsdFO7AdaQ1693eJ40CLm/s
qGiHQmSZLGORj9zRsvpA/l9bl+NDAMKISyfZbG1xlAhF62UiDfZi925mpZ6fMFmiYcG/rMxJrhX4
hjsa4MADmxxOI7sIdeZd/s8+7SdLNPDlb4x4xez5EgBK0JJ8n5bYk7HgUL2Zw7j51ZCZpu8bXWeJ
5G8+ys1LO5KWe7zQLmSVu6byxD4PHDdFQNWR5T39L9VmSj+3NG3yEZex7AesTn13Pd2GOsuB63Ws
Uy6nGvZEKPOohCmPpn/7PTmJ8hDk1gQCRaQ14e5gW+1/PbPvpqZRLH/k4ZKWJ3bqCyx457HJP8xx
kHB3f4a7nw5Dn/Wx2DI78o/572jdp4qH6omK8avBpvQSFdtutRUxsrvHswD97sYJd8Qr+RLUtGxM
oKGL9ad3DZxanEsf4uVlydAUgs+LBxLRd2yPY6aQZ7SJV1ELmkNCxG7bKAdzNuX3gYKSf3HjlSrO
uEig7902nZXBXocVruv/QVoF5yPCM22q/or2c8/Eg2RdiuYQjNzpfSOyLUpG0e9/VnQrRD/yRb9n
0YWrEw9921vfiFElUlT+ql08LE23DPerhN5YmT4LiGs3NwNESIfX5pNcysvES0wfcicl20mpLelJ
y9T/Z1mTyg6G0bCGx+Ck8/z+Rs4n3ZIDdD/8a/KVw1JU0jkJA2tER5KSayifdwgt1pSACwtq39rg
tez4aasyTqDYBhsSeIHhU5VkaoAsnr43eIR5chZ00dg86PATzT/RxOn231PUWh4MZK78h/qhXxOX
xdbgEv+sJguKSHqy15JySPwIqACaDisBL66mF1DJ9QKrk4tlFFhPYR2O/7jSDO0/dY/xP+XCyo51
GkdDDYPma/50tPfg1rXEq0jnw3nmrYzebjRbLTi0j2+7qcnjPRm9EvCosUOJ7buFwxH0TdQweKFr
kcX3rhoAAKk/4uf4B96mltuQBUfwnYs3AEELfhzROd0cobzWsYBLy57giA4vPGiTvASBbdu3IuVd
B6zX+TS89LsReA3hyX3b0qHLneEAtH72e15gLXctqRNA1H82OyKDkdsJxNyYWUDifCXl2L2imB2X
TPwAoEvZJ7W5NuoDRCmN/z3xfLSr/6V78TDk8xzmFa+L4CPUwoRhFsYnBEk+soPBLMmZDbM9+J3W
z9JDCizzTvPORsjid46Esfe19wwloqBbbphPS51VPA2RCkYaBR62WpzQdV1ncOhhBZEwfBn7J0Ph
CU5+X8f6lBie5gRhhln1bdmi4lBeY/yLURXtyiO+mge0FLZDDZ0q2UtatERcS1tg1cZh4pGIoqy6
ZONRRX4cmSFhFWKmxHm7ofXr2M+6uDxyc1J2xaoZUeVvRsVfKIXNfszCG5S0zef7W1TkPiu6yTbk
t1Cwua6c5NaqwRo3+b1KrLRSGc8oY9rFSnMPQma+8S5JzcqQlxvoAd5vGgSZkaNFOrGpMpOlqn3T
VdrNMtyg8+z8fvR494gxp7i3a9DxgD2hki1rTWRyjbtwW+NbAnv75mjSck/uImbGq3tz1r4+pSiY
6BfhgVSg7zEybmIssGl8a/hDwv3e9Y29qAD+vCd3ktHNsTKMqKLvz57sMaSLKdtcOBk0mBw9WGgh
iMSeXeL7Qpx4Br3llOc8bxNvvYmTmAgsbQxYjVs3C83eRXsWZvNKUWEuuBWHvzRhk2Tsqo2CQlRq
PH/N5yXauo+le/lAzQW5iK4Yfrmxmo3RgUhQPVRDQwPTabU9MwDKnKNCheX6H9ps+4+tKCvtzazb
uEhyxBC3pyvvtoGbrZY2/taueP/FhCtk59qrVrZOKD+iPtAPbD0PwJruDvh/bGz595YrD7OW7wUK
m9w5hNA7o4nY8BK5MkNH30k30kGzqTUd6i5NZgl+07lZQsqLPyztH6CIxJBc/yuusnDEWmZzMX6T
03LttVGrxjA2xAj+lTxkUc5P7HO1oMln4UHR4xUt/epL1fImpDWgg4J7spila0MUsaUUgT35w0t/
ReTUJkKdxFfhVBtVPKhxTTFSo29KtRtEvtC0hEj5jkESHMotVArHz0euey/jKYOF8hCpR/YrKHq1
LYI5X1EIaOy9jp7v7K1PZW3i1Tywu9RsOMLSM9Nfr/w80yRA3aFwNctK6Zn/EtnxsRTpw423UwdK
DOWyVmBbuvri+MlTgdRcBnYusac7ewMvChbTU76BAyt+GFPcY3iG/D2pw6lAGmwwRuaeYhOts4g1
gkEsBbjSCtrcO9ALbRWsLUN6AZFEHKudFucixsMZmFPSl6OPupbNy4xvWK8BuOFFwMbUPK1z5c4r
XpYqR/ixBZeQ43Q1h9N7hmh+GqtYgRAl7TVI0M9mZAPFS46eJ7zCi+g2mNgD8LxXwYjWl1qKmSc2
TUdOimM3uACw39ENVXGjbgSFdkxdH56Pkn/vEjOBkn39Gp4f/3VQP9gw1iSSooDUwr2sgMyxqkfl
Tm2Vo1TGnU4W2La7FE5Ufu7YfaaQm8151/rzjUPUssqYGfI9uhW9anFUND96/FOZ9cX8K6E0yB0k
f+mqz4GaVoAEZdwisu2Auh1RDZFRaQWVtQER00gz3jjPIcM6cutdfKvkALWZzfqHgn39kTIfPdx0
UqpFiOO9P9Yr70eQyyxQRmvBiiJluSDr4LWrWR68rAB/IuQhxNHMpH/JYXPcook23J6iUJvKslVX
WXi1uHvdb6liDeR27vZdAVatzQxS3C4BohTV+52MU67naPGebM9/fVY6gDE0QNPfNKBQomlEn746
nY7qmlrdU5myv/xkDuhcx6Yxq2QeDUnsUJHVtCjKbaA9vHd75r/tkubfu+GmDB4Rg+apeeEwjDNb
WRLQ6skfCAHBSMwmijkL1/8Mt/T9pQZ5bdsy0ohXMo1K9s9fVMDh2ZYyPZFaZVBGGa5SYwqQ0RTY
LmN5pZE7YtZ8dtt4t64xM6j0cCcIEaykr26ae6LM1q8enQChvrzdHa6ABlaL7TFpVpYw9erwmT/0
BORJhNvQg150yetBYjCDN6rSN2IKUS8QYl91fP+ygJC9bTbn+Nr74FSSmMIPCsLJZmH9kwTTXZTc
pL4gZTWznuCNELWc7Y53RANcG9uPUJDRe9i0xqKxSRucN2EMn6KhfQ52TWdbsqzhJR6BkOSeT9YG
Ht/bAmwvCCBCgYXQU/cERFVE4aqkOAcWm6qw0BUlyXKvW+s37sO4dRPa2ly3NxTVRlqn0nCJdoas
lSaHK+NrXEAsd4GBg8hNxvDfqucPCcDNwSzJfx9Wo5zqnV8i4IkA7qPxlLOrdiJtY71ealmHiDe2
EUb35ATw+sSuK1qCRq2e+IK2636/bnkrvY9/Xc5nDMkNLgLz/+28DooWukhTzKkcV5vCvLgQB6Vg
rG922O/C+bIEUKjxCWS5Bo19PRXuUARq8kq+HvJR2QiQJHI5Dbb0Bh2RPmHaC/uJ0CzGwWuuINNF
kSIcCl4fJyIyY/fZfWk8gBQqzrd/shR27TJutHtskwKy2umF2jULafmkZc45HiZtCMw6kvvoCE0a
2SPJYpesbm4oVMDxGa1Vj4x1h4g9gsF0/xYJQCVNe+BFtH64ZCIa2TOLkfkG7kbre/SPDctTa3BE
gBXfmITwUAi8Izn9LylDAw43VuPahmTrp/vecX9vJ0xmH5+x197Q06/hUuM7r6Fxxf+qj0+gIJnO
9i/fpx4Vg5XXZU7Bet+cqSE9EYYl1yjSzAUQ9eBXkc3JCfG64xWy9zyUZW6HmYePDCUiGsHtrpBH
WoFrsUumu8PhJxQPpGnz2lxUg7W2ei91wqF6kx2FiJiKWz23NMjQKWkHFo6m84NrC784B5spxfAL
EIHW6WcerafwVnOe+eF53OZvPMeQavwj2urzAasflOigXbTeG1YrJnBekei1ssaoWzj0qPoSypDu
UpOsak0hylgiCx526JYVuvvj+YbF1qNWTsrFiDhcD53s2GDta+N8IKoKtSw5F2jJJEw6wu7BYBjR
hZnjRgNdyX9EYRZTue/jZdbttOEoH9eLqVFweaw9CwHaxvYi7TVvFB5AetqIo1o8CKWgn+AhNpE2
oiigiE30ny/uWGUxI07BPgFe4MCNDMbaWVDWa5hAurXICSnbUUzFYKKlcXTCqODCkkVtwI3Mq2On
0rY9Ed+6lTq9EgxhzA9bRttFdFitZ9zu9pxtCr4AbUiULtVgrOg3ljVyqtxQAEJhN3NBpCSUqODP
3fjHZceRT+StxBXWwsA2dY7dpsipIxprfeB1/KzmJ/g5O6CwFp6ediudR3nCCcko8f9uxKpgnXCL
u59+q12iT51iyEW0JJDZRGQHlwCpg1DbTk97B4HNW6AcSO2XBhV4Xs4uujQWBAztEnEKRdLEELqH
1LYyAOWhFtIUvX6paTomVzM8QpTWe7QZ8JSnlX0huk9mRarS6vrC+woFeGKn6w1Mm428TXddgHjx
EE4xDzAp4c/jLaCG/PkmXLE0f/uvCSQSVBXzLVeJu5CVkZ0z3NPhgbl10UhVYhCTMUaKbgEgBEEP
LQ2RWVcpO264W6b+LZFf5UJ806SCJ1w3MwvkUC7FsVz6oNm+DOF4Tm/Y5kGv1MVijNMlrxFrb5t4
/xsBIrbD67UJyN8egRT0Zm88E+ttJWVuMBsfe6h3f/FuGEL2WhcnzpgOEQfRJ6IrqxMUrvolGnZh
Jv6wjcIm0N9ku8BBhB2NwUDfsRqDdadtDl8GQWyW7fPg037M4ex6n4hDmzaW1L84DtDSO05Ney61
PdYXg/UvTGoVm925NrjBQmsvMSR4Y/AbBomd5oLuPMyf5yTstQrHw7FFEXJqRzD989UDW4cZzDtB
fpuwLz7K82k+kzg5BVCWxp4Xcho+ESZC7u2hNoZIFTwGfDSJodjbfmcxkM3Q0+QbmJyMj6aI/kLD
Ogc8CSauABBemUsxg4YqFPqo90CjLu5YNstourhDjg/txkt+GQv2ZueDzc6/GgT8wPvjuaGrYpy8
qs0C9rihZABGlXBMyXnoBBSVt+ZtodrFIobFRs7nZlNJgtHqcpQOSzbDYPoIAV5X6dqFaL/ihLr4
Zz76eR0m7S85i85KEOkbtVK1DX1ysVxGpMLLBqv0ntyvSooJRXEt9L4PDTVdIYXJtyc8OxWxLLzY
ZGH8I6EmvxKfl3otqlbph81fFBYls+OX9O8fznckE6JKYnI2w/hw7l72H5OVCO2vI40SXohgde2o
hoe1REfDo0N4q7fPxJz/kUmzOsPuh9tMqgBXmsyFndoQIKvxWWAfNATQh7ZYU+Jx9yBcHFKzVu0l
fuQzWRvO+Lg1GISjLo8UbigfMYmVpztc/qKbq2pGQWUs46uYJPUVSbvXoAtWihFnY6Kub87mf86S
kmYXVNJYDMt7WGss2rjA8SoYZKw25XQKwHPA8rVwMJzbTlyzFK25mDVXlWKMDm68h44vUY+yVNcU
5cdRdzu1zXruq+udRM/3qWi4VkHX+3iEUPuerCuC8VRJA8ecgQZ0SZWy4PXKICxFiFhbCFtqHTJu
YdCs0QhPgnhR9Op4cy84osha8z+XPqf3FDF5e5PArF4tR7t1aATDOC91lBVDix8m9MeWhbcPC6kU
Sw5L9m57QDEJjN1TorSCt/8Ql7T3jqYoHVzoshAj1B7bIguglzYDo7NqLk1vXCRbT82S0dUmZE55
o9lyxPh0/wwJMgb3MqySoPsDRCHrj+eNP30AJQmXNNioo2OCrhJ/2YDz4NTzNnEi3jJEjBdNweKs
USBrLsoN4SvaVkhBVjTXActgJdtqdpQoNCzHK5HYNlIIPuG9tdkl1BW1JChDiyT9SA73q56zOE1T
PWaK9CTI9uF+NbSR1JbYPFPligSs0Tmo2ABdgPCm6mzxpO2809YkGQp/XG6L4+o+S1JYUSmEBck0
u6d/ExAo1QL38ZD0mXh45/wHnRRBAxHWrcsrWf92EaYr6QQKiZCAdpNrr5xlhySDp+GUx7N+2YBl
fS5N1nsOe1Rg31kpyHiMqsFpnR6aXxB9FCF4W0mwnGROelf18RBjOlEVgKg8yBwMVTzP0gI63O+O
aMfn9tBlQcP2iDolSone6YJTMAcNOeixo3klLd/o2L9fH0uXy8t0BSjSiXR7D/aUWCW3QyDsCzcM
b1NfGM7GeguR2lNngSZHUiGtebpI0vr7MWQ9VUaEslsc9l2VI+ZSANfJvlYNwl9paBGTgQNKO6Sw
CLDU/teIZpSS09TR0c1LeCAqQGjLHLli9F1RgSGLPFIEe90azqCnZTjOZZZL1BPAOIhj/ZihAOOF
4fCDet4abqhCWDw8tgx2kbW37pnco9g5c83DolNFjjFPr2jxEhtiH+0YRP5EEUQXT+Uz3izPsIAB
Be62qVXBlbNoXBaUXYIQkkcNJRiHFZeQpvbrxPEgJq3GTbx/VxSWdmc7jx6hF19+I+ttiQAVYSXP
zEKxirLB4N1Lco73HnNyA3av0bn3cSPj/u+4Swe9k4GI4ZV3gjJwxWBik6oo2Fkp4F15VZUdsB5e
zNz209hoV/+zalCeH2EbDJnedoJIs+nspxa/d9ZhJUgMMPT7/kXeW4nDqyFdGjwKGxCnqyznABZr
xvgn/lUx0tLVVCdsMFQfGyf7C8gdpsHKxWd4W2j3DUPLLhbrpTytXmH7FFjrgBC70/kGunrtqxwC
fMzzjknSNZp0fibxDMio/s8EK2kB5h6et+kQzABKOqafxPY0XwwMHEEFcFTtgUQzDSHduu9tfTNN
W224+zmDVDEOElYW6Wta+GvCsFakun/WSPyoNJXVYuVeK5Sr+KL5XdN0D8h0v88fY3VkHKp9PEt5
a4dftQN4O6LV3OforzTf8SQceG8hHbPnV+EtFcBencxbEVNiT+St1SwboI54bTYRgs6Dn/QSr0mH
+czxNBa/02uMX4rXI9Mdv7j6NvfkiIQUkQPLRqK04YDnv7OWvKP6lkkS8pCGzf8FxsIFVDmD354U
dgC9vPz9qhXGsuMvltK1QClhWFiNlMYkaNINupQJlF0tLtZmM2vHhRJ6N0Sc+oK4uknod3jvE9fJ
YFSwKe4i0zyNKlPz9hqlpk76r2vMXTZGpA10uM9ii/kqc8YRDO1eQGXzLZeuh+9T05WWHCLd+M3S
6fpIA8anT9gNr4lWvb7hZwWkfJ92k5EtVygwxmO3t0D+O4aax/GQQYsyT7IDweLqrXmjbwT5C3Fi
YIDSe1mUD4od5tj5NkzEaBT8yD+9xU/Y7bGzsHzu6669X2GPvnLxy6raO67TJmFjQVmATeslOkCB
OTPPMw7WBHa3bTHi09BQ9I3HFYTIWh+TfTmy8FeA5hpl5J6GLxYjCriCcaL5gxnB9RX2+6wazP04
wIQOIk2n0EZgjLtdAiYrHVBpmUWO1TLrhhubNxX15K1GtJrExma+yb2E/zYiSvBVW3/A3zlNqUym
P4Vyw0Yoy3RDwKofRxO6p6xy9XTxzFGvRxRAcS8vaqO2VhIeuP/B75/8p5JGaB3p9Y/ICsvkqe6G
FbDgKXd5e9/Wr6CwVKUAbdCa942ZZfrwzGgeTyRscpPi8rXjuUcQFCCo/zwveVEZl6tpNEywZFxQ
t+dI7KWGYtQMcgVZB+qhfIVgxoL1zpS4iI12LDaUz0yiPMi1vbkqGqY3Ofx2nNIo+de4NR0+HWe+
YoKdRfEG2Ob1aHaBM6pjxp4gWE3S4YxNbskLihS4NwFipI29CPVjSmbBw6yxkumPi5hDwVq44e21
kBrlTyC+0qAzykv9LU6J2mmtuBaPAC09yNCUo0/nw2nlvl6aQoCgXGaH87V0KuNgnxwv0CS/G3xk
HB9YJGRbBy52dWtWwceKcj8pLZO9QtnotLAG3KCeUTGFDiEu66bd1qMoAPqRvrDGbo3jGFf+TpGq
uVUi6+JDTguHcYBn78WLERd2zP9rV664EL9s2hJLGuAmRyOvopGi49P3v+h/udM4/tKWC9KeSfR0
WQs7b6Ybltu5LwSzQRfa6iOx++yGD+R6LQ0zoXovvPcH3OuTeR9IVuvpiKaNs7vKtISzLdLg84Xw
LTqOq9pvTTjNySAmlD2BCXnz6swVFK1yo3or7GO7j/WyP/JyOZYnILmmU1RVO37TEBNqMbLf1L/+
SOpH/CgiFoglsxY+QoY5/J9uVTELM2AagVzfgfM4gWrzg0BppYhFeRFKf7GEaj61tCLmgfEhZGid
KVy9b4ikGIiGcCfvpdcAIldjoKpZPqDDee47Y3ytKE/1SjMHSk9UmB/s3Hyb5uzuWERSL+2zM3HX
ze4v5WOJF6gUqk5h7bvjAWYeQrK8uiwtr1ziZr0XKMV5/M6ZY4dIeY5sNpr9iWLfB1gEGF6lKRdN
nYQUlOg4AOORc1HWBZNS8mprAQDFD+2tl6EsMonX7HGsrmSPcokzVgvqX9igjjbK8+jW8pBDeYzL
uVGP6bJLRLNWoKld0pkRHDOirIm50/XJdEFh/m8Ri1nQmdTEAdC/ZiA4tHapLpFOYhrhdJLYjM9D
ltEgJ03LP4gzThDmfWLdrqx00IbGIQdmUgfaVO81FJWavB1x5CQ9AdG+wEba1eZWaX9cuhC26eCV
TJXqwlPylhpZBNpRb0iU+aG5OoxnOaEZzd2FHDBHyfoFV64c4VoMW6H678hDE0KRAt1xcE5d3cC5
eL3YI524ggrjOR9xW4QgnR1BXE+Nymbj1bRIi1BBBogJ6s6SvsT+sQ5iItuAFJYS9c9Bdz5eQ99h
YZti7LJjiOWjNiiM09+bCYBF0OFTHVjFYtmdDtqA3vlDEf9gs/dcAFt5Xp9I2L80Z+mxeCS/3ymn
N25GjyONitqATSPFiSKbIHo8KXAFlD8zCSC6Z1iLZmvZrNFVvyj5Qf4QyboX7mOqe26IUueWnVWC
ws2wp249nxQ67vOT5wxY6dimPmDXnSc2EP0Czy/FHYVDM3YWKb0p/0iJCnGCb36a00aTAGChUpmj
JKvEwcMUuL2aISeO6KNtJaDqC7u0CJ+6YUc3CraVDy3e6X+lLTcssPric1C2t34o4oB7vdyrNdJX
5OG9+tSFeV1zbbLTu9TEiVLfs0i7RkFL5CrnzmWBoUzVWCwcEsVRW+DAYe3CB/+9dHmbyvGp2ctK
IKPWYywnMX158XXb0TFs4E9PvSU9HrUSk1nJ+E/xsztw444fVqC6Djcav73hJ1ogNq+251IflFGm
KfZPRa+LFhzXDU/B0Srrk9t4hHW5wcsP/KytN8wF2qE7Zwv4N87hEAhoR5mITdi/8C2z3JGakPwF
acG0Z4Si6bmyDgieZsGQtwxTtZPwRDw0wIOzGIe4ZnjR1M0BJfOcPDX+UUEOzybDBtvt5LknciMi
1MJPGlv4yAYHnkiy80jnWBNdyGvwVmnFBEK3M456draZE+EMLSS0r3tVMQJrcOsgU648F9K2bKpi
o2fD0BDWp/ujVghHmHOahnVPWvSzThiJKrHWLb8KwoEnb18eHZyEnITnM9ZKyKrVF/EFGps6VTUJ
m9yMs6tVosB7KB8K31rKYL4Pl3ra9XP/sT53uLIp3EZf5vmywJGzMNYIobZji8rUVf89hbHkW73j
5ivTgZjA0BCoMPtNTuiBwnywbkojsbS0Rs7w3PhD0USoIHTS2aq8Dm7D43w7t2+ySN1DAgo14UvZ
nJGTcCMdQ6nBx/4v/pFOeZd4No4b2uyP7xd9rFivkLSlucQcEmbqeS5hqO+9ejlQ5JgtPZ9PXj7k
vgaAu2kYV6PVu+Tg3Z43cEQegGOTGGyj+caezFEMKhqqTThJT6EyQLwROoIqmWjT+pIj4KiDYLxO
dQHTahyI8nfaok5KV1vEQE2CcEDLdm/3ljj7tgL9Npdx3pXOQ++I+b6zTVbc0vXovugCpaaAZgoT
VmXhebativiVcObROu+/M7OaDMbkWYKkaq1q00XyWVjiH/7HyeYKQprGuY4Ea9FyaF8QaS9To9fK
UDl2G6mEVotTCpWR+0Wx0FIv7moNRBMlz561hXBPqr/+4Kr05hf7TB7A2jOOcW7f7jST4Xq2BHpS
QYeDidZTgd6PIjZVar9eAKZOijaPZTSW+wFTSMf7xFLMlmTUEz1BHx5C5hWaTomt9l6fsJUE5dL8
g4/52+4fQa5dKfv4pq7YbcsQ5zYIZh+jCmFY7KotBO88RjisCx/Ch46V1Hz9QSqOwSHingZaKT8N
huXcmEEDAD2eYBZOCxh09r7b0uBde5IlGqzHfdr2HE5JuQmxo+Y/Fh0aPo+2dtyU1miNGWv8yGVi
oZCmn7o4xT13/G/GrJVIx3yCjdj/TuJZfR//UhrR20X7T8KbmdkiNKaR/LeAqA8pZL+/TnD0oB9W
yc6qccgKDY5tCvM6uQd7MiRBbAmsP8Ytawg8zmZbW+Ha0T+d971S3y+IclzZfUGxFSBABk7JQ94P
UFZfdsnlGTckmZSnfXPL7LKoT6ub7bap9sV6FshcgwBiVC3zod51e5O0mpBfVi6X/mcnET0m0rfY
ZgSAixnSoFN/Nkvp6dvjIpXa2iWwIBclpES1j3I0OBfNp+ZwYNspF1oJMJdoeJfMD65cCYzt//N8
gItm6nCnf8ad6aWup0dptWBWdO4jtTWyHEpGhh2xRyyr0V2tj7EBR7xiTSixVamdvve+RhpV6ZG8
cNEPEQAd0qi/xjhAnKuIVOsvuVIXfydrq9/GcFaOfKiH3Tj9qDMIjqgf/vOJfomAWB/IEHvR8evF
7AWksK78e7ie/M86BUx8B+KpJPihXRS/tlSV3YuJFjHZiIprDiy8QfaPK46T6gu1PutHLXCLP+36
dbNPrgKno4mdS0gttFrtTScmEHwZlwrksTYo2lXdzbeQ1JoTHcY/EMHUlvdRvqrJGvCmzH8iW8eH
qii0jbwqZ2jnfSyyxLpkZUQ5cx8dH2iSvHAvR6lGfPitm3VqoC4OI2iKxmnRH1Mu0uREa2C3BIdV
Aq89dF09T20PSdIMTE03g0awsEmsH2F6L87+DFjY0zm9jvZBOn8mjX+/nRo1wi8wT1L4RqMLDfsZ
pSVQ3afRHzYLl3by3bYDZqUHrIoYpKg981vIJTNXjE6GQ3Wkgc1C1ml/q85lpoLXdQcl+RxnXi5W
H0Xvu0FN7nB3CGK+po66Ljv4On66TEQMkxRA9Cfmll7JRSOw6R+OZ+lJ7A55RHswGFNRaA/ywbpe
t1dzMs504/F5Cp5WH1FzafVeebjxmDZI+P+ghW/uUAicK2ruWVxiCesjCR//wgRl4bU3p49h7ug1
fPC09kdxxVIsIiDKsRuFnJJEtQy0Sm2OsvHXBgom/Vap+4Z3q0MDySlnTzeOlq4L1MqKzoTaKqMb
btSCeJv5CP1LCGYbT0mGcmruNYGb3U1Qc/znk/LlhY/w59HK02o6dJadQmBycpTwjYY4+n7kU7el
taK963Ws2ZS5kPaA+Apjo/gKPIxJ3bC/qfQxV/Q1etxV9yYDuA4xYt6d2fkX4u0ZN6nU/+J9vvDv
hUYx6XokrXwhSG0Kis5mSSGwNImRGcRY9jRwZ/8BFYFS1KGqVK6lSIs/3d9+4ZQ3b9mIhKgnsQIv
bwtKiYg5jbekjlpnR/twvVfOiwrelDEwp5jrvtamdiq4H1aeQIqxR+liSWe0iF8+iEBtSboUcK7E
2B6gZ2xS41MHmuT4g3PUQpZRUmnEGW4+bdhaaAPwBxHed4lT1tNsJS+Psj8o2x/uwlDxXIPkGWIQ
Z2gTIoati5+6ep+XJZ2BC3vvqopd+POxh0s+8yLd9Dgbj8Skg8cooTmyRK/l6u0RfJqe2Q1to6wO
wPdLuUq9TN/GPjR/GZ0e01PrIMd8dYXEcfv9mO4gRQOksawWFQQ5UQcc2UXpcOHlhX0+z2OCVXSP
6BOJjLVhovKxRRkhLpVgkZMEUTWMpE+d1UXeJZaqq+mU80i2Pg0YUo5fQieOo28ExJQMiiVb+SUQ
lPbHLeTRYhtP+Q88O1qCKbX9aFNzRu5DGGb/Hm7rSgWNAIUIGAzqX0PLsWa2+YtjdW9o6lFoxr9J
PdniOZJ4aPnl12RHP8N9p6eF2pXVCbEFjmP8leH+tKREfdqkg2IzYS+hxVnIXfUiF9jhUM/klLdA
G0Gn3wljD8Q2Ryz39ElfyiKSKPrkH1eND7vpyMV71YNU9yvuRNPrPSy8BNwHbr036doSQe2tv5IK
oJqVRnzVbzREtIghXKUvGhVRyD0oXNX5/aL6GbeJTyTOGggFms301RJrkOo8Q7zusDCc0Ze2xJkE
gKQ7Y1lu9EWFSKQrKHPIAV8zUDUAg6OPx8bsLMPqvFePk9EfM6lzv8rB+dDdCgg4A4Wa6oCYDFIF
EPnLlbzwcOSDOXXIzBpNQNrlxmS1gA0+PqO9CWlTUuyQNQIznelTsBUD33VBDa83QdawB7qKDyQ/
eJUQGhaEkRasErdC7JeVABDi/ifGSt5N0VEAT/YyTVA3TkHykRhx/KX3xvYoG5qNA10JwZDGgEzP
ySHO9LfqMs6GOVR2bPkE7ZVSQjog/ocx1mPDTikLkjyStf96DZeKamBFfPTHuy2mDUFpYQlcs0hm
Guc/dfT2nIF1iuP5tMAr2dGvECXl2NdIO6QoZsQuAKm5BOMQf5GWio9w/6DupTqFBfadeg8NkgaP
W7GykG2+JdbFO01Sj0oSY7s/JF2cFjHghGOKbaOGivMlalmftJFJgSKv7Ir1gURcJGM/0IGtG+X6
pvGgdqVpfbQeGt/luTriZMvw8TnCdRCAAOiOL+KYfuvnCZSluWAE2mHa6yy72lFFP3tlKAwUYCzJ
USGRz3+kwcOZXytoVKd0fPDfE2P8ST2RpAekCVDKOs+3D+MJkONB0A57rJ1q1IkwO2JYa0IXHZYC
gT+w2gZVNjPO39p8NcSHqrDW+1Z82mNZFw3uUgk6OEH71+CilgyRu64swkRub2pr0u1hLdhOf9So
b4DGgd0Oh82vj93blRv2Yd1oM3PBlpwTogNbq1neBEtvls9FS7IGeNRxZuNa7fLWP4YscMlsyB5C
jzAyDpDRC3dhd33NLYg6Rfy2Acs5VelniDSybtsj/nazx1C5cTLFky0LvjNHxGSy3k95p0Boybrr
bRcWaJLn9E2OjaFwdqV4kIRKSK7grkkIMhTHBGUX7FSuPEo/rqGjCm5TxIc2F1D5cvU1ApTTFsM7
vNjtlUeCkoiDCewvyYMffYakyVXrUZBhA6YR6ajb/tDQh/kGb5E1u/xXe+IqvQvVJ6N4nuY8ysYF
bKZeHBREDz+70avaGhvJFNQP3Ihzy4xDCLnfX+p76a/S3H7p+MES0lO3IhhKZifG7yi/87q9Wghe
wx2Lo7CWjBnpHSqjMQ0yImhuN+TaC8tng0UASApe/Q8Awt9rh9Sg700Yk+mAgMcalMVrOqO9fnk9
EKeupxz2V4r5jLR+RnK/fhWp/UwOzfdMtZlOtw6cGYUP9AJsw3DuZsuHJHhkRCXFdYW+Y87uDT4N
WZvawmRmZGePzUcLNkbiQfH0YGszdPJxyafMUerVNWj0rnBop5zLoYjts4rWY8cqSSFz04nWohOv
I95O+Gtytbsq92jilycz/CDdu1zntx3kal2YcQE6wBoztVz/laQxxNOWeaiLLN9lJoFHQOd7k39M
B2UvC0SwJa5mZzTzQifXELrZR1q98ntUp4FsaYJGtt8yKW9u/FxNYkIypJmG6IxmZyeBXLUTJ5SR
cSVoh7TFugz64Q7Tw5ZLsQjMv21ohN4yQzuTqsa8GwayJv1WXXPxKQmDqxxhOdP8QROj9yjUQ8UK
Tvr63hHrgOMoD7MpS7qb+LgTcQh+EbImED8KMEx8bH9Glu/Upx7NCGy3NgMG12ta+yDre9ltSNQ5
Rnh/Fvn8qtHflhSlwxLKDeGGmYyouivz0kFSf+QEzpV+w0WHYVzzgzQkZfXphjL84n3alo3P6T8G
toch85cUsEf8r0OMw3fjMHVxAUD5ZJ6l+UCp9rHi346/2b1LwZ/Xg3F6STKxr61ccnPSJoxeBQNv
9dRmA6yg7vU3sZlKZyNsTy3q00+7Nwgp9RPYGmZqhXv0G1vfKY7b66Ul8ZXsU3MqzmuCuMeCbuFs
vKip4Tpo3R+qFBgHzJW/2CDFh9MPCf7ziK32y92OpKgakIAPvoZs1tLtIJqZD70BK0O6EvtYPBDZ
7rbyU92js4UfL9mjIOZiw6NWaR6qlMBNMIjajmtlaehjS1Pm7oRdRArpio93Q3GrpmjZy7yEWoyF
LiriCBYpb8a9KTnHtnEHr+SLsJCDQ3Qri3gFou1MFdrSfSivkkTHYVGNuEtReIFP/yDDcq0vuVNy
cdiVWYXtTDyMuKoG1+HdNCqQ1E0GeG+K3jRambRHaJYuUQhd2Pl+MMMF5w2nkJ5HT4pozBmdylZ2
L9oomwkJqer+7st+haVcWSs2NYFaFi2eS5pwIEFbC71s8hV0xp9lrdmabDQRvr9OJ9kzVkPoefKQ
YxhgXUZ/HMHKmndatoFi64gIrkcCVUfypVdNNx4iH/tAoyoL3wH6brlWIORwSQJNwkPNi5JU4a5N
yhJNhkXWMVHRXitAtU71ukNHISurWPGk0uzv5p1YVtbmIRrFxWIyHLIZXdHrjcZ5LpwoOQOaZ8+A
xj3uvM0dyxDY+q7myhlmDBVfStJTXmqXB/J1UQ0f4sASiYssXJh1q/IrbwGiyff+6JlK49AF4a+y
ppcjsAJcBKLgzZQ1Ky2JfpOneLK+xpvVJQSLQgUBcr6L8097olHpzQoQA3R/yAp+Zl+Ofd81nbci
3jXUeIL/4HI9CO8/efSkouSG9qFh/jb172pwbNHWe4cvUIVL4kQ5YpuWzP3l85XBobuWkC0fqBrl
jmpzpbfanpwcAHYf5KzNAJj+45oom9wew3qcdIO9FHYLPdlDu2cgdaVIr3cAWyUCpdBKFqRlK1J/
4JV9X8qcv8CPqGKGm0U9v5T28srrAsc8qw+dYdsXqqtrWtjjz2UsKobpQA8tBYpmEUDqSI8/5/zm
rK8gbpVTE/t+8TH+JElXgJKsE9NRaUVigFitgMy3v8bSJml5sGmO2yI0BfF1vX3SlRn/JYSHsjmA
602QNXg5wI3UPXMabFq7IhPB5jbVgJcJb7F69RmtVhGscQjsZAPz4i/3VtYn3pF3cwft1BmO6QJ5
XMNvQCkEh+N6U64ykEjaY1QF5wG5wdFh/t5sToJ11MEle9iYv6ZGM/5BfhYoXfPVRLthKAejM0oJ
7Art2oxUa9QDS6Muda2lbVFZQkmtPr/pNUrzxFgnVbkWf+Vs0l5XHj29QE6xEWN0SlyL5Q8EmbUk
0S4iv7jlwr/7faCUuyzILSGWd4Ou4pVlQNxtfqA+Yk4G1wnAl8Ss4qgeoNBHScboqHvtHmqR+XFg
GPLCJb95Yxk3bne9aR68scvBDZ2cmo0FxBJoajyGnn7NwrdSqG3WkN/1JcBCkdFl1JdBErjoWa9C
L2+gPIeT2iQKmW1grhPF4Mf9ibtosuubHymFThgsOHrkU5xCEjcjMvl1jS7ls1FXmBkrzeG2fAdb
r/i41Es25I3HWcSmBEaSFUcmgjtvWahUTBW9xorx82PrhPEr+iYh/s8cE1Fj9q6Zj5pjO43SMtr2
cZW2lEyTMEKFhc35ihQnCqhvrLXBIcJ5q/aZh4NTczuWmmcc6YfzFJUBh686/fO/fCspsUkPSAWK
Pw6QNXf0HktRaDknzZeBQDNsOpmk8eT+Qu29Aavh6XMRDRM6NA7WlgBg3Eac49BtCEDzhn/vgVI/
PlM76oTAoU0Ou4yw1YNbgz15Fw9LH4stBASkUnZ6YA8tOpbOXO17nUjdJXO4NYV1X985LCtn2A1T
bYhxpmRAB9+UspOUYXm0eGD67b1IcoNUNYeMGEnzNiVoBKx1KUkfX1EKPBPZCgXPSXYH3t1cs2lc
TKs8MAx7AzOxA8+Tb9w28IzZflrBrOKwzU+kLvo3BV4UK/yl5kQeemL0zpahva86fXReq+GPg3S+
xPF1Qszj70uDwQ9RyTOgPSIvfMzTGE660nWyZJ/FzlJiDWDa8mpWc6S9qqCkVsV8T0tzfF7SpCBC
3sHAXGi/Zv2SC6ZGNNK3sODmAD3bWhEiz04oMQoIebdDSpS5B6QTMSTTybTSSc0c0oKhDTMtIiUj
eSxTeglR8IPZ03ONkW1EPdz55nj/6KP1mq+vdqDJM4iuiQNUizdvjN3b6lcSwfWHyGkYdyudacb8
0s7oavt9g0FKEAA7lftjjpAf6pTE25SvmiUigF9sq1UrSdQiuDheJjOgzyDPTvobU2OkdiR9GShz
Rk1Q0y943+vSoB4HGbvmSV9QhGyUKMIpDxW/94kT31ZfPJisAkT0qOFj33YtTcu4cHDApp6DXoFT
YXIqyoIOVdgsla53BsnAs6OUhTHsAxZdVFqTIOLiPII+CasEqESHmssotVZOqufgWMchEv/UYWma
291CpeaWDG6TplnSDHxWrTq94EBjSJFZa2Pqp+bzmGZaCx9UPgmKybYS0a6Z8kotN/PvSZfaaK5c
98afKsHii67PoPW16czyd8VDJKZqpvRiqVZ1tCFWPyBDaPokKC3jmnwJbXAtpdncSLI8VH3Lss3L
Eew6wX/Kfea3hJgYL1RRSswjqxc9/ALquAEXyiCaLh+HzIzdPkO9y/afzEd1PlyIjjgbi2hop7NE
cqXVy14jB3DRFe3NadxzckRWtEREd2587yQdNVtj7RAdqcAO4ASkBF5mF37uTI8C4ZyYjKoKu+6q
qj1VGoq8lPwgiATMPdRC5R+SDn4NgOSExpAgpb3mQ9L7WeZD+sanI5/onM9h1UM5ZOFkz8XnItvf
oApKNRZ5w7OMqLocOFCC4ELL8lCDwXcc0PZruN35kQhJOPnmLfNoX7y+EV3UxbvJ5Tnag6XE7Qzz
/fEt4Y8wVlm6WXS3hGPEgw7gOPL1KM99rYTmqRqXMgADzm97Sv9Aj7hjLYWyWaNIbZw+VJNun3Bk
VC7p4/vjlTgYOg5ytuzp4VmaX0jxWdP1oSZvbDi3xv3b8HBEGoVMi9qfpBCgtGq4LezMsrRiuBBX
V+ul9VJkd+f8vLnEH6RMj4KHeMCv9RuDKr3cWtrwEWJNcjNWrz0VBvD5bUTLAh0XJXYpXeOpCuVj
Z3PHwqAy/0e4hv0TrRdH4VaPJfvzKIZ/g1sO75WHh9yvbUnb9iu44r2rhzUmDoNYeP6iPoaQOeSa
TQpo/dQdXhVeqchIJw68h7mGgwDNso+DdtwmYd5o6FYAwbmRAfxzAM1pgBvXJ7fK0l7nnqPbZ+Ek
UXOPfu6mV1AOnrq2lefetDwvoikaU4ftvAGZ0ff5EjxIx+TWXpAN3Ax3iMlBUXis2vDT9Utg3xHd
AlCkxNLpvHTAorAatpgPW6IntAdTSgKtciQuA1YAhT/kC2cTCboIFyAxEuh5ZV7eq1u7gw6FKpvU
o3gBN+7MYR1UnTPNO7gO6zH9B0VGU41eWVKzsux9S8aKfhuA6+ubP2fKxEVzrDsVzUHlaJ7OLkxt
CXo5Yw/iQMivo6O/8VusTD/PaEcFIdRGaHJJ7TwIY7eCFPDlQLEI5L1wsqTKftKc1TQXdMZGWKN3
LM+p8ijDiylLLO+T6ivfyW0xfQcmgHa8jc8YnXL3Ak1WrPjJShCwME/8NSaHtit6MIMacGrxGKSs
ZU9DQxe1ZkCGCpant+bv4Zt3zBRDo8K09f39SG2D6eti89DiF8NwB0RKByX6TBdcaoD4si5KHliX
gTT9eTh64fWpjFewpPoPes6pKA8TiaHsQTMVTLMwMbLhXNo1mw7zIMQIHllnos89Cv2fbJYj6q31
MqSqN31Ollzcm6Wr5rE6FOSyIRzey3q7FFPPyEeatCoPFRgQJ0KTtCGmfKxqohFrzCylGtc5IH3j
bp32cf0PdjBLiH7WJsbjYbLjSEKM4e++1WGgvf7y+IDkf3Qf46YsAWf8YCLVuXIiFHl7FKd2WTM2
jl8bfRsaQHzGFYSf1Slzc+AX+etLr/8f5KexfJLzj1H2whl3lQe/VpAfPyJnqA8vQ0Ev51oLbUFX
FtInKGLQ5x52rm+KKyYSJ4qwiquvJMhubEZl12kJFs14olU87JnNm8SPi980/P5EVsWx2YcPsMXd
FQ1jmJ4l3ahqePrWAlKOAgZQklrreRF8eieBt4AYViHRaYPzjyKk5kpwRtoCDAaocWAP1MCU5Bfj
kxF73qWiSzP+YFqTWsXJqARDIPMo3RsUnkIybSToYRE0g4slClYdUXxd7q1Nlgxr7Hzq1SCJZIdx
nUH4hh7jLALNp3Z7eVap4ireJyMcabKWc3nYpSTMVyip2MVHcVYTJGSWCw0RF159cQwbNBc9Wsdk
AWgoJs3QDR3s/6bq/8PHHzNT0SLqOkzyKRtgLz5dqhC8Sra1d/0LqVbtJsn4kysi8PlmYEJgXe4P
LsNAF9r23Ua38haqBTSf+BFERVc2Ed072k7HvHyPDErtMoPPG29i1Pi38BYQE/JeeYM7rYh/SOH9
XPB4LmgpSt2uZcGcMhv0c5OBVi52W4UbATKwnQvW6i0dChCjIhwqavIX7t6KvmwL1DI1nlBRYksW
xU5hEikdklD8Sf83feymTd+o+xsxmDmVoS7vc/0gO0Gp7thktULGC9xS61COZTIVfxWn14pLFoY1
e2tLJpsFKL9klU237CfAIFa9U5U+dhX9M/IFaAvigVWNo2itGi57fswXkw/TsCG2T+C5pldHs0Ra
5tj6Y535nsHN5hQL/sdZz1s5XWbasvLMv2hIiew1aXNyArqIjgxdvcCqI0W0tzdelG6IlsRTQ3R0
EP95R5nKf4noXP59NHgOxNqxYrf+EnaWO/iCEYZ2MxBOrmuG5BH2X1CWmYdZapDURW0UYW9haA3y
OXR+kFSmWPaBltKaDOGbvofmlHWQa2CS32kzHMMWxX/GZ1WxeUku6y0iZHyorm8cT4zfsDWJbHBv
YSUECmzICF9Bu7VqIoNuVc19WVxgQVy1G7iTAoY/BC+Oymi/MPhsRFOkgkj/CRyBjY+0/m+O1kl0
+nq1914A0bLE9GDiaI73+ASA8CYHalMAKZtKJPOBRfa4PgSaJ+pQLIQuiDZfy++I0NMLIbGpm/a7
Hdo/HBZbTaSnrrjAb6+fNOv1qju0jSeAAeIqNZkURlBtmcSUqw2S2iuu3M5Bfx71B5URgpVtHe0q
f3LVHGBxZzDyoRDAWEqSJX9d/eHSbuhlAmy6+mpprmPSuPMoZDPF3gz57AkwiV3v/QCdRHSSYVUK
I5JiWjMS4YNsBYOaYUjNmkyAId6dqkS8xjf4fYHxyMkO1TRDPrOQCF38zisctDjkZ7VFxaQ7RVx1
xRHyUmrrtZpLHpS6ra4wRCyO6XRdg3UuvZxlXDM27aZtk9gXcGIJONCyXEyCc/RnSepQWuHvodJK
CdguLf0GGD4QuG2TGSp5HFcCLvPGa0pU461Qs7s5CHdQ4McLK8NM9wJSLu3+48CIvumd0tCcWjgd
NLJiA9aS6h6ukG+Ckmpul+x4HaYjMgqPDXOIHWGNQUTZVX72dV2wWTNCmymPoNm/K3mjXZX3YKAs
8jctjUjhxFj/AqfkPT9tEIrC3PAEvydU6ZWhrAIIt0QU92xeM/FVrjlCCWesc8+nDsmCroXr+LXH
P1s1vgekzp+nno/qeq9YxhRCFr5MSjhwRR/w0dBOJO6u4mGEf9kN6OWKjpzxJGmJzIeMm61OMdOp
z4qMuRa9YtnF8NnI4gYwY5KdzJtadu4uG21Yjoi/7EG40Vw+yWqYDvfuyhnVTZh+titNA7zHM0qJ
ThiJ0/qKfAE8HT8zipAsKtrlCc/VgSJE3UdXKbEeP2CFo/7xaMj5MaCW0isW6MpL2mWqRu1LtjKV
mtTcDm6qMB+Nw/7MJNkm5WCZjTNijlMJk9/Ijn4s191s18FULhdc7Uw9K5TYfXp9s2LoWee0tzDW
ZxxoPdmNOQSrSeveiSVOicFBZBP2xY720xmIPBf0NDXL2LGyV5L9/UgfKCaINoTwY4p8qO+Z2BVk
YoROgM4on78fQEDg1dv/rOf3K8VfUXQOvtutkXj7oJPvCDSNRPYmf29kXiEEbkh7YliJQ8DdbBhm
5hNpA5V2KofqKxjXJhOwkz9lICujDdjP1c9SJEDZxRfouhvt52e2QxruzQCT1wOCDEiYhZdYL9xZ
jEmtUSkfN2QQ6/oucBk5R/sqCzU47wp3sNH/4emZiK8DJKQS9nbPSjTlR5rphpxj3RaVVnUfEdwM
8Q9ol/F+kd6l9GlMAG4nYnsWKqHTisBFUPOuhbZdjgrsrtD3VRtYix7vyg+bfsj4SmR7GTHUnApY
BLzGiZxFnFY+3z4WmVTW5CoSHBevwftbryMd/E1MfClyeZEEi9rIUPpDTda5yt5rlOgO6Km2FI1D
KCQRfOJ8EM6VN0fUDcloV1dTScmbgUHJ6HOqEDx8F64fA6CM3pVXx5iUuHvVLmSe286+Scae3dSN
HapeirCkpfYdyGyqNUC9tAZAQIbBbsEnEAf59HgIMqU32wp/z8UtPl7naUJ7fHu3oE5wQU+G9fEX
I9QR3KIkuAZ9NQ0c4Hg2xSHrfWx1yYwDJsM2xuGsXbqxqy3PJmqyoxA8Xz9rOxS8dnnFzXWGgsX4
NFXtySacro6n0+rF3oOLgqb+W8dNBu1F3C5RfjzV9yoofgRbsZt0/fGThCjHdopgUI+/juY8JVyc
4AqNuZEzHGyV/O9qQYHmw3QmuyLQiKN0qlM+ItFW+r5uhyXAqSuNxJy/JqSo+Nd1wFim6x7Bm+TV
PDgO2CJy8aboKbAcpk6icNJvyhGBBQfUmitj9xzAZh18xIzrJijf21MpXcwxebfGYRrRCokoMeBT
qfWZOFkuEXiayNba2o1G54KEiN76T/EbkI58FXfprPdfwp9IJcW7IUSGLQPwI2YLiPOp+c5+TloK
+ESb737vHAQFjibXc+hfDxGUwRzbuTaeq3ckyUfJP9r3jkRhSvCG7BBoUFFc2bawp3pJtqsOk86F
nAvUguysdTV+OirofqB8y/Yj2/tdYioTwbpat0qWQyl8ef6uAfzMvfkhfVEZsKnVJOXkf/qnD47h
x/YumBMjOq4B1gY1nJ7ruup85LroDbA5AtpRkR3zDMT21i3ct/HWVLawt5H2hJ92gVs24d4dBXxW
CbZsFZhCa0/ALoh1ka4/UtSA+Lhc/tHF82Cm3SjjaHiA9zU5ym4VndqJE+vwY7He7qqx81SpY0m8
38WDK8NLoJKCOKTlr1QSPMeozYKHdiAS/8EEgQnRGIC8RHbTZvLMtVyOciXHb+cn8OSk/m2s8PL6
TZrciqjNCKONWbkJcE0DBi7K6hWsxP7RZXBj54Z+Kw/HDClYTdsnOOkpp/ma/QhLKHeTVdW5hN51
WRTISfRlbeNEVvZ2RCc7kF9N7mvshSX1oMhah7JZIUqRuaa6jYe2wKX6MMlxRcZAlH4KdDe0iWvP
JYhxsueczaUPlP8OryX3gdZ3vWGeJKUPQz9/ve3dARNYTf5LYgIcxNZNaUZa3y8CPdqQq+ne6qqg
KyUJ8hib8+DLew0n9BEcxPtucsiVeM7I4qWWLCUiV5uywF++Fhp85/TF8veSp4zF+Z1IugpoQyeO
vSzJHqJxPZmBWa5c6djh7Au7g+Krs4hiUbbMRicd+4iRO0ISv9v3BbtaxGTlLq+KH4nhugvdRj4L
OpoygfD8RJevl8y7gDh7XaLUrLfSeFpkG45Q4A2aDcowy1C5SIf8oUKbUA0sg9OzG6NLZvsB4gr6
Pyo4n3GycjYBP8w+PrQvMStbVnTLKwAP6w9Y7gMHGv5HOOY1jr4rx3+4KEcyFJLlhiRWsV+rstNI
U3tdPnDjdHvDorMdarhMGxkQfSi+Rp88jUTQIZODf3he6Apuy7tsIDQOvSoW8Zel55EZiseM4/cr
nlV+wvkYkJd5taFgTfU6gZwX1TC5ohxcpwd/g2FKF0VS2LAJOi7lACjWRGcFXb31TJ9JfbPsSQwu
gk+m+4UMtUG4CQlh1lsPn8Vvfxd/hvIXNOoEVbbszkyiWr3TLYn31kaMHQEQ25Ifiuz1v956qrsl
sbZSsX8rRdpF8wXbeHByzzPzgazLr18aBfc8t2nLgM+IlWe2f9ZjymiMP8d7CzYPMk9icJgqWey0
njnRFe2Kf/tYjBPPJpxK9R0k/yGv1JnFSXknf+FtUcKVj1gLTsDE/POpGF4VoEGXpxn2MLFcwIxI
hTP/bHkLHnz06x+p0CPhQ+RbwyjMRIwCCovE+cZeJXVv+62L4JgyQNkLiIDOEKYB192mmSnQToMD
mpj6k/XpbvR20CMIn1bveb8gTHmgADbuXnZLE1u6p07285fnMvY21cQbxGlpYya9/zf+tCoyUgMr
jC78cpSWY/a+ElCHcTb5hJDxEKsf2ekTBCDg48kGOu179CaBcKO3E3Bp11lw/Xt3l4B/XZa1ntkr
ynTDHhXN9VKlKjiK5cWuGG5XBXmaRAI7gEBy1J9KTCeEgsVo0qtpGsOCmVi3PjjXsG24DkAXiYdP
6oBgxv+B81qwWWYdklYWdRkrerXxsoy1518DAvcC20Y3ou5BBgq3mdGsfWghOZF0b8keoGW/NXxC
BZZzdx16qgRT446pw6HSPuDxa8I2eNLu8Bs4ysCLMrOUYsL1BAjgmMmxfQtzfi6zzMifiMIPANiV
5mreYlWnZStxjpPJmSN98no+jbMjN/oVVXoL4rf1dbufNBTAsjxOOn5tgUp7DaxDM4wOQ+2NjBSx
TmLrfJzMUqrb6+DfuvRQt/8BBCOrhd5d2ORtzKk0rvGfejyl/G4+0uBAUsEk/3Bcp/L4VOeLwOP7
7G/2fDEIRaqV1iDzW6/ud851Gv4npMcAijNu3ub3WLduJgbOXpnTOhz9b7Pv7mCHxVa7BPApwi3Z
jamL9iwyFYarDaM+Lp8qfoWra1UXJZMUlN2XVPnzKODs147Cu/BByXnuVxDuNDFUF0A9gMcl0hI3
3RJcdHEMscv6vQwEAIcET4QLvXIDxSjBVrQTc9atUlkz92rzWvoFwB/veH5raDchHSGD29wde805
B7/rENlz6kQ652+xFRsTCm4sgGBAL/tkdlxexyHzNb8VPbHTpmlaHaLyVTyIx9qVsR2Ty/cFWhdl
9DUYoNt3pMNANxRIoERQ7zP/6YagsFgXRX0b++6F3m2RN4vijyDcM2uh2YqFasVC2KJSk4R81iLh
zpMAVoItSpfZOffkO0QsqDaz/nrUAh9pvKVWcXbn6qSSlWrNZzY1ZjJc4Geq5EbQc4OXDhLk0/yQ
YCyArxhywuedw5Jemdax6h1gahS+3oVNSQpmN0PXD0atwGhAlq5mUGBSwdimzkoBL5bPMDy9wCDA
2Nel3qqxI7PyaOQB714GWu9l47wIBweywj1xPaASp0IrFOhcOMB0oV7pjHnhWzqrxSXxjHkXb8RP
SuWe9HoPpDWNIfsqvhQd1kkmv4KEk1XgylyuT8GwGNxiyPbYX3VMqGOJMzvTpk23sZ1BoKEDTXE9
EqOlJuI3ojtLh+jHQosNZ0gXLz+aJY5LtunU6bsigz1/PnwRXdFig7LIBPq+moDiggb+kiHoy2Z6
sy5xwqXOiQ/yisJLPFvK991pRj4xlGPT9n5Xl1XwR3grC+LmeacsMpKBNAmL8+MEAjApUwDo0oxh
w5lhZjaIli02I2b5kQ64B8tc4zpW1aN/aqPI+mu/uEXsp3kZDGsQw8aB+ncOEM3Je5VQIml0JVxh
5DOJWArGmGxGYiPbjzKQzBkxRciLuQM4JKTYRrLgXQiSP8CfyR8Y2tmjmMaaU8Uwijjk8d7kbtdB
y/lpstUna/7lLoz0RjL8VmvKPIqUY1ggbpMbWygz8d0KM4FgaPv1Cwn0WtlyV+MPGDpdjwaoP0qT
ytJKLkz7MDmTZGsjvkXIv0R+QGdzYe4IRjx7Jj5k0nVh7RJvD+xTGwfla8Se73dNjPRWm9ie9utd
a+TG832/GDW/J+9eEAw2AnuhcV8Q+jPZE0/QQeh6aVOE4GMxdELyv03n7blb54yCcTIjs1VtD/Ty
UQlIELyQPj4+g6oW27lhUeq6b26DBxRRf4RPL/q4RZ/t4NmcH+ff/rNl4gvfI7DwcsStGpyzMDM2
cLqmmYzAM75XqJbT2znOIPn9iQqsnAJqktHPRNrpaSvbzd1s2/v+doPMpjEoz4YenF7K2r2SuFEk
KaaHyTnZ73CKirkOf9Dm61IrpynReH/ta1g2k9KOhsP2FkZbHbETbOAgVdagcdynTEusesHPSUFe
QBJeBvJFhi9LOltsqbbKOVjWFu9eB9UmcIv7Vh3a0kRNVr0OZ752xNdZOXmPa/rloMrhOidvK5d0
LKcZBFFoUuqR3X/LyPIHUa1c+EH9BmL6E7YuGUkJ0mB0B2WecJwt8O+4bTA1GimkY5utOKIsfXg8
tnprh5O5FPhYfRYnVLlu/fUl0SIFQmYB/oMLvhbP0YZStqxayXctWn0dixSYtPAUwezYR6656G6r
AoQHK2phTPrSId5s4db7jiCXFEnW/TAeto3xZOEpZX1mPPe9JJxho9iJAQX4F8A/gZdAmR655fEr
Uf5Tg/LJLubAb1JV5F+G88ZetZaLO/0HYB+1j71R4QV98+UGqZi9OqaSkN7hZpDeYcrdEZkopr5o
NuzlaZcENPO46i+y1jwfQ1MtETYB9C95LtW2agTDCIEyk7ike8OvOyJlYRCn2rHZ58tkrrj0BgN2
tr3O5DmYyF58wMdlypTgZtAyrT6DP7jHwM3vX0zKJyCatAGkntsx2+uDsyM7jWrgYz0P0TdNTVFq
o/NvCJmNXfYk7XVEN3E6JMCcbXGvci9kxLn2EY4Tj/MR2EsqH82DzeFiDBBVW6/SqncUrWaw88Uz
KWg0lNUvhy8DAqVYWMjJ/b8pfIQBONCYPxA+wEzQ6xKd1JXtL/CtL2zdPOQrBcdJ+QQ+XB7NxnBp
Uc29MRtPWKSvKmV6WsYm9xZmAU9h9pBHVolEKlyQXXCpuGL4L8oCtfDGd8gsdjzb0LFyJ4PnyYjj
kAMWu+k6TkraAH+QEP3VQVQZ12ZGZLSWNHPbq0YKqK68+lXQU4o6rk/pzA3lCvFk8uyGgKYdmCRj
YgJFL+KYGSaIGRTlm/1zwLeWAmep7EUnjpstzXtHLWYmgJwDQ1LUwqEoldhIMK9YtX7x4ftvOBHq
LQsQS1jBRrXf5C15FIBpP3pL7R4Gt5CMJ0XO0pc8wRAbfmvRJ5tLgo7bjXPWiqv3eksRWy9QFwPb
CQ3Ogw1o9MlZaQlf/7Maojm+gJBpBrQJMGKJmTpVcZw3KfP+O0j6LTkaWXuAOwVkFTmW+/R2kC1r
8iXQKwjf0Yx2va8MLBcVhde9/0SJiaCTx/pRqu9wGksC9mB7LNmR1xeEQYogTS2fnyLmUPAvzdkM
8ywHrMd4ZxdebMsDjDwBN06wXxZr97wpG2YY+CRSBbY1OgXlr++5bzkISTTrNfQ/Va6PnENjkpXr
652rACEPE7U7s7fBgnb7CvnKlT6WPG8yQF3ODpHUdEIDJWW3MGxwLDfaQXJSk6KMbCb+ztN0BvHN
Le0dJ6ze2MDq1+BTzxU+76/evobEq9XqhXOP6zo2mzsZySVCCTA/l4K2tezZxGyT7f4iL85vODcz
FRoK6U2s+yrTQeizkI+vwZHoURsxpxlSrFU4iUQytezddm0rehSz+ysqasA/jEYvLoSjJuwDo/t7
luGUFzcPaaL35FTgbiWhjj0c1LUNdAXmancAje7n6wD0S/YZtYYfv15GxYJSLp6RZKKwQQk90wWn
dBrAdSLnMoGLWjVBLbSQwWYZoGityjvBPU6ZD6uaAynKANKIIU0NORa0OTmInPqHS8hlmHA1zrGV
hJfylfQY+kUFQlpImHHJHKxztVXhbWJfyDsuVNh9IgluZklYWoK/kgqSuWstpoG0J2oAkE4EJCDA
07PnFQj+uQE9ytrh369CZAh9rTXYrwTZwLZmZaiXtn9k9Q4Wz7ykckAbPlipXA46yuBabUUZOmaI
U2oZaVf9s21Os39I47gdW5tQae8ol9zi3jZWi23xnkpUl+5sbFpEdEnuklKFAmckgJ1W/iQi6Me/
4JhZPWFHtWybMj921RCThRafAWRHkosu6urAAimXBVUEwz98JIaprzzN0FfmbrDqi7vE4FkxjHng
1Cm/ps06G1wD66LHCOYaTtXviqyXFwRok4EXUn892aJnbgWJLctKmBnFW9h52seHKDKgJ52EPk4j
ya1+pA1LbH7hsaDnkY1Acf8fsrbNEkppDD7ZLZlJj0BlDmPL/LnGZRQAJKTV4a3fOBikUw9oAWK9
7GVZZGRVgddVFrhZKLotPlzveK9qiTTnS+U8vMULmP+1K4eDjDGnGpHMvAmDzjuXwxS2ljOxEcGl
6iRlw5DkAh543sAbm9D5Zy0i8iXU6Z3Cl2ca1ewaXUUoSSfkyrWw6Pf+5iYW7LlTw16ne/5h3tQX
isRVWkTUfRQ6msz2PHaCun46ezWq7Lf10FRsb1WHSd8ri/lve6Y+CKDdPUq9ugL0tThjiGuetUd7
mUEnRok9S6KAXZaNKUS2ZOSbjQK8R6Fucg0Ibn/8MBIGHnW1sMxFMzNJTWEcAacjkpOy3RRzRd9z
l1zUleaW+Sf37K8kNt+/w1z+XCRSTlGaeMPnCW9g9XmRowjh2+jBeCILigNEFVWtxotUyjOTXyhI
q0/lTgCkgKRuuapD49d9Dn2sh9naxr2kUHnJUU9LIatXGk7XKIMhl0IJaSIKTRy+knO4eBVtkH9t
+0WgiKmcxnNKM0gbnPD9jnUncWpDD6o+Uji2FD90WWcMHcL6rtMZDYt/pZqH8peOBP5vX5HVhN/f
m3YUUYLTDcDLiBLiG682qISGaJXwJ4tdfLeeWpQHi370hJvy2Ym6wsNI3KgdAHQFnAocuYvlXwGf
+Q6SWxC8bEEVe+NI8+S75KqpzBvAHbtl9s6GUMpVlZPTbyhvbITyeqmbeTLMYBciB+8oJVj07smm
pyU/bpj1UK5se4gOA0Q86PKaKdpZpoZClC+DGZ7aGjMssc3C7qdEyFbnRRwluc7MO2XIhCN2uwVj
SBFI2eVxToPKSLNwF0WqPV7ooS8axQtU1gvPR4uz03fwtJ/Qn3dgqWa8P3H/UNx9jDkp+Nn8cDPC
LfIyHOkHLxWm23fp0lULkeaXni/WzqzDcHHtVaQ/KL88gy7MEAVI7wI5sqmrbu+sDjMu7ULahZYk
DENp8xZE7BGjIDmWcgW860Cbn3Ef7CirT+pafPyj3ON0FQK4GD3qVOGhnEPRg4UyGwRNmEyPcp2P
cQrQTHSDWcGtnpUQBQnhtJhkKchD6nZ5/SE6ZTUaLrQ9ddQK5Wd5HPzdfZNS3xJEmSarNq67JItj
3oK0piHOXvkmBvgl5T75pA8Ojn40Ro1pewE4uQIwIkf9SI+KXbboJv4tG5b2YOUnUCGtyID/GvcE
7oJFC6qnUvMFSDYnom6Ewv9nWMkrrSnkudKvYjs797Dflc415TkFeTwLE+79fkOi88itV0Azob6Z
95RMmCX6JooC5bmKGh/2GbHXVJbGqrrWLdU9Dti4sTRrZHjqEJyPOyUDqbkrlNHEGenCn+bjrNay
EE7r/Dd70F6nU83Pm6+G1V7+i2akbLd0p6O2r9QN3m2bSrg9wGW6O+qWrCXkJCrnE7cjIvbZ1erX
i6IVxbDn2a3KCfnPqVX/i2GSLwTipdj0brauYmvFAfR/SWKjgoyuhrASYR25AKy0DFQ2GpbnaX7S
zajlS0Bl/FQxMLGqtpn//wGsl13X/XoK0V9SBSQIS/bvdaGJejrGIJtSmrBwCOrmujDavybt1GlW
gnrOrgpPr+TEe8z/zk46d0n4F+PIyjRwVFi4oYF8bA6pXrrBpvSobLxCGZ0TxtY8abhXYrcy1bRR
qHu56AuCQorK7HyKQ8BOvaJAVRDjCboqmngKYKeaa92uLse+KDqAvPAYgILR9bRiAYz9a9myrqr8
2RSGQV/0Rs6P9zPGOK18BvIT7ZRn+iJjqL3No7qFkfKYf7Y+yN5Hmke5/Q1Mn+Ni95YREaOrRTeV
UN85zCw5d0JW3S/BJP/LWUZ3Hspull5iYpKqZ3ZPlzDjTzGQOZzJzqAMrFFdnuYyL5Os17ViH1xS
RJAOR7+o4kEM3eN0/9473r43ZlNbsl/4wqgca+MlFVZBInSF3/jgrjRIGqCuIFrc4YK1wZU74969
WWWCqvf9Otk94HDjjDxLVRPi8DEGdjg6SSV5PsxYN6qNAlIcAu7TX90eSqhdNEhePgtOGOcEKlst
XJipxVV9AXinFC2/0xKJQLVM+bHwp5I516XEcImbSlbV0B7OkBLUg8cG7CjE4h27g8sXg1IxZrho
pTq88F+/pI6EWKWtBzNHnty2eoCglAusVVLkXCgWQyPr08Nt6QMvbMb+4j1r/fJKIPQB4vevNu3/
6H+BDILpJxOr8JuLecHLngYHFWprshoHE6RQCH0MOG0adT90kN0/K58ZJwpkUiekSx9jPxO3vs2l
01EX6813h8zvFbU6h7Qv/eODuDbQJZLxr0MfACWeHfmIa2LmtGCMB/VUAUAWKcCpgFqmx0ubTyzl
X4L6BK4QjlCGdLLt8gZ7LNd//b/t9psOXwAsSBxq40W7NUSSib15O5TA42vy7GH6ekJP5HaFJh3J
8GPTDmN386/loE4yI7f6KboekPHV8ZRbAyeAEMk+O0UwfdjLWMASUqtehB8iNEDApy2b7FvyG/bP
ujQ+pjedNAabVBfL1GAAcoEASUMpP28XiiuxwsNFW/rM/DnXXxKXnhOAruEVqrOYEUqoL2bnVUGZ
1pTsjOb3G6sEqYiFO0pS0samRMrvMoP/YwwFlR7HwmAP2PSgOZbmMA9dfxNeSwR40nrPBmy2XiAi
E9E+Yw4XbdoTSFSJckSU9+pMBPwKYQeQGWw/TN87tA5j3VPBC5PKwP+vHOuSC26l7G730AQWgKPE
tZB4JHWVFK0tk1Kzn0OSkh2UJmsnbnaGQFGfT7BXaF5JiY4ZdNrvPIXQYNUbzCnCsw2m90aNJ1rH
hnc8tCbW40fzDJRbEG4riu20E47nRfA2uRxqNWhBoxmfWnVbJgPrTA0xC6S8RKeQfmUxLq7qgNIJ
HexDV5buDzCOs8e6XUfu+SBd6BlJtjh6Zl0+ZmBcHFm1MX3/3srva4Aj0/moCCr6MB5ROG9YVubE
/5GYY/DtDuisJ8uZfm90NL2HRjxOfA48pQCqonvDk4Aj1YD2K60CvKMiObO7u1qZH0nRHog3dfg8
2o/Mcurbh0xacz11Kw2Nr/uFNb6Z1q1QIPlFNjselEmVNDaqgXNDRYY2ZbTA1uyrYrTTWVHQ+faC
cgFFEEfstsZZ9bTtw1h6C/lkx99sBVdHxC/xB6DicqSXnRdDAiDRICWhMoOIXe/wT/uc29vqwkj0
aO6SzrLBiSiqMge7m01NI8/ISeiyq794ompXUJ9Q72FYbJd5J1JNPd8muJpEiYbpKBjoi6ae1t1o
TD9GHhF7NHCBM6NHgCdCnRtM8nIvkT2LVHOHT79Owau/G/86hleS16ufZuuuZeqi+4iqGNbMb6zH
N6rz/0/uxp6Foa/2UCJjo8GsHdmCBYWzUQ78GnlHCzhtWFUkYX0BDC86IaxhpZzo3ESINdfsI0i/
RYfzrOVLmgrxukz0garSiypjcdnELsQm2Sqshjui6FEgImBEbp3VYeinNWi9dJdRpd/vDeQT7s90
FQSmimJkWD4NJPnFNFXKPbyPE2i2vZmfGniOZbf03JY4t4pxoCbZ/qdeYMur6Og56vXDpXs8MuII
T9OkXW458Long0mea6RNotVQ/LETTqE28UEDztyPcOlulqbB4wOGGVh+RR6+gZS14NmRZqCgpd57
lX6uKNUGuCUkZmhwcWo3v0eK+jsp4UqwM6bk+2se6sqZNpf/20ZeYirDKV17gWIg7O/acQ9RquaH
W+dvtpQuoRRGDYsXOwq3Ze80RIMNg1KfgMae5mkOc4VGMPiV5aRTeAElY3KpfZ619lYDp6a45FFf
rs3FfNoOyQjX/+TZgFGX71XuuTe11/yyWcT5tveYhYOKJ+x2j1chQIY2DnGTqJkvzHWQtmdxh63N
7BoPiKHRBy03UkurrQU5dkGBGXrQqpRrx9mRQAEskEMGf4r+h2so3goikMNaYdN3KNV7RqLqk3GB
P1S/AsZpjPKvBWDrCeeeajN2RWCRlRuBWJlaFh0VuiMGEeu9skjDHJRNatMkYooXNdIAPmkp1y1w
oj+Z+4XF8VX345OMvowbeVG7YpxtXXTwCHoqW4ds5a3+I96ncuFp1xThECPl8rkpZ2WOepaxx3yA
Fzgo2FZ+UlbGRKs/M3tpBtmULm/Ns4MQZ7oxAsB897NMSHDoOrbYtn/tjbMjg3RaGYZ6j1/8tXBu
9vt0zhChjk2ZFyTqMUbq4CK53+9nrRU/0VT1P8X0BGe44mSgssp6049Sjn6WWi0i+sKgpGe5Wt44
fLwhJQyu0+5HISslKlS9fyNsGDoh/3oJtFKk2uGJ7NSzOXQiluulpvxyTlRSUIyxHpo1IpspYqSW
K4TR2ERyfqYu/Vy/FkUnY8uQLEUe+2fcAVWbAb44bF+YIMftRK9kKWW14Vt4p2cuI3rqPT65d2dW
GtDsJko779UKOKKyaxhtvryo0tvAMuZbqnYJcSmVQr6QfibIalzPP3/d5y5MbHad1r/3UWfokKgq
WkwvMwF+f6Ak1JYPy/Gffv6XU9Rud3MRNeRR5b+btnDHF4UP5H8xgpbURVTsYW/+/8KFhuJXAJ7Z
gTEf3Qfv4tmj1Sipg+NLTh44RK1SHPePLtJQm4Brxk1aW9VUhLcYqtnx+aSswiDYzJcfqrCJLuFh
dIupOgznMLmY7RWELA9XqoCnYf7issCPtOF9OF8nfylan9kqo+OFNaF1LFcsm4Qw/8Q7lv8mWPgj
k6NqfZ2N3fep6lSUUbzxuhrl74Hqz8rApEvrn5x3TPgd3ZFnZk3jFffL1aD+4CJtyt09zyjFtri/
1NpjX2MiI266mSIw40oe/4wOGGDGHjBtkeouU2SktnHcN11ok9zirSA9ohA82AD2iv/pu1jTNh8S
HuXg/e4Xq0vkcZW4zBXUf55M3u5d5Ru4i9M/l5wa3uU2336q+UsGyTgKEb063/Q6zzusx0YL+9te
mmmuN6zLucIoMjeAv9Q94zXyeh1TQSBZPz0rFVz6odqBRWqikZ/U1wmM437DI3Y2cfBzASX9HkOK
DyLMoKXk33yIRZ/6j69w33PTpI7KNDMLSn4vOVQ9FRsY4AnwAMueon7IKPgmFp0CadF/tu3Ml2oR
+qFatOLn6yj9KVLFkZODRK3eTfwhk97KfjqBjtiX87a2N7yKeH3C8vgS9VFc6PYn2/wT7LgDn/Am
xIh0DbIsg/pAOnGP3uWV5xQnGLpfdiz3MCKadN5EElVaU8DOGvHSHfUZdITQJqP/82hLfo1l5qAK
FD0Nn7Df0fK2rcr1JPIZ07MPLKuRGV+1oQZ6D6to7LVLjczQ3BSthhcqxQ8bD8f+03S3b+kAvYCR
3aLPL/Qc2F80S3UK/LDxzI8UuJmAQcxGYllZHOxe9ePNjDE6FcitQq9uqhmGNuUAH/wm96jGP/9J
8uEYOOCyActGMKu76laH9jui/J44QOQMtur2VPIO4lp87UIHv87UUmYGkHq/T8BWCQ2IzZNUaUwk
FfcxRWMiPVk/EEvHkFKlkSKIQm8vKmGPzoVEj49IY1E9LwpLX0tDjL3N7/bXIun+avNTTe+s+TiO
GeqqxmqPnewQ3A0jtBhrJTCJ3MeEwVjdKeBTViGx1rqJGu993fiHL+IXqKW5+18FK1Mt9iVA3cXd
ZZL1YveghI8uBnwNGNJIfDwHQsLtgLuzuijDuW/23vn5MxFhO8GpdtpY+34xGKLMicOzvBxhe14Q
5FLrZ5twWfZi3h2dNR+/BdGSdtQZAuCZ8+fRJPni95SWkpumejHqa7ZxLa4WKb2tG3Psyb5QLNHE
0OIIsas6Z7prCo6nae0edVc962YGhL9PFnrEjHwW2fr+J426OJX7tyiUm0p0AqafSDVm/DpR2xbw
DNpNOlRfQNarPvSA4AAW/k5qg4mQY99ghBeITeJqvgRaJQEnaofyQM97Aa5jQn9vDQYPR7aVvtQk
4gMYKw6DPY0ycnblRA/tjJCeh4Wpf2mn9rKWZi6YYmGY1EVC3xWLE+bfeTzp+KZK5EMFqupC2j4k
E15HHZ/8a1jg92UYlfoUFox7h3GQH354aBi3TauzIrA5hFsbfApfVrF6kzVf86ZCJPFn4gr5Na6U
87OvQ3yi3m/RV58ecuGdLVfLJ9EQQvtv0Ae/4gJYJFRHZXd8KwfL5cRgyW3JslM2DM1qvuTLH1zB
F6rItPRESrGUGN/vAy0mejeoluQKMKi1Xz0OIcSRSBtYmSmlKtbUgPZ+fCHUju0Vus5uXyTl5k0t
qZLVsvVhxDShJcX1AuAyckH8GaHjLxdbG3NrfnThQrX3Llb/BixUAwzqKKTpWyEEAEJ1opGvfr88
TvR571SgwYoe4ZYVpW2EokrblSmh4pjHpI4Gqp1mRNnjX9+UGNYOq9p+xD6YP04xkBnMY252VTxu
CQPntadAq/yljtHFxNa1xGEt8L/t88uQsuYbb6tG+9O9ff3O2L/2sdsKxJc9hz5F+g7YtdwWy/6e
dWQNxqp6wsB70aDre5+3mibrYXPw20bpvSYirfQ2EP7LwKqiMxZBX+cx1i6DakaTpVhTKKF+q6zm
QKoClgGZ8NH+5iqh5+RpNiTPIbEmhRXgtZJR/Z2ZsPNO1Pef3JgogibRD+mnr6ujQ/mJYqqbijOs
uPKgGFincVjJ2aKI7tvF+uwMiVRD/GmuORj+HkgmsLEDtonflVJdzFICFl/ClwWpiQB3yQx8pRrt
uknjVXTtZp2oyvsehY/pXRT4WSPd9Xs21x7kjSsqYrkvdeXZCiSo2oLKj7JHASyvaXY8zEoHeGXK
pod/6uBj9GzixX+9ksfSWzQ1Vq/klpp9wCtRYYdlyFtTPqzttJphOR6VPUv9UZNBhHDC/gB01Vtl
cFI8hLEgzD4sG2qgSNPeAz0KDtiQkPMDXbCF0dP/Gg4gdS+3FjQslsIwCqEX/uwlNfQivU+IZ/wW
d8veG8oKg9b9/5r2MLAZ0+0LlM9Ed+nfLlZgvxkEO7EXFOCTC0RQhG2K1xcEfgoC33Cutm4MJhzT
eW23D2eV6sWktPqekgBTwaNt1e3FPAqyNM87Q+TO0/ipzlpknczows3piXlPRKtf+PRQu3ygJm4C
oeK/LdxPmP+ZwTObikUK8pUQNe+C/6PU83u27fiJZHVLvT9WW0djaQXG2zG44z6JXrqwuyPk6wuH
4KgujwDS2nnWT0E2At4tIuwl6WHIT9Q5GfKsArJ+6+RaomfT8kbJIgZdg93zWcGF0vDmCwIolxKe
N968lZGI+8XhvQHEEKmprbvV11rhpr/6ML13JeeemLEWi3wr/Blz7rUvOsjIXj8v+Dit+F24Z5Qo
bdWheYBykrDSxJvwXJob2O2Mo35CpMUsGXpO8IAhZETEDtfhTo1v160YHgWifuWy/GmPFmGIc96r
JKy0Nh8mQV3k0d7rV4VtMiDfrpxNC9doLJsifwwFd9kDinpp6Wl0+ZplF1nygJ9HODqtpbR0671N
BOaSN90DHK5DH0yb97v8GfGZD++ee5knEKeifRHXaKccB/HiK1abu2qZYL33GGdI3sa90FCMNme2
RSuOUoQSb9DwqSDB755kMPZ7LkbEaS9rem206WF3eQxi3bPEnh3kFkAM9efSiPsJPt3WIphKvS2E
8PzP8lCz3CEImUnqxp0pKDEHhC4NWzTHl5rUQK+QkcYoGECsf/OOZcjBUowI/qTF1pKxyAti9fv5
4gyGa6K0LHp4fQtiymnd4vPpqkWb4MwZ+1JK6+ffE0v5I2PUB56ltdcY7xOXuPG20U3+4Xy/XyeC
VEUMmpmFX4+ihtHHZ3eH65pqyJANzSv7G4uC7F6/kas30MBemoMDNceXXaIL8YFzhiYhby5uFSP3
4iAMltGBVWG7KtvkxU5KmBhYBJfLfer+KTuTx5Yet0bloqhAuDn431+fJY2PYeOmIGldX9PfiOyI
GJpevrqgi34EOkVFOcmulzDiWxqzhh5iN/uJKTw9tJTTWBy8fZrW2P0pveE0ElAKc925xBxHE9fb
psP8mWLNp0/hTuYmWNM4a8MCMMmLDaL5ks9ODg9TaZCahm0snt12RzblKlvPoll5H+IhfNMJDzvo
ULmi8Ek0SyvpXIWNqCeT8VySiDIa/rZIvHd+MfTSybx3o43NhRKG8AQDuPd7En3TeX2HCehbvw+4
lZFaF5h1p/iVE7Lk3SrS1ko2vptJ+0caJojOTmA1zdkRnhaKKQJPWlD35hUicD2D0pfY3KrWHEar
zNRfp+7GURsk+k23ihA6A3u2UUhF9OIPP6Xl5xuQ15iejawFBKSRBDxYNLUVvjs3OOCz2QHMRhK3
J3TGTgt0ljLon0pjV214Eki/HuyqpMJlRP6ZR0Jf4ll+06rfLnRlfQ4pu/Z45gq8YZGVONCe5fvR
vwwQh5QkKUweYIoSs9SjKjQ/1ki9pui21hOL45svQZ6GSAs3zEUvhW+1NIDZSjFWhycHup+QIYNu
HmXflxj55ixI7BFfrPN1/gsAuSlPSWSXZn1MKBhGn3rj3MS2xJJEnP4ZtQ+Eh7UIWZcdGFGNJrXb
kUD5qt/G/PUAJjMtp08t145PQ25BAIXuwcui6AKcnWOqUDPIlkMVxs8UgtVPAqnai9xagPPkLzde
DR1ETtSJDlbJkuJs7omdcC0ofFNP6TUbVDV/iFsA98yGYiIT4ZtbKf8LO3TeKv9CGpMlqNIxN783
iNqkxw39nQbn328/3O4HBkkAHNGmgsch5mtbkIJoc6QglHHO91z5huuxCeSxhWrx+TpnlqjdMV49
50aaUgE/mk3cEOGK3XPYfS9qAtpP9T+i5CHPLj/MsRmV1aPiejFovkf0a85uhB7e3ufH2xzYjaua
a4/i0Fd6C5x5vsk0vWlIidYIolM5VmMzQskuyW1Jn8LcSJ1dGbYiotv7gwRyx6UzGDLBX5uu1PBe
SX7lT52dgfSfu6iIbQxTzEXZxGoW4J8SGm3rhvVIpAWgPQtxkPdSyiGNBaTIC0+l/7uSSl6MuR1s
qp4uvRYEmEfVvAOsZkeNiTt7LQtBBISUTvEv+olP8r86bfFl29bmC+d3eK+YB0HOSfHw1uGyorQq
B5K5Y7M8o0NAkVg/uoULOEMhpEX2FTxZBW8XbqP8lab73emJTjiLS9ZeLnpznK0QAT5fYLrY8mtC
B+nD6gd31rwuQMMgYvXSueZNInBSg1XjpMuPYG24HQ/gr5x3ExIQXAGkMb7lMNOObooVCYROIrap
PksXIVPgCOSNBYlm650upr+5kM+LyFI9jSRqm3rMOrCfGtDwsrXtWOWb8GHMcuNG1cJJr5e6HYVq
traxuMaL3mTwRViNDNEYIoapD/YKUM7sPTcDJKfP4yeIuDm1MqCcTOsV7I25/Njez5X2nVdKhn/h
7iozmgY5rFgcvmnW8xAU3J6t5GALErslPdCxqS3UnNDubeHqrfDcGFwo6P8Ns2fIiH7tlmHvPLmV
mfYUK9iJDacODkb04quk5GL9HlATbnanYRp8cdfhQxtBsY24M0V0pc6uroJwqctnB2CzgJUNVllN
HJcD9EN3aDI0GndpDgP+oFxjpaImHbqPnGPov7WERoF/2hGcHtyUaKwS+159s1gYYC2HjTUd2lv/
yiacT9KwPbpirNSJA7JtR15xD+rPABnftJL6wZ05OyNYN9AMYCi6rkw/fDcy5hyF/0LstWUffZyP
s7dYd1oHBi2vWRFxVxB6nebLNo8vA0IfS7qY+zB0CIkQ06w2e4t109z+GDYuCoeq4welYTREmW3N
kxqeUor8FOtm5HgXoMmFHTHnvK+4JR5+TmVe5AOr+56asZSB9Af76mWPGRph0wm5PCflowo2TaCA
UHHD/NHQ5OECQjJMZ30hATW2pjHkyKVpwIYHRzEw4EsnC5xJG1Uwgrg8z0Oy9zawTluVtexH/5mW
mSs3jXRj2Owyqgkiyzscall4xME1IKX1j6rPIfKD/oYPdPGYvRGVLfs6tUKQgwvHvezlCVRMj0jd
jVsdd9mcyPDzJFCCSMaP0BHHgxxUEC8h7wotS81+8G4htDdppmoJ4uRbzrNu4WVnWG1yQd91en95
yj/WFpy4nwvdpFRsce2oL5PkJttBk3ORwDQO0mHvvJnKQteAOpo83GgNMRltZyKxwIoC+qA7xUh6
pToW5za4x+PjBDzmk5XKD0XSF+FhYQ4gjLXuHGhOb3O/HWWLy82C/7v3G65vQPqxMZ0MBaZmPQEZ
vE4m1Mzt2IsgZNYDRQgycrWa0i5ONnsOPIoT2Bk4Dx4sHaCZZUK5funCjEDYoVZDtEOy/MgzmBRb
9ZOquXgCsaYU1Kp49BIyc+0asiybWWXFcxVr4NEOwiDUUqrTeyWgs8GU8P0l/8jeTWvsYrYrb9YR
bBEoCvZH0ToqTQUqaAPGSK4mm3i9j5U7gre+Nglhindjl/be/1+RI2offWqsAzfbOA3oIOtwAD3Y
6XsHusJ2qQIBPbnikcOABoynOiIZtSfJHn4UxcJPqjzyaPZK9wxgelXAkrjCXN5tSSnV2Eg8LQV4
sf+FTJY0CSpepGN1eMgn1iLvuATGpRZUsFm111howh8H+Q/mhrosopTU+CprL2L7XOr2+d6Corjk
LiRCi1X9ICChftApytJOMyjyzajIjWA29onDAiX3VQcbxdL3B1kQfMVBml/RoqqhqrX3oqD9I14d
7Po4EHTwH01K3RQ19KRltTA18ODR1ykFoZXL155wpnB0t01lOwAujfinBrjC6g5wFVueWS7oNrs+
vF9g7RYpKe2bGb7vacLKunsPdtTEYiLs9q4Z0k3ATDkTfiABUzC6tPqP/SpYwlovLtNUDTZgJ2ZI
VTWaPE+cAvPpq3JKYtpY+wlT05LAL3h5BAP2tlhtS8n3MFyIAbk1nnEVfOquySJ8awpOOsG1YrAE
JOVxRAdZWa+0ZqHgaXqDSQxlipwUxZ9cYNS0M3eZcLBcVGsp07qUCedQDyGwg5nCLL7jszS7YYcz
qUmT866xDy0ifp2ERW25QaM+9tdjMiWCVR1hAAWYDCOrm01ajXsV1cIuwnZv8ofJ5p0jxw4c30VR
bHMNYEJuQPT5DpIrt5j1f1mBt45HLUmXK/wk1U5UnBv40otosacpzV26XOH9GHuUyeGu8y0VaYkM
G8LTEC2vtDjAzg5lDvRRLAv+HETWR/npfsTZGP3B1PNStwdUjMDMflGoQLw8DSzphdGvhxbLi3Ob
II7soMZG+qCIfSwh9hY5F5EYy8Pp3BVsaFGk+o+9Xm9vPnYHjZTWfAuEgWA827F5zW7iRh3UTRNp
QtYNo6/N25OJ51FTz7+Ufaww7gyQA6GCME0TnPvy/C4qzs/1cTa94by1yJvRj0w47y5aeUl+ZTTY
Kkr+B0kBw46hVS5GkuscKNMVrIR7W/LUlHimDkySX7+tYyvE+i+KEg3uf2O4p6nnQz2S0bSFqnet
zyvjKj5S+XIYhd8DllAaC6Z8Mj4HjrT8C2aliqKmLawydq63fs4HS/6BAZi8I8Pq55Lz1eSiOjBe
ctuU87+ADSAB5fjJ5buP5pv+53xg3Y6IGwArb9ZWG9nN805y3Hrot9d6gn9ynzRhKYh6hjza1Cx2
A2zaIxT0qBVf0x+B5i2W+2rRqrFlCDbNXLI+ecr5CeTdmj/d0SUOmmx3HLZ6HUjjc3zPL1x1xAnz
zmEr2vN2vwGxIbW5XeUWtiol1Kr059DdX3g8rSnJ3mACCphKwpBvBZ4qdKLoCIZyv54IIwKJKI3s
eXrhs30OhvPtndCFMTlvmIvii+HLQvqz87O4vBoE7pLQcyCqSZwtB1JNalF7gmvL4HpU208jhWoR
PlvMXFqpN077maJyN96axnILLcufQ56DT2rKYFw/OjV1+pKPjg1Pl7ybWlXOvFywtBWbJpYoLZsb
NNrdaUvEQheitfDWJLTYwjVqb2gWkk1YmzLtlPt6zrMFiUT1ykClr4/FAXTufKNcFqOxwdQUD6Q2
SNAasbUD2VWI/aG521kmAeig6vuXdpeBCkcJ5eT8FJ7OtMJGOP99sBraSHLhOYInI/j+0kQ5yXJw
mpjNVLJ4TnORRjrzsH+A+P6aoKaWw2uGVAGbaapIKjYkyCosZ4GkZ1EdnYTVIvoXx9D8KEdmvTSa
BOOgT0dQp0W38PJQhoEMBHxoMNxWKigISe43UF/7xceA1zbnhsGX/Tf2N/Iqq7XL8RubUzQIjH58
U8G2/sf/vKeTxaZZBLO6MYX4oCatigLZ/l2vAss0KUORjI8oV09RSIWBnmO7F6mCz2xt5X4/ixEn
rUBqy9pnxI3qyBcK+B1WuJ9HDEBZguDKjj5pLTQf5zADTZPxQGMVG+04q4fIVhAYkxXOh6PD+1Ms
G+VFpDVdjIf2qTZZ1dS4OVxmbdhrqo6wIteTxE2uU8eMGqcydamkuB2AzkOJxNDbeKgZzAWwxw+K
TzYSbS/XO/R6ZVxJtzRYChEgF7RWlRibZwrsVwcFAmm+xr4SBEDG4P4utuxMhyr6sabkpX5N+592
oublhuFEKnt764mhwSkhCrQk86hQlHmAan5aYfuyJjPQcNzNK0Dk7MO1fgYEoq05b5+7z/RI+oTg
ghBxUjVkj4Y2QDsYlNUYRtFD0Ap4TvZrvO9hx/UzQ6EIKsEl2kkX0Xj6Oiwg8xZ+BTDajYdJJRhT
uWUMb1YFcSNH1HGv3iU2Vvvp+QM58KAOQwPdiQ8PZy5C9+5+lp+z6C5chZHPfLMLUxUqjgQ3IB7t
juY5NgFkSzkqwNRzPDLl2tLDvSNVphZrcVQiJVh+od2W1/i+4yLmMmNvdlNjSF7sT3t8JKm7Pbtc
dTFYcMj8cSw3ampfRAMFq7MkMJkJozQTl+Mzhq3lpv0ojAFoPoyKXd/OgNCsoQ6LIqSZhg4SFt2t
JhWI27Pg+xmr/gUwShpeKNzCx0xxw5aIrhas1VkAnFRUZwweaknhJ3tC4C1hWPjHZkJ/LVX8USnq
LspaQcVbVDDIb1C8j2gFHMzodWplt5qKbgZHwuMfr5o0v6q/idJ8v4QGCypLi5Wh5i6Ko39N9AJh
ZaRFLWdujd9yNKGNERNOeqjFtWpzgQA0tCOF5zZ08xtmQ2Fw3nKV7ctnbZaq5mbgqVwHJXU5pPT0
t2UaffqBKrOOZ647RewekHoQQUjnFisyx7gFQdknmXJWRfeUilqkuhy0UPdw4dIAQpugJLbD6KfK
AmkPniD/WE5YkQsO8FoGxP5DIilIwAo6ZPwF0qOZXnYFOil0wUU4dQinmUiX3OQ8yGpjWcdTsYOd
40ZbiCv1TreBYlzh4SOhKl4l3wM5p93gxCaeathfVtd2hAv0rWXcrDuGjrHRWke6vgxWl9LO+naU
QpvdZ/7IMfHjiROqj50dfUr9ESLsVyX+liqHRaIr0nKw8U4B0ox7u3vn4DvdUdCkFF7Dvce6ze0u
y2V+a/mPDvfUo/zWEmDLS/X41F1kQx4Ip3f5DV4V/kZKVdVNRh+ShPa4vgdgYrR19o4oQNkt/Ahn
VLCL/Gm5jyrcGNdmYqNQ9OEJnjyY3iJatviaHj3vmo7p7SOLNU3lMZxelv/+YlK1dzzsXK2nZdtu
oeDOK1pjVZlgS4KyaSVvkgX3x2KohwQDn9aUZQgzDC6BAoiwBwhKtgDyTTiqLVr26Do3MEHFkGTl
EMP0uKCw7H48rbiRydOiyOU3uYpxLMCSZY2Mpi2ljrQ6Kh8ff+eLIUbyM2w4trUb1Ubk4MB3YtmW
JAHtTbGtiucBh/7qNzqULrjzjf+qTAZCgPS5iBoBwa/SZtdHQuhmPGO/x/7oCe6e/bvSBqPoh4Zn
LnqDw8L9kBgyhRqwYAD+qKckXpHGL+syXWEbHXnwOMxU6yjRg2WVqUAahKu+Cb1Rb5tAZ9skETG2
5Flmpx5tlb9TSDYjhxwxbgCz2rIaJJndRZV22wBp5Q/gpfprU9n+hkRJyfOotHNu+vqsQAfdUSUe
5Vw3ynIhxlSdRDLQYVIZZGHNjlPfxha3M9p/MW1zhLFo2tbPT9C6QTEMdLtKofY4FKkGORMTVek5
7daj+lPBgDRYEzSf1psqB+X51L388xkM+guWvm0rulySPwjEGfF1qVHI7ccYqqsJLzSkKsdno18A
jBJDFNaJ8yKux/ST2JJpsDb0iUrN3bY6h1zsOfzvvmSxs7GvWY6Uwjp0QPOMMr3gHAMZQuQHill1
vPyTCtteSGb5j13xgEvutYsK+ylYWa7EXs3M/0N5vpQVoXizVVtZuvHImlVH2i1k5YNtsQ3hIQHI
3TpdXcHHYNmGOQNyPtTptdMeTdkGfrNnZLNvh/lO4qjO9CKmtxDs9abd8apusrwnbFBed5YH+99g
K1+9anEJ3xaUv8ddVQfdHogRQ/XVH4Xenvo9kSQs0Z1dURujnQxlzuogtwsb5g0hIDrOv/moVLE6
MhR9p6x8TI1qQORh7ZtQPFOB5hkGSupmN1qmxp95rvYkCoBXAHG4u5hZ4eZ5sQMQZatnPAufNO29
RMs2alCW9sPjdsqR9LajfOMEhWKcHZZG7gtTkYcP1ysq1tojcWDd73IYrsZ3t4xX3FUqA21GXpuk
k/5j7xh6BllNQmKaQiCju8TmteGleQPfBJ/Z73arsWyI4Y0mj707SpW5dFnYPppv4DMpTpUCUgu8
hlwK5BNuF5+WYU7L4wMwVwlQDZmvEKGWQJVmz1+zQz8iU+xNra4g5mEKSAD5HFpgNMRKDDt/J2QX
tq+Rc+awEOC+A1U7KK3JA9iEVVQIZgQ1x1OoQvU+Ms4r7MDXKr69mT9fxhXxTiMWX1npptwXvsDE
+KqFV2ovCU3EwLuQhnVnLxfw+DY/M8OUyf3iFQgLN1fVJPNgROfzg1dMj5pO4raDmqX71BxAgVKx
cb3qBhUyRNbZgQvgz3aXYIMhFHyfDsCDxBOBE5xsD+xAAwF2cHlcfqqA8ivrYQss0PP6xnmUoruB
8wKFQy2F6K74k6RG4pyTBxNtj5RiYQH7uitMKLpzlrWhA9Wwq8siezfRBmaVqb03L0Es5uvJht23
HrgetA+YbiwZY/ydQRd0S8yWxHrDyfula9FOrkWnHMyBZ8ALCZmRcZtxlG/tFKQzxrZ4fNTeJ+Nl
UOV7bqyQfFvHxXfM0Lq3whWHO4yuCnKz8RPDRH4SyTjPstfFg9uzmeqU1CKqFSR42DSYBfOUOFNH
Fx0vKmQoywP/ro3QroauPK9i+CORdRHSp3tL5SGbFpQF8D9wDLCZASXPTYZP7VW8JWrokkb6Gtye
/WLbhViPjhGNN/1JLyQhYn/NTuuL1cD5lfvi1/Lzu89yQ54NIc5UgrKl1gJICIokazlkVd35gT/2
S7muei4RwRtpYsV+rDYKY3M8jFZI8GieZAJOCHyvpVxJarU7Wud3TDhuvVuVsXd1eV5yoHiwy54e
GqymQCTt9qMpaL+/MX7XmWssoT/h9hLIO/OV3d3hPDzPCCnQ1FQLyJFQyB5v1rlxbK1547QU1r+A
sKbU8L3D/7EYzp3cHx/ZLjBBMCxZRa2yiT0eNaRmSjwjEfrCz6TbEKDzHOBq9k4QJX9Z2oZ9y5J0
2FTfF+r4ycyq0nKIGzsFZ/lx/M1leH3ocjqHt2RNZt9wuBTVL5cHGw09+bjfxebkQ4557u0fUBzl
n2UrmH1LpTkjXyo++0xv/Nnip0lUZ/6ZLywYmd/smGJQNflHM1X39BWDrb3LysniUgLhGbD6L/Iy
dIWHIgl5N/4BjWpkRpNRuDOpmzBi+1D75xbIfVrrUGB4x+UKYiQ6ErWPHN+trF7vJuBKDTobglML
9tihA0BOPt6O6evMMP7FZ6hawI1Jl0gXVESJHb39lFT2POvbFjcxenHkLRsnznLhkyzP4Hmha/EM
qugXCpRetEMgIvsbh82g5G4KzGFjeJmq+OZDYg9Xqcnm/1jldSeXcb4O+IwsL+2kiWawsuCoc2/b
/LgUSdYwN5fpA5N00R7OtfMI+cnfitpQ7yH0DVjtbEXWnVVHrYcxjJMGBRCBNwvqhIw8qLCjHWmR
jO/CbTCoKUc4hPmNi9Cg+ovqfs2I6X0u7WD8oKPmYG54/DJq1TURIPjNqlMTkdFZbEVZZcv/mbLu
azsqbcK0xUKHAirOo2cUfZ3CdDu/uVUnzlvkdqYAsk8orRDYmOFg7O4ozUQEgwUsOxeqaEWsyLzn
p+LKs91JQtDgHXEcw4Or0Ey3d+v9e2RUkhpZoEgCgapGAkQYWsITZZf4umy4mEIdinq8vdu2G36Y
imqyoCWUHJ9wMFXtc5peVIfDU/oGiAXqPzGPUmP/SAi3CWwzgwPuWko1T61pkHal2dA8QBLKSOS9
+f3ZnGh9TDPcwC17XNZiebbbG+W/jj9UKebzo5/KaO5lIGWDwNSJiNRP93eR0vsBSIkKTwowkWA4
vW2RyiJP6PoXjUpfPEVo8Gbib4QBERAuPedhbMGlZV11zcJ/k47bM4Ezav1/Tzqf3SKU4JmoqVys
kwk4IX4SZV/fnD5FRpshPiGQpYZooiwG291vY44lPnnXA21jYJbLQWgwh3hhUEA7FpnFd/eMok9D
IiRBvvwRe47jP7LK0qIk6+0EZcH2PYzxfUdbljoj9D882+mIkXCloS1SpIwbAGaslVRY3YarigTR
ewbZDHeKrTN/DQb9piJdZHwnqB2QR26CA1wkbdhSF16K/tQApd259qRsXywkS4f2iTfAA3lowOxW
DvDtBnDKk5dm9NoxPo/WQoe9JXWJ930k4/v3a0GE8r/lP0R1BUGIaIgoE6ZRpvnIYRAd0r/Zo01/
xl7VvFTaB53W1xPnvL3/tN+KMwI8i180cnch1LZ16AQdcjjt6VDHPdHL3j1UfqJ8euNg7Z/X4FAI
y62TS/rhIXxVAi+XANotoFg7yESsbGlr4z2p8hR96WuE2+ll77vjkVZ/3dhKWlDAQH0eBjqMPQKt
NammvjkfF7GgGSMzxNc4S6VShLSWAN7RgK5jAp8+LG+B+CPltpgoxuYOMioO66TPmbRC8P6euXI9
YNDImW+Xm3z70C4aEZ1gHxIOfP2lwLYi9MTWViGjFC7HYSLWc6CfNbvUipcjnhN8FZsmB2d0ajGJ
8rIAd/6Zb3Lh6gKwUjnsONpytvH7dSR/+MCL07iby+P1UYRrwljPWxCw3jA3hrvVFK978BWQ3BKp
+u9B6Asr5EmE4Ggj2txQYHTyg6aXiXFRmhHzguL2Gnhc6ISgxysSb+qqAlcdnA2ST6KFe/hKI/Z+
b2JdWsKMxhib0ukeLbu1rCQ/S0kGUbcb5eTgt+SyjIzcMc5Tqq2DTq7xZDBMN7sM5BNSn8XXwJnF
XdEo1zazB62dpmd4YON/qrB23iB4r0uytK0LOPa7zC1qO+G7mUUcjGVwF0DJHDB1Xq32mUks/zon
T6419LxcegVNfRmmjYV8BAlkTlyXKymyk5c9pXbgofRlQIXFzve5TbOy5fLNCaWj9dfsSdIR8Poh
iV0VgL00IvDfxbQXIYZ9xn77opQBcjUHXZacpnX7Gsmsozs5ZF9k/EBFnfV6bw+WRLFb7GcRnG2i
ztGm0qtiCZjXFH7BvNzNsJNpPSlaDG6pcFyOh1flAeigg6EZKcSqk99W5eHaAe66Vxak5YqP/73T
eI+IfROLy5oopcuZAf+nh7XjqJEUbEf+OfwXO3FzxRH4VanT4TIU6TiCpa3lL91XIM+n4EvXCUsF
9o/xlaIJFzXaoCxpioUur3jfWwFC/pqdM5rKOxd2ixdL6z8vd/3XiyLwxkKl1Gi7UpOaXGAYhJEI
NmYG4yUeSuO+RvS4PjMqJAZPzS9ZNl2wIO0dm+irj4Su/dcyWnBb8/nC6XO3PGWOgI9ANjatAYDj
7HoXfgOUsNWX52J3GoyHHkk8ftlho0VSWsnPRTEX/U1jgBVMzm8lQD+c4CrGCcWIhkFLafTd9aXJ
nUEKI/W8JHp1qv9+PL1/Jw/yAJJqTq4+/25JI8easPwzW66MPs7Ib/QX6OxtO0ksOGTY4NzVp6rA
3ZxR2EJ87dLEzOcIReyJVLxdB2ba+8CfCtYSjNvPAYghuYCsVce1HeKtDYJ+Yky/+uulIsLD3xQ8
/tYxz1JNTHhB913KtaRddzT1+jbMe2/2/bS80SeWc2heMGAW37XK+BFaA2k3LaK+rWRg8pM8Kbb3
UOewR/7JQvGUOP1h9mcOTH0oHFOpPz/0RBKHGtjlms/Tdcmy7NiF3Ehpqr1sCWrIJvuCon6PVaxh
4Kcn9A6VpyaqQ/sFC5QSttZdYfjBs4mzoSiO+95MnVkMAXxz8QwEoekoY1SB4z8vzg1u9De/5cj1
30ZP+BZ61zPxrhV7vdKbnJfLElAhkZBMnvEK3P/xtnYKLRtY7a7/LgZ6fbDiUOn6W11VV86vEY0i
ci3KbL69jCPQq80CD1ajUhxcgLRS0iWqLADs//F/gPFYtx24nuulcY7/pA6DTzlTAAHAHXdip7z6
BPX41DZQnDmKZ7u9Ji1hzsY+anccTEYGlCyzILjWmUBALjXMn2X0eVjlg5kUo9Xgl+zppCAELGnK
AFChkqLshYZbcgGv17kJaJaljJv4/4nCRgHp5u4plEzuhkkmR7jAya7BFCh4mVj2/45kmyrfw55L
D4yEtXfY61TXtcT/U3hZbyjFS+IkeWTmR1LeKlNFD3aGo726/TNDswTK634yZH4D631Xa8+2P0+I
zc2eF2gCdQPHba1hunBSGc+RXIqAhjeBgZ4cCTrkCnRKDYaPXN4N085ZXmzv38TtIzI2dfEc7XmE
3Ie8dW9V+KGsTq1bgEhLLaaB0XOE3os0xfcRrIBH8J4sBJ8/Kua+er9wmnnlqi4ZVU6ced5xrGDE
RddRWdbcGMoWCtrXaFzK2NWqz2eB8UhfKdD6fZKeqQ0cOsJocmCrpKrCuVIya6Q0lHGnZEV+PFFs
JBGlNolYNgQpF6gpQCcxznln8dHG4Dhj4CgZLBlzSBpnd0JGYfrpWrCbn5txkQF+n/wKhhGtYBT9
SHzUdot6bDNgWg6u3yjNzK4eT10OwrBcWsySDvfugpzPfk8V7fbBerZoITQp1qHQdlxZQ/QaX98c
R1lU3Ot+ZJEAzsJRsfQeL1ChIhC5FoDPpehrJqQles/Jlmvo5w67KTmGaZj8NfrphieI3wwThHBe
PTB5l/WB2MIu8nzUzsTba0MIB5grs8e+CP7GdsJi445PmHybflktFTVQiPVGIYlHNf1o6hP7+5ZG
iYqKE4FCxKLLXEq5q+kuwpK/q1TlabVyCJlBzZsFOWoDgYJO75x3AlfXAAePdY6JLrmvXvDAl3zi
xbqx/FlmelchUlesFd2Q+OFWkgXaJZfqixm3owQgk9ocNSCWDAUmAcw5vC2zGzlpn7WIXCs95n8N
bHDaAa05c5LjE/iwRo5QoARhIwvHEzCHo611ab0s/hEPdfvdUIBEx0UQU08FC7iD5dRUYB7qctVD
5SpM2M/ew50kkCi83dBGrSMO255AIl/el8Aa1M3zKtPA1IP48QVvukdfy6Bt87NguuvhLSaxVs8z
MVusNX6S7L+UGSqJrUm1AsVu6ltLe0Nxr6O3i5D1nP/rz7kR4lGg/CTl1Sc8RUbugjgBXM6f3zOD
hP2aq7cupOENSqa5KXmwfIPFueWo4trUf3L9ocXAd5j0de5nq1D7a9X4LH5wQ+qcxF3UEter6FFj
uyve4IkHoguhW/HkZ7X6285GTHupjwDrUD2Ss0aT8LKuN0eKZG4z+AvDATD4v/IsgJUbIbJksUmF
Vg9tPPP6OhNaLrAzf1rzeCHnCiTJ4i8+R7vAAYih+7bQEi+KddokDrqf9tfA6yynBkVW8sEDWYGc
FuW0vPDgniGiHT9+QHT6V2z7VInelZsTNSp7lJcsE8IYobA/Na2FtoVEIavjCy1xn25HVAJDtKAg
X1D/qJLDCpNuzXs1meAQNiycGOiUktBRw583l+1cxw2hzlt1soCkhnW63yJNVzl6/5GX020ocGvo
7WDy+pXX6wlwi645d1vnoE6NBHdEp9Wb1AEEcPJ541IPSTLTn+GZfU+V8h2aCJzrd5SVahoX3oZf
7RIHtOiEM+sgttvNAMaMtJb7S6U/QQ1ad5MDEvQ//aanJjonQG8oXiFpDDVIfJIexStvkdX8m6OM
h1/Zv9qlbIUjk82aPV0h5whx+mVWlC3gOVR/Fi3bw1FQFYSWqXZ9kzD66rJC+BIQeBQHTttfVemI
Kk7jNBN8qglxG568YppQVBTpbXnqpRcpYA6+G4SSkFmc9dwP8OSOwBWveBgEafn20oMFsmHq3lrf
8JPN/KsRnptzrK09xRqhF7JB9eJpKB9StzRsBj3BpmhJl5Xx1FM0LZ/NDU/0sZENVi7LqNlEMKP2
sUx4o39XuO0ndZN4ylPO8cCZ/fUJD71shkRJlDQ1srdCUKQo0FX3AKGxpGTVkHcCYPIFeSnu4rK4
n643htbh55tyeNjQ/EOOJYD3LhPQBeHsJxvjZnozsdE/MS+Gacj1iQC+nGyG4iTPOyVgjBwV9Jyi
RKspgwHHl227zFmfjpic8ks5Knk6sEhXIYOYtzfCWE5Ig7iJk7j6QKt/F3gzdvajLFHxgNsX4utg
rR7OD0JeBkb+JxnpQYkwPjKfoMr5AFaB+tY5d+FvMtBcag5cN5yn+3jkDc16YUpr5F0Y4gnQGVI1
NrurznJYOJKgqR61XbL1Hm+GAVDIUY/qaa2a7DbgfeBLlcPUAjsQK64N1sFCS+vIXth3F863SzT4
uRxaPtKSfpzE0NzzIWURHAaEQjP5kPDqYq1oYDk/YTuTBWuCc9uZEaFoUeRgVtwmG0fbmPG333nC
/D1gib0YhGEaz6uNYX2E+BTgA2702XmTsJmwBUSVHGxzgOIjL6y5IAepeozJ6+a2KyvUjabgMYW1
icX/zjPp/AvtNVF+GnJj9vgETwXUZh+EtThTzjn4e9mG8Fu61sBKf2D72pilO30/s8S3n1jb2g7W
ixK+dbC+Jtt20f+sqG5vs3sOIBfQCbmnK6LG80o9ZPbvhs8l4A8uEH6mTZhPX7ehahfIdXWbciBd
GO92EmYqKEvBbnBPnfYBgQrQoimy8PToAsI3088gdLsBiKzGcYljT9TDYyEkLYleRjl1JXkV016g
DopixN/bgug+LO4Jw3t30nuwRM1PZp4ZCryX5r+clNQCz4wa0YRVV92bFOBHzCd0Pg7/r3zQy3Nl
izb78mVjauXdfbLT+HxSr2yWkO75D9AEG8bPVM3LJQSsjzibAuHTchCMnLyo7J89BKesM37w+n/S
3wjg1fxORV3VqoCqRZdilOrC1Y/RBXh0UOfW7iZgoz1KveSA8Aq064ixaIUBD/cqbhyT4fdiMzS6
KI9eHsbLf5OWjd1WOxrFMPwurnCXUss5Yp8DggLPYRH1IeqOFz7QBE7H9n05/tukMJGy9wB2IDxu
cgMBrMZkPt3T7Qtt7ODGXJShg1K0mzAHCZXXqXHFRBeswcfB6F3ASTR+yBXDtbQTsup928VQHgNy
qipYbGGGnuixg8TGA/NHyvl1OTG6BYfHwC/csgqcWYCMCtEF4qSZNLmzj7rqBDLRN3b1HLxPSOn0
mQr1kJZMmjaXo5tck1wJIAMIztwm7CLSIcFAkxtthr6bj3ikmGtHj2C6kUqVk+ZWPhkC2dkXysq4
8qnUEn1ygXFqnMDotsfJvYSdLyTp8vOUM4ESwIAcSne1X3ocGXekkmo2TCoheZr+DQ+y+NIjXCib
0xSo6QCsv8ty1XBgIgj8v5lQ3zycVd+YL9r25+ZfyEWhQuCUHCRW8alCd1pORtnEVZesAo4TIe3V
cUJq/yN51XzLe8UFrCqyYbPFkh/wwZXhgV1k5VE/iJYt8shGlvIy23g3426H/4MJH0+ms1enizyc
7e48+02KzduIFTpxuNMpM+GUsA3VVhG7OpTuWO2SHsrtbZf5dKaVpJ8uIPZNxWyTNV6+FIFFqX1h
HSrNtuS863WYciZQi/3W6DemmhOjBlG99LWC/8Jdr1ORUuWFhexU1aCkgnMkiy7MxHJ1rde66XXp
E2yJuY+0icgn1E8W7jKlJvoqVa+DjqhikKvF4LRS8bSdcRJAmnNPrOm7fikIS2ocLN2FKUtKIX6X
mYXMyWHGUvC66UQ/ik8sH9Z388SB4P58oZaFRD+gPfdGNzFodlSuGzktU5c/dsuLCwyvkvZVL9//
1HnavERePEtkHF++r5I+T5HmBxuIrC6iZpOayesT45lFF8DZ6/tK7w/Vvyhl/fleEtebEh2PInax
p1rYP/7A3VCkT9J3t8SvYn34QfTQPfH95HO5/pSOsmsx4xLwpvrdHP3AcRPTtkqG79xKl4Zh5uZr
gY9WkDSBsogqAMnOqBB5sveccku8U+w6Tp9gntKBXrF5MWnKFYD/6b6PrMbT3Gu1XOwOVrthuAuu
cd10aDLwhGoKQhcvN49yk+j1HcmPi19wvMcNqkndzmUMAC32/pkDSeSTpwBmzv07f1tZv8A9Os5q
v16YBvea8CmuvXJU7sjbdaNEStVMkjuLObv4hg0RLt4afc2UKhAvzP7nvlu0fFztSBCHMVEx5VEE
cK8dnLrUOFRhX1AYhzycJ0CCbCMz5MeOPpbSQokNwdLQ6lALy4khAbxsnLUbx2lO0xroJCZyLR98
vadt/jrbRDmElAX/Hj5lZ40UyhReTFqZGWQfdW2fmql6wMP/pkkwbFw/bZt1YdknEAwa2zoa6coo
869KH4bdpTc8dOC4t9US94jpnOpD7a8Hnp68d96voPbuDWKI1jvkIlKham8V04S5SIeqzC7/Zo0m
ONQqSVMS0sRK5rSya2OR6+syZlpd4VDbErax1UJlVTqwoARV9ZwYyacLWCRWgWGjI0k0qzN6U3kC
z45FskvMgHM+MNDdirO9piGtr+YuRK3AxuNqIvnfs7oON17L7K9t0m3gmqu3ddgzBtcVuCBZn7BO
xCO2+r27jEPpI2NypO6gtrn6vAbwKDV+YZ0wJpvoKCUxeg/aC3yDiXnFcw7JxhOdePQnb6yHPkOE
SmC8Z6mdQQjCOSPp6Rza0fopbsJ017mkFSBbKa1t5rjNejN9A2fqsAw8ZN/0hWeta5xBMJQeetoq
x1KqS9rC8gv8z6KYNehxtWUGI64goYarKL5bo3J3QjeQTD8DhxvecPfq1X4vhrb/JTa8zvHbB9hN
ArsEqI0ehYLuJ8tzKeDLEtto3dyqsXLQu1Om2bc8wpX5XBbVEOpJ+09KN1Q4Qau04VT+Q3IIAdLc
2Fwi5lO2e2JiowB6CUwBLyyPdhlwXXwIuAUeVEW/CkNE2h3uCiXotC3nfWFAEKE8lbbKwE/gA5kA
69wr7C7cSRWORmTFdSy81eHE+9X/LDe+xiAGX/ngOQmPzTjO2yvAD4ailAID/Pxgtngl7OXx5xBX
TDAt7dAG1VUlmdNZOkpLKMZ/T4wSlrfvG+fSn4/NwxasCRPMG9yNyuPHBf74h0qg9aVYYVckKQcr
eCMb52lRRW+4bLokEbWY8AYS6bAf9jKqlPxIk5VRkFN6coKJetJk38a5sAB81QRvIbdE84CWtxtZ
scdk2LTDWshxe7ZLsCKdKA6lz/AxqGRNV6jcSgBZ5P+LfHXhIMFsG8Dh30pB3KKGCkp18+7vEsDF
zJf/bYRODABUbjwuyfRd/RdylhgaO2IRxe+T6vcIasPpDZ18FvNLZfL5ICjST0o8MTs1KaM/Dnhw
xyF9sxGIYGSdfq/UGDaIWOadmBJxZh/ANF4iFWyUpCYmewX/ZqJh5XJ5F71aeFZYwaGVFO8c/sNM
LcYDv2ub6N+Ua5lNy+d/rHfS+ZnErOYpVGw2Sxha9wq1NYKukTlPjOMO8W3mexaBNZ8aIuqZLPT8
PSXtHbFTGPtSSnsrrJvdLddZLZVY/TdjWxWtOf3J82rLaDaqp4xoy+OovKO32y4cmI88iVGukdAb
uKKSUUiUNHAVbMDZrTnZgBnrSR402pdf7G/2gCHVI0zp1vWMjcJ1xnWrBAtY1glxMEmzS8rAeieC
rU4V2HoEZjILHZIcDgW1jXHU/mNxgDGhXYetamDRAoz4i4WuV1RMkM8+74wV1bhMCI0Vsql25PTH
n3t3HQPh8xK4c3To8VbZ/7YN5pkS4wYGZdl+afgK5rrtUr8haZZb9HC1PHvgcfkIBze15XP7IOtA
b1Dd9w6UOrH+BNL/OaWCz9uzPgTh1uuamKa3+u6wJysFvSkOJiual27edCMKdWlJREo4EXI9ET3b
WFdWJ8E4fAj+7Dt8ZyJ5bFHoHfCT4uB4kP2iPiSjww03143UG8cRqQ+Pty2xRgmnm6UWZaD3NVI2
eyXQgRvPB8EV/Ah8o7z9WzDa45e7pz6DWY43F9pL6ISICTWM0lWP5z5o/ZYix7QM+5DJ3JDLb2d3
fH2OWG4MR2A15cf5SfjYx6Ag8tDfQroO4MUnANNfQTvSD0+K4V8dbKR0/FRUQc1Cn92Z+3QyyZKh
cVQMu11cqwoaUaTRXwLcrX1utmicT9t3XA/lhrpmwWAG8R07iclkv9Twp+sZE954jePtJTbZmcah
OKdTRYwN7zBB3o+XqgORxe9JreU61oC6aOR+ymnAEid678oye7wgi7h2Hj01MIjbjK3EEbE0OzNj
f8tGF1nNccoRUkn6niPQS+Ra1NAzORwoXd8h479fhzs5CoUFr1vJmbrRUieF61ukNVzvw1BsV1tT
mg7vq/HI/inUjv+jPlX86FLudbyPAMgVJz2lflNu4QCzClelX+mtDsgkKzg8DditJRDxEEJO2g4P
rtRtHE4w9cARVQuCjawLO87PrNrxxTDnlqIpqRK/RmFm/jo3y/ljIf8VtEzAhPd8eYEf6RCrDlLP
vlEYnr7n/LRCN34at2arGO7rZz+sfYa9v9sIa7iwoOE/9Qn7XxOC1Lt6urFpAAmN83OwAljl2K5s
Gv9IWZ8z9OGc9ruF1tbXstvOLEaGyTMLP9colm9u7JojgmdDmoonhjhDHJ9Ok7ZHjSokmjdVtVAa
/nfC8FMlblQkmUwZqf7SQ9MK2KttwnWRkQ+J+dZPEe30MYTNLE1hfWDL5PPiRzueGL+b2ipi/ex8
+wze4qu2XhlsTOJx9CfTdN1tUToyYFrDtLDzzzxUGvFKLhlDJ6YPTZfzinPRSi4Rutr3mhE5RGUy
6GTlytwihQ7uqebTFTkLlsH7x5mxUv05TdtzH4WQuWaabdeKZUgU6+8tkIQFBOaAtSvxpDcufWHc
FNjjGIlKV2wEDJzSApTMlp877ZqrsJ6II7vds2pKNW9oAm/p3oos4OTlsYALGGRvpPjF+zmn+mjP
RMbHP5S9ct3kbCmIv+pzNzuz624OEgzgRa/NcFDD7C99Ah0yeb8cbciQLPwYXjAwwBLuwyKKRmRt
IyD09YQYFoOxVnI/Mo+wQVGgs0az3pymG828S2w5Jn9lqEXT0GacfPb6HyAhpqioGnlVdFQIGB+j
r50lYtPNswT203wtlbdit4b7ZLOetWwqpVykWUdEOzYiUNbvYn84DlBIxHK7dT2B7fbZHGWuEBsi
pS9CXrpjx+yIttlhvLxzjgmP3zcdQ5UL6sPZ1o8d8o2ZDGwCv4iRYUMfc4Udc/z2kMRRr5Ez/WbS
c4PQ2HxGHLPhaWd1Uyw4Zy1e24MKgGvvOFR/ULhQZzhlcj70oq4pGi90M3npMzzMm8XCIQEmLy8X
eefWg1FLPN924b+JkOi+1FFjHWY1E2TYF+wHg3jIkrD+2n/V0mglyvV4oQEiXIHjNJCpsAsDOtbw
Zq04id4xK9OCXbVBGdqOXO4r7z4qLDTaHPnuYiTtrcVTc78bWpeCXu5CzEot4AodCgx25qxlm4We
nc9HvY5z+Zcy+3VX5E1/HUNFm7vZtkyAHq5VGNfUTXgwqodxHaS/V/ZRPRggCkLrOiFvv34hAv4G
5CAzy6ZCp+6xOj88LZ6RgSDxw56YeoH4KDqH0YQiXSmooqqPEwLOqJ/nsqsHuLGW7jGxugZrlu06
wigJb5IFP9nvBhCO4jMrqiTC9MWo/uSZhq0u+XoTXM4M42IzsTvQpvvrtBt2uASu61VopwVAoHDh
+um6C1pJH7oKphuWh7cQj8JZi8q7n4TCD2PUnumR8lZBasGs6iIxK2kIzAQoL5/EmfMYoMEJs403
DwW9lIcT1M3RIjAPIEEQNU6p9wxi8VYmDcrQZ+Vp5VGce6LiohN7YvgdrHQcRQ73Pb+n7ZQgbzj9
327NjOXY57Il025hnBRM/WfVCNPiQZC9mBQZe3drc3++ODtfSqI+7JPArgwUHy0NXD042Q3l4jZ/
PjaE+cYNfA0WGTWXlH6sYKk4/dBj/yrvA+4XoQmXTs8dplxddPrpjaoBQQJfx8shachvOLBI8TcW
uvnFNLrlQoV9qxc88ePNpsjarAvUcnRRxxO9rMGqwtH7gFVT6qO/qLsopr54U9pRWPWcFgLXW4Om
YUY0Kj6rWJmsZLwN69o0b6WgwEeKUyGYdE8F1nGkBqInzDl63fs5kd3K2jjhvPw2+GnG33zY5L27
pxU3+izYAj/p6XRayc3UQmfHrl5iv13WQQGVIF1mYJ8AQmFobiIKDDzvS+xNZA1UEBzaRvYeQaJw
VvCpWgTnjl6yPwR25N1WRKKDBG3n5EmQM9fYSZVFvz6ONO1i4GC0DgHyJZHmyTMU2XwDBIMLF2D5
DlbyfW7lxHMvioElTTUlfyrF011Ww/iM0FkrBTvmkadzUkatOt7Eai7/SZNoLA9XW182Bxbe9BM8
UmLoIJgOSx1kETqgsLxxKxgEkA12yAwob6iO4wRd2T+bV/EGdgq+GVhXdqEw324AjalqaBiGzzTN
z/fTTQrXpd3rloFr4SH7USg8UkzKy/aaIf5SYafx98U0D9bLPwDoJ11gr/j0hWR6cbtejPCn+RTQ
B8njcbVYCbrh9hr+LIej7y/0kue5QidQlPHHQb66rZJCOziTMd7b2w/HqvBkMGBJiJr0IlJt9rfc
yXzv3+vO3445D932tjMSYl437en2kSMqICd2TPmqIar+DHpRtxXrkFj3Fw9RD1s/om2uqKJ/ndOl
zWn6CugdCmkBchbNk4kopvvrV19jJn3jcHLuNOs71nq23fvIeSMsRkW8ylXNG3bjOFscaBD9uQ/y
OI0mE+jgGyxWeiNbAcCbutavDq0+mUE+sHNnmPo+MnrZc7qp4z02fh7kmDdA279yWgb8BRFG5Kg6
j5B3/Z7J9QjdZMjFtCBtY78SzpFwpMXwz+H4AXF7yUdYX4IRKeewPqVlJVdQWLlO60RGgh4Dlnau
odfHBbE55qZQ5KXo3gW/1VLHp9Rxbh5TZz8UPRkACPUMiEi3CRBbNxalliRtGbS5AbbYz47+XsIp
K66/z37iJ/L6kRCTNoVpsxJkiIRehbkfLBZqnT84oWUA6oq0yD7NF3e0FBWo6QM5GrEhbXbMQCEZ
8MzZSr8F2uFQhMeQT+7OJ6l4VfAN6ObMKhZ0nS+4GxG5EvlqwaCVkMVHl2+9lYjys1RpJSbWzsNf
rKU6DD84T/qh2/ivUJ/NMG2Sgpodt5aqc39c0xLyGK5jiBh1pVFYFRgfk3KNnXcM1mAPWZsG8UB7
4LmAIEVHK9kFB+/+1brXiOUymoE5F/0wQCxvBrlR0QdjWxpgZfKB9tvEP//0ZUi59EN3p3wkEjlS
6ZmOfkd999HniNfvx6mAsb7NSdoVgw9pd+J/YxCHT/FrqWUvV6JRzSOrOd9KJqPdaN7thm70VTcX
+Vu7ogK8Wgbh7p4PgdupJ19Od7oIDACnj0IshiZrw8hQ9gwLxb470gw5eok4WZontgnZqvmKzscE
jBL5ZWeiWRe3gM9BlI+J4nmxjFYS6kwWZWpA/GewE/1iX8+vJ3whxL9DqeHkQXdIv3sgPZNOhrHA
NDOCNXRjQ1o+U2F+iTV1P1VesICOvG5IP6Fxw8/ETGFppFDZEVBWnaIkEljMceX4GcZcOjj1dWrS
lW3+4SX768OGF+sF9b4skjdS1/y0mjSSj12s89mDyCidx8MA61BiGap0dcQcajjkTq/QqqxCKUtC
VKaskg38LKTHhLDUPYF2fVIlixwdzlpIoqAKcSAsS3lirj3GqGZpvcg8aXJECE4Y58UeAVolXGWj
fjM8k5Wz2U8k5te5+dnRkyMweiJ8py7oJ48NnaqS87Nfo9CgwVwgCwyOXYEhDeAJ2ecc7SjqL4d+
fUGz71Kq/w1SF7TLLRPsZuMlvHErETYxp5ngQTtk+qh2ewORqlW16rNzpCvLqbcfNj8SkbCGTjHl
kEiRKZrqcINqc9cYWJoV89+BpDkqxM5DsF1WnF10tqKKq1qIkFU4U2UyvO3C9FXHigvHIVU4AfFl
vIP4udDnGq3aPOVNaI5kklHsN0tAEG95Fh0ZgrJkvbQvUq5Ynqea0iYOIS/4hiY6IlGuYcrg/9MF
bRQZBmrBRFWXurqvJ2GGkGz78W7Ld3V8hDuslcZdYtmSdF1C3qAxy+56Ws95PeUWnEHsaAySrarz
UKjzU6yraAUnG3Z9eOzGMB/8rtbd3qHcYK+sKoCo093Bxtd0HDaZNHVRkaX/gFL3ilVCjfYgupRN
iChXPZHxfnjFw8Lmd93eWELdPM23UG3Zksa0cPq4LqtLdZZYu32tZGztYDB6BgxYkoMHWLmgthK4
mqKbaauoqqxzJUt109zWSoAJ0BaATELQKCYGGc54wz8H3zRP4xHMOw5da58W2OGBvv1vqU8NS0Jy
ZCSkxDleRHM9zsbmsPLQ1dA5caYJJS4YKbVL20ztp7i/7MecaMPtyOobwFKsdsKYuKIjzYQ/m/hf
0K0XTbcHX60yx5QVT+xtuYrMdVZtltG4tfctK4o8oqhsKpR7wigpshTUGThIk7m9CqBwPVjugW1W
YinRwAiEze8b2yoZ7bnjJ07R8ohyp2ZukOTMqQC7N5b8TDmVeyBP/fMaszT2EKltj1N8UyeUHYzZ
SC6V2wWmGXQsUpf+RORcn2s+gJ+RzAhnj8HRFHRMilehN07h6KD/Mc0cGCf77eZRDRadxaBlBL1M
4EHVCbU+VXCX6p17URYCIpck4PqKA+cXUTgYbaymxbCoQlmXo5T29fleOmZ4/+m0nAGK6SBE6kUB
JTG1yDCcAfQXPICPRj9GcZaThcdvSDNm1njMedyiNfcRM8Bz2ZNdVfyb5eXMlimiL6qzBHOx4xoc
ux295DBcuwkCmJQ3gmvPL3iUmV2xPferLDO16ip1uilQKUE4VW1dg9EG+6Pe5yR56fY2ACNdQu9h
9mn+7jqZi1oSrQ5YQWEb+C5sxMOBLozTIwN6XLR/yjitU4SHFFdQTunsU007EFGMeCj7jEAEuF6i
auDe2RtccmdgaAk+YS69EyX7pmg33IlVamvXV2VSYEy7K+GS0hQqqaEk1xbKoWBgOy0hFypYA/6d
5rXg76PDeSbf8oIAttRnfST/tdaaQcxe+okNXLvmcgrAibOV/7vBMNGkRBKWYtn+DN2YIJYTkXFO
4YaZbthZIa86IGCPdUSiKQJGbVtkL55YM8zsUdtVHF2VGHUEIDs+uLlPwLLRdmHkP5ZFre1Ai3TO
uzeomuzaG38pOJbUGorYJzY7S5NbKn6GXQlg6jROeeDkw7Y12P0yLAH1tsaFa2dnXwA8Ds7uhwcd
HGP6iocx0q0J/erQBqXLhJDvsHhCFlQqLs4ibTtsRqfX1fwQGsRmW8q0xA/K2IcKZXo1BfQcXYIF
uReW9vilqQbJLgYn5MTuc7YEM7Kpk7QhW6s1YegwFjiyx66v6gKM9hXIlb+PbX0MonYmorlxchI8
CWnXTzJLTofHtwnsf0ipEl82g6ai4l5p2J4HKFL6kqcAODJc/6wrOmTpFkSK0H1bduT7zUdEwHjc
mz6pNzOKwqBLIXrXEUQMC3a2Tn1kZxhQ1fdBt/rvqiVBKn3ymcJF/TH3uACyH+M7HLAYgIgrGaKg
gHII1cecvlok7kMJr0CGiFXv0rJTxZMWO7pafTmdkUgpTmklpuxoK1QGXPlBJ7L1CnyFfRbYwdTy
7tVjJfCW9SQhPVAo7vdr6EOKbgw0oDEd+UpQGafu0l3I4ZBN3NZ3qqVr2QHk6l3a+lzMTYG7U5SW
1jBMPUGg0OU8ZJEV93wMQswMpXQbk1Yt8jfjKGR/7XUq+2vesdEprx/h9kjgv4GWwuMZ2aqpNnC8
j435n/2yD5iBZTWARI/beBeNfV2QBgQC4lo/qkprB6//Zka0WDcIJxp53r8Felhvz5T4TLmqjuuU
fA9MCWAXkT8ureH23QlUTY4MKtsPbmkk390CtnxdNdZ10WfMZsuhvECH4Q/vzL61tijrSvzmNpKI
HWIr2l0mVTHo0OFdUkzvYs6vzqWswzi2GI13Kwix9OSdUAj4awaWZLAO5O2M1jo7VPoCV5dmbkwF
Vh4X1hypsxH77ft9Bgy4zomv9wSJs2F93rLFRhpUBi/gcCuiyXJY5bHL6gOR1THzBeSEbaI7CZaH
14kUI33ygkFtDk/raLa2y2t5SUEZMr4T6AJ3IDJ5k+S98kX6uw1uAjoBD1bic65tAOXIlBmUIKc2
+wMToqK1dNvq0kceZIyZUQU84SZn2/VczOCrx0pzKXdCabcyV6kWvxczZ4dwYjUPmE8nhr/d9edr
9MQyF3x8TTIZ04ufMD+gghyi9+T4L98PPtVMgnfhAOFqhu6NpQNXJ/ZoRy3mvHZjb0Ew7rQwuT4i
UMfhz8McD4ivRuVp7SWliNOEo6+DLxEwdtm+k9ZOZBKdm2KwoFIsud1yy2BSaortgMVg0bPxk59X
emuqHPKMLIW5U8mIuLmWc7DwspW7l8gZUE4eEK5fxcHvNpXt8mzhUnxjoKGO9g018kUSjAa765mg
tJ134i6+vYDfo0Wl3laQgfmU8CpwO9Khw5ixcGKg0yGnKm5q6AG/LC32YMxjkN4TWiVeEqRG0ALI
bvAGT08/Nk+5fXHPsDnhJJ2TVS0RkDYWMAZA6svZDNNq2bcUiGQLoGXO9hurz5O9eSc9KzzCHcfR
KFPJfuQ/fRpULgLAdau6juw8hZL1c3+I3/AloWRSI+fOY2cydsLuIO5rtaaEj0gURJsWsDbwMwjv
cg1uTfaf0T5d9EYkdigc5Ck2cE2kmK6D6xI11qkiQvlIDF+gqnOAaACjjP8SuAyjagBb5nFg+5WH
vQDnw7PLkl9DsqaE60WbcLVGq6lvo9MnhrOSCiac+3iBGlAE8ptHr/PQ16vA6NI+GZ7tLbNaEJte
UJruEtoH5drVkARO+sJFUABHOlfTSsInt034F+Q8DLwWweYjoKaJnA0XgnCBsrUdZsQArc2X7J2F
hIaEp/3yDAtq2Q25MUZWlDWKihJhwdSWyu8dIwZNi+9YbmgLDgMg6SEnWZ4Ilk3996HepqHfBHBk
eDEiCgOPDNLk/DIm8pHDT3EMUbMWBF6YZJ1pf1qymxHn7Eq68Cx53QfteKxiIaRjETSVbTqQ+oLK
Dns/82LmAm1EsposIwP17zLy7XJEAROQR3KKs3GQayKpba+MBYl6eBcOshfYXpAZ5LiAtwXn4ld1
Ofz25BMcOqAuqmAGVQHa2R9tiYrd0tJYRP9/hzay0e9dpyefXEb9J4YgR4RpAWYnJZrQmay4TXD9
tbudgcg084XB7/Vv8FDoKfE7EtWoZY5CjcN6RA4Bq7JnhODkoWfbrpLIy9gZRAl3QpR0pRwNRsCk
In1IE7hs9uCQNnA1+zCqFfZjHCq7HwYULB+EbKpq2J/XmVadx4cJxfIu6LE848R+WXzIfCL6FZtH
GFDgvja8CcB63oxLTgJOiKrLk3o9DO4it3Xvs+JGoBbLQBPmJZ9rFY4hlAHyiehxhT8eBvLoo432
rDvgm1z3mo2v8jh9UVFjIrw3wL93OWkLrN4jklJr1Hss1pRWzolGFZP2sBggiTX9XLewtJQT8vvQ
tZtAyq25nqNzVPU80yLQFdwN3Rfe7ssncRqCz0T4YrkAkCECVJIqf8PiDH5H4MVD6mnJC8rriYzk
iQTxlZdQPjdxFU0rYlpFEKnu6f01HtrrO/VbiLBZ0r4e+tR2elMq6ycBL95MJMItsS8Gx7FLLIap
zg9jKlv8AuR6D1GBbisKxmuS6wLi+BlkZb9acq0AqnkNLJ04R77fFmlo32cnUQDBTt0up6mbyfd9
I/MMYY3z0hLSY/rDwIBHWYXbrGm+u6EmOuasWpf4QAL0k1Fvcd3nrCHQSedNm9B8R6KweJYu//tu
eUEIkxnFdFEioYEjXJpeTcwTq60LJ78ZeX+BICZdZN2g9WTanPKVzFfmtqOIKwX06156BO7acz8F
8OW5v8VJJVTGaC30WP3gX2hGbPSyco3lx9+i+kr6HLos/9pSw0E+mrl+aTihB2aplul+2idZuda3
wJi2eu8JGRhFQNMk1hMmQ0WtGh9bJ0/UJdpeYP1vwkZIxI3xHYXxTwT4yDq09+HHYILDe2ipseVS
WQWeRJnjitVLHmbIHBeifQOA3ebUk3NChqG6KH2hUZf1/pdr/p9zOE3WUjwLUpz297hwT3fRJVKb
b8Kafm0gV9F7Kis44KnJzIIrxxbzykaIDq4I9npYRCNtjrIuZ3rz27punmANO6bFPYrTcFWngY55
B24AknjqAxX9/NCkFAXDRmPOlGWsfimkOtpdExttxB/O/5aNOcrjQsvtp+YD+GaYYbH+Kb/dzdgt
fS+RWzknh02dmzpDQCZBQjMC0INU5LbkCTWDgGmD0moVW4P3Jpl5TRiH8Uj/7FHOirnf6Cbd1cK9
fRAHdNyohGv7SHjJW38MBHg1BlzANaEk6vBBLMNli67TiKsKJ8iassBy2k+1QhRc7yNFQbBFyB0d
COHU8CEsKGzYKD11tdl5C3DXNMu/I8kv8oaWZaTteKcE105yttwi1l3gBVsAOvR6rPUw7uzVKtRe
zIVk3usisKzt/NUFf6LOv0m/8/QWg6/RDJKTuDmuIUcjL74fo1kqcfPIQDWXABT2pMrDZr5i/SyE
X4FJwvSSNAW/zdGwKerRNnUhnUS214+rSN401Ay2Riw2J1zbFG/MdQwcA5Mi2M4rUzzHqlGv23zV
EHARD/JdaBvdhBmSyvb6zyQFdVQfiipfOZ7SpWE5TRL8+1SHbz8VlzgALkgxly9UrD2tvYu0wZNC
rO32c2r0vCOUR2/rR91q/3CMAAFC0ZZL1/jEA+/49az2QGIb3Yb007hcfJq8QRwsqx8o7Zr+N6fa
uV8PdkeZ9psbhVnIvtny4eBP4tHX90cHopxlgcA3s0VrEVgFyBNTw1WoFVB/KHPwtcOm7K23A9wc
EA8k2KKEcsT50Fb0gRYS1I/2Z68ZA4e+Qg85XrElRg7goDNjtc0hNsy0YhcgsP8Akvl65MkHPC+o
5QzQIZlx+JwGFwxJbf6P/D0Wr101krVY4Bl2/Oj7+ZrY4pOtwhyPVDexm9pTHPpZvT5QCXdXWLy3
VS+vdf9p032TqZ71KHnwWMONZxByUhAHgmPuP/hx0WUt9dWdGoltGZAQfn5g53eBy/ssowsVQ9ze
XqwmEB533Od81DUWolM9BypQjVjJMdD8lfT70qLSU40pPDwVsGq/UOryRQ7AEsQxFO72TeufDPb7
TMD61+EDJ0S7lTrUIrHfb2V4bRk1G+u8+zn71vZ9dK5YXh5zrhhZN29di9+8XuF1wBQ2opPfzpak
SHUaJcmqZUcXvXArbU4N5/oiKqOY7yoENQGR04vKFxOu4XY14919of1/Yzxm2LpIp65cDuWb+HXb
1bmMggKZIlRkPYr1MR+Jxhm2RtFpIgo0pBNoOYwY8k6XNa6aVNXUlYz6UjIzmxq2IjlqykP/pRwD
gTELhHLoORLL5guqTgnBlR/o1fvRO5ne3QvohD3oZhaDyxQedk2wGuB9FVu9e88WIrY9cxjZx1Ew
4UMfOiy0Eltd+VO9BmABd3JGthw3QVjCk1pSchk7tqpt+L2q39CoFbrmQ9TuO2OWUIp5xusqi6M8
0KBX6kDZDUe7G8l7V8mc1fAt7jfb2bRlflkBAqMh45rMOXMrQW7NwDBeqBPlEJEVAv5KH6Tqq9qK
rEO8to2XFboDrluXVo8WLjUDmOcDTUSgjN3QkfZ3ssiad/2H4iK1YcP6h4UDpykScY6ViQpGTwhE
+fd1/dS7KSC0T9mmWuJucna5nZkCgc6I4q4pIWJCwKt+gVoay61SnqJs0BT84mlMZ67J2vPmI9j+
2izcMW1ZCCSXy9xdJEFpYJGl2duqEcygQ34HWBIHJPVNZ7cNgb/UJZl35RHyDuQcVajW6e2edzL2
Wa0yIw7wE0IHAGEitiqasl9COAdxIAQrX50j3hnxfuvUKxlmbZEz9S1XGayM/EqM3qEztIAI9db9
c7w9eNzkpVHARvOKwa8siO3PR/piB79uWgq2XosVoKUeAraPxeN4dZWJ8PJei6pT/a3jbCw6m8K2
sTXdZDHHxc9aQsVd7Zjj+hraypBX7c7EOmul2mbfiAvZqdP6h4KTSOmNztzZlo7Z89V7d64tRBWH
G2j7Qxvy5IBnG+xKkjrB39aX5zGPtNsKEnVx4BkFCC0rz3+BMExr2jSBcWTc+fvBW1QK/7sPROcw
uwSm5di8tAppVKOG2lXCPuAM7Dv4yQj5rsiNMdIDlrzyIcr2ZC3wrMF0G1yPJlAV63WzWHUWmibA
bZO4YS6pIoJSKInUuEOEScLrkidG3s3l6sl4sogGwIqsWpWhJATWxwDjsA+aeivMle9jtBdXGDse
dSmClytfj+nXBb18dVwgnxb6VnQyqVXbhwbURni2BImqlJIT1WxSxPxigz/5pFZywCkDawgocTuj
IG76tineJ3CwTYgc0t/IubwzNCX7i6mwwpCUYM2NxHKsf81+QdORdVLAJPGDPkjRM2xK+zr1Qkxm
QULw/AuE68hLI24lIBq1TvqjqO9P+X2QIqttC3HxKeg1Ch/0cGGGOQ/0CUdvKNfF2bwXFJbCnHVt
i+1V5OU+GKeNv9tQAwvrQ2jMKRm44wuWTCG5Na8DLAE7ulhjVUDaqqqYrjB0uHb80tPGgV7H7QD1
n7cH2A6tH9ZAGja4yLaxQMsQtbJm/eZ9EPVTu3Le13MilZXkUWou36rns1OH4E1HVlhnQSDwRxVl
xdYzjDo9UhNFkUzWSiC9jLucCZn1qcK4FKOigZbp1qkQq7ak/nIHqNpGKV5dKAIK35Sd9k59J2EW
uJ8ygcT73e9KYQ+6q1j7vPbRmqAL0MkqMcgYNx3lpX2PZuty0oXSHAT68z9rnVsFSCN4/YyTfDH/
DKU2kQ3t651pACUhFQmoB1YuInmAMorbb+Ow7vjUJeRTGS/GmVrRorXvuV71Tfk+cikMiOKsYOHL
2UoyRbBrzYHrPIUA6tSL8S3B4Lph32F+k2y02vscQxBe0EmiJC2sVdGZUPpGZpHR9G0KK7ofsGDo
fA/xi3LqPFZo8GO9T8I+rgwCaVd+UxHe8zgrMnEDwitJbDAEOzh9HRoTUEbw5f+Z74wh4XFOiXro
Kxk9HR5iTa3Zh7fkqzGQUUB35Tr+R0Wned738Nzukb/DuksUm3j6H6rY2hzE7BMkzqP93o65AGES
mn7XBYf5GpBGuplOg0li9fjzyZsKN4pFhFalIKlXCiM5Y/zCEggK8iABsctl9V4L/CVW/fSnKG/I
zzfGutvfR/ZCYtZAIfIPbiraNtncccozzldA1MbbuwPcEmOXcaVh6jeHz0Hx5ll3tdsDJHoSaHdP
B7hMGqGTzgct7X23EMbmHrvWFLYMeca93xFnga/tFlr+SeL0AUUrf9Kl1xkYQjau9C2X0/bGiflf
4f4r1y+iJKq9CzAvzyQ1+qAyzsM/IcoDVHtkT/e0TP99zHaHRQe2au5bqlkEewarrLmAhGej0w1d
90La1qKG/l3elcy3dAJDwGP4oG9c3oHcoJPk5UkmqyCQKXYMJjuvU4/UBeiGnV0x5RDCASUxhvp8
lrxQ0cxDwN1G9Iv4Y6rNdZCsO2N33OHTjZKjDowWF7Q5trQoUDNI0A3pAlOI+t1hvQlwn7x6GUmm
VpPdHficBGMtot9Eu0lfPAr0kHLMzdU4BeuNXbGncrQNmTcARPBm2jV6DZ3XeZ8cMQL86Bg7fYwo
Q56+GVpRQey1UkY6E2+lEN1/fsb/3O8/7UwwmJmeMFaFL++wOLEhFWPzI5jPO95OGJtSSQYlprI9
KQ7GCpjzP9LoODqEDnO2LkARiszQcZe9LofdaN5/SpTS4tIt/5xXc9hS2cNo+KWrvsAtW+jOcD1Q
SnWJzKeulDWntBAzZF2xcnJcybmrNrPkG6asTXho1B42OTsEHgFqQFrbpMsfjV/Y4xvGnSUnyQNu
kVnU56XySJCkK96M3cSZWHR60tvmiTfWoN02ffKE1ODf2tVvCXxQGQQQIilFBCUUMsMwG1JZ6qOX
ssGsT6gUZ2FGLMJ9nJvBPENkLWfzVO9dALS1mm8UoiJgeiuNdhKVNUTzUqQTOKmutEBSKi7GaxLJ
MZvQ2KMp5zm5Jq4rzkYoEgj2citeCnR1qxzd4w/sVgYrvdnB7dqxcyqtCGxZYLIPz6H26gILkv0r
iYvR4FAn7u6B9+fc9ynjiFtzqxFcIc1hDC3m0KbKJXzx+2hqm9sEKrpusXsCFMR9onMiffT3cWgY
Cecc7jb2kIQuCvwEjGoXyBX9OqjYvAP33b15tHc1yjbelG0mJIMgbcEgd4LR7Sg6yWxrSmvRo7of
R0Yd5R8TW+0+HSi0CtWaicAMeNhpRVIEoBD0ooBlOu3Q2gDFQXy01bz37aj12twF/RVvRO5IJCQt
us8KGouL75Pu7iX6QJucLFLYxF8zVMkdAmi212DVFrDMLNxQ7HhlunS/4SRbSImXqfmzS7elVXKX
z9ESfy2ML85asWNp5KtJa35ruSaMoQqWmL6m5/zXwq0NxjcEytuzatHnX97QeqVXdQLwR3s+ElxT
edgJq15hmKIxD7g2ghuh1Be5r2r+CZ8ss1o6f8gHaLFjlODhADAdJnhwKId5nwkxRGQCArJohhY5
+8a9AlRJmghOI/2cbrLLxHRTxYd8NZLOtDBe9eFDu5vIVIYnX0jK81a7Xbz1HBhhaRNXTu/wLiDQ
M6s5sbLZkmHXOgnOgPiJx+CbQ9hDeCKtPibz7J0MJA29B1iNhuBLBWPyoxly0V2f9czJaegbhjGu
gKhjoM2Zjosafcb1x9PukO6M1OqbSseAoEKgwLDzFP2Abpcva8tYVo156ppLEL5c0s4GFTFZkSOl
Nmbj0VU2zj8BPUZxj1+XPLKaGUky5K6eVEkJiWY/B4zJ3sCiHm+G3rLlNXnESSUp0J+nmwm+KUqT
hBQtOU7d2xdQAClHrSfJvBbJ/mL49ti/F2Gp+LryFG7jhUaS6o/suttiVsoo6wYyoZQG/cPjae4K
0AHYlNro7qXxL173WMtGIIoYBz5cHFGoaHLndnlemgokv+tYkgttBa7Im22AoFH8/IUeMMJFZ/wG
NfkuprjtiNOUMMyuk/Hjn2kVRRxHAT2TCGI0byCdH4jkRNN23ihJ/wlziuyFcgXVTj5m0bA4Tqbh
b5XgnbNnQEIQT4nhd3ExAnBhZddf8b2V6UUX840TA/p56NymlKJdnQ8qW7HczdpI6Q4R7Uj4ZDtU
rwqjSZMrmdwkGRPOLfnkDOAAoxO1AX4cw6C4T6bZFcukOZ/T0p/V3l36ixx3tvKoRG06dSkMaSx3
S1N8+lCiTVfIjCxAf4eYhVmxA8ccQFwHH00tzjAO8beUuNDURIR9PCQZNUDlgyVlok9Dlh0yTnBQ
peN8xD71JBsXAHjnMvFcaS0VB77FyEhGLo+hdy9G7qoy7kZPl/ZUYuOOYReadbSzirQ8XNL0rkQf
1t9PGgRLCHTATiX3DkND+uvoF9c3mbbb2IF5KgpDtMzboVbST87lxs70usXRuOjdsu3gh20Fm26V
itww/wuBFIZhTxH3ksOm7xaiq9YNXQWZ1AuIQ4yYbdjSyP+Bf+79uaf+iz6+83S1rl1COF51uw5X
oUZKvIrR+SaxLMUpypAbqINhpSwW6UuEBT9qbKcPIJe+2pjhTSOeQkvGDLwossB8L03Pg9oYIH0W
Pm/79reY6aPcYtoJelgUdf3LnuY0G1FZUu6cTnH5KivrYZ2VrOGsqhMwjeUVljeE5vO3Ovbi8Xmt
5AA8r8z3p4uGz4ce0oDfAKgM8Z2FKZst1BnjaJYdBnTdQjXN06ARmJFBePPGnNJGOQPCSYhyxTcq
QgdG1hgK8f4Stf5ZO1mpq+UG5o5spPIJjh8ZjGOG1DCBM7lT+oObLcFUezV+bLmKkQ/iGcUHBRrx
cMUjbEY/66Y5rIVkc72ihJISw6Ec7hOKLn5ANcE2LaPTPMeyzui/LzGFqEHW8SNLxo2oBTc7iO6Y
TNtXFWDGmzw4UCrBlARTSlHd98F8Lig76py4b0Xp8iwJ+apMgS4glTRvztdySUdvL1FGU8WmgFyj
tG0lbmb1RjUl5hXMjNGOmtJDYhjfxcohpls4MKZbxukiTU4sJiuaFQKK9as2izJ233dW+dqvSYoP
FhnkC3i6xJjOArYIk4MyaQykKkmlIpJUYSoTcfRikDo/qZkEuF4LYDd4+5olv9q5xM7YKfJ+regk
Oy+BV4CRsYyhJapCDlDRdEscp4O9LiN7Uqf3g+J2YaQFzuNaMsZVA7LNcW2QJoarbjiIYgcimV5q
C08D04OSH0PdSx7vFsZ6WTHLl7s4cFQa090OoVgiAkLBwMJaYPC6HaOT9mBmXHsHZL1ofI9fmM8g
QuXUtlfQqQgtNi5s/ZVuNCtFupao5kxKwMJKaH9n0SeTBVRW10lPd/DrB+h6m4dg1W7yWTNCo6FU
4Ln6RDH8qpIiEiy1UoIBYlXE06rYhxzk2H0CQlYjGwPJl22mvmCQsHloAM7WDgFzhgmbiFZre3HX
oqnF3vbP+3ZD1MRt32FEjauDeSY6J8PgBIU9GhY11+WTIyDdJ9LFbB2v+otRnrmVSu5ow2mTp1gG
4yt9yt7a0k0IselbyM28MngR9k/PyB+iHn2NRPhXiTawIT5ss4CuoMmCHKyThQvIbL78VdpIBQ0i
BXPd+JnvZji1uG1K+AUngG/+WGJoQfm6rMBC846CWyjwkf26BCXv8HLWiw9ucq9VwUFH0ObZLqKE
vVvvOuBdweoYMyUbbDIfX1lcZwKK6WYEoJ1AAybWP08HJXV21orP/NGmiTVceFTfUCtt1IkIeWuh
afwejAhhFN1zIG89vy77SUDXpiV0CGLPcSvHPefhlmtdWXXQHGlY+dsEVDKcrYn28oTbwFwWxham
fzoJ+HfQJVoS/chZHCYfVdaG6ClCB/0JM1fQFbX5KEdtrnU5aVsb5bQkvApBnlzKwcWDZPacWk8f
huA6LRQ4fyhtDKL/e44xzzdEQNG7S+mEWHfcM0Tk+w8uYsXb6uhoXXBIKGqhA5tiXpVOmSXqAA2P
Y2q5O0jWAMnit+Bj0w+ZMtX7b8sQXo71+cjruNs1ml1F+JEXh5uObE0/gJqPbG0p0FLRhGi47jVZ
ss4XYIrHvkA/z1CUmAEB9tzaKsdlT90nJ7/F16jLET7zV0GOOVQ1FXZ+sOr5YAGkztbs4FcfFmh1
XU4iosEgrBKKi/cG9oXfiWaSxJVGOF40rDSDQhNY3QbjED5APX4+15NeP6QTI0/b204F//n5uIdk
TqEuRPY+DhxsnDaMfAARqBnYByr2YKTXW7dg8s9mVeA4bKWetWu4e0JAu63lwZ5EIOlIdBvYfXCA
EGqTD1xdrFWDfJGClnj2iCzNnTJs2XW8GaSHA8oiXkD0BqV9OQGLAGHM8KRp6SbovE8e7bhOoVHs
z40F3eg3EUE7MEeuXSSuxoLEfSh+rmfxNRVgp408bzPr1F3+uM6okXoT9BWnvIY62i2TaA1RaK7+
h3jLWcpEimQAhy2ym+zjsDZ89aUxY+BN3PvXaMh5Zy5FTH8R2e0m5YMf/ahZDIh35FzIQ0FM+l4n
PLEFz+Fr3wTZUpx+VbYHnV+MTCwWZBaiFeZoyF4I295eFF3JayJHnDao1mh5sGuBJC8zdJMTAleo
RxGo5nWzzzoxWSVAX3cO5hkgfQ4DjLSlDniBEJUoiak2RCSaajDJdeIQ+ZMZd57MlBslCuH2GMDl
7cWOX3MtWzV7BJCrHKL5mf4IMurSWGxyc02LlRJ1mwLsTtNREAI+2yvWLmMqMGEwH9orXHLlulcl
cqm1H0NDYURCxu/n5QrmzE3WNT/UVD9kjWnA7nHGr6TpCByi/pgc28llLgXSD2X+4kJMiGFhfwa9
I9HQjltIM6TqijfW7lxx8xgkJpgbiNihxcPeNFXFxe1BuzF6H/E9RmTGSRgfvkUXkK7Cvp4T6soI
eXk/5+UDkW3AkVZdZ4JnHesPnlQ6/v+q8hDkW9rAHTWnNvLbMk1S9wsPsVI8MrAKaT6oQaUNEaic
WQ287H8Md4cbxlrsLGl77OkH0u4fenz1c9v4OJkUl9Q2NYGdDKFdWHmKcffop2JpFUKwR1C/pZTY
n6e6cFTcDrpqQ9vjRpdOlgN1Ud2aBohQXKXQIXARTZnKVOHUs+WwK+IbhVq2ooGmIxaWvyofnrTH
1aBnheT0IQCpNUyOmn2Vv/QGsbDVjlfQ2Srkz97tviJQsmF59mIDB0qFk98+ts/7+PfMiFfN7C/r
zOYMSohda9l6ST4fjkKxok7G4fclhtOHaA3brtKoTLTPIqQDOcte900AWmxXNmOa94ySM/SxxmoQ
YonPcT9mjD++pNAIoTcjKDOstRDrK5Nk2hpRi9XS08ansVHQLJ4YfDjvrW1ZPKVuW4+0K3yHRG7M
6cCOOqcbqNKYGpkqhUBTnBLflSUpGn9UJCGbMA486cRtlGd2Ir47z7yFl53VrWaFzVrr7a1pFW3O
Pbta6Mq6Bx3ytc4FyR+/Zr+is7FO5C2S/UMGSeTTxeOZkazIntaxkA35eQRjEPUWk/qv3G0y0BRj
wUKzxnspyuFV2IPFhC0gi5eSpJRK5mySR82Fkc1aqwYpHExebmuxwjZC1+Q7BrEfihtT8Ur9fYph
M1kGWta4diT+Z6oSkcmKHPwGeZFDdp6KG70NQ1htPT3nTBzcKjqmsAloAmWJd0PlmzzT8f2fYWEs
oiiw19mFQrTNfkEOxuJnmUjJzIkGgUVi4cZba73Ql8aT/x9B0b8dVel3eTcAMrhy4mX4jQQpS0Me
4sut75LJjVh37POaPJJsNrn4y+GSBpQSocEZMFTa2E0r40h75guhKR8iMMwZSAQvIxLiaquNL8Kx
W74Ho7fIp5mh7DZoPJfx9mNE+9tXSRnbvnpC4S2pDQMJnG0sKCvED0l+okA9WQKCe1SbEbrkLmpy
Cg+iBbBN5XHlokQbYcSa+Kl1LN4CPkHC5WW9QUDrA/ULf3tnWFVz3G1HQwwbKzwu8nGIOhALmePN
6yL8OUtnJqN2Q19g5I14nXGPir8bnOlsMcK+b6d65Ois10URtq5KsUqnuZS6jMGjspQ4sp2+zdd8
UGISlbtQvQfapCN97E9i06jbQgDXNrURxzTw/XQbBrmlUkNsyWkmU0yFh2sFJObhh7Jhjjwq3s50
RLYUFOQXR7CFzfeIWprN8buuBwKcM1+QjE7sr7SEkpa0FFH/1U0wLNZRor9WI6l2PJs2uA7H5nhU
hnD6ZApbYk3f4hYzlZfJNmSiGQzdn6Y+L6zTLTycjXRwiToUKp1azKxNqTKsfPYjCjKAIA/LA1h/
hi/pRVnFfoy2xxh5rT678derW9d+DYN9SUJFBjTk7Tv3oYxvnb1R1sonIKzL5u/bXMjgaoPp1c7j
hT4LHDJ+XiFiYRXiS3SgZopnulyFX6IwbYhO2mZ0cy8g7Q0+cQ+mG+1DkoijMuRJsC3BqENH1508
8fzCMiF7Jw2ktH9Yhobh/leq9eJ4znsOnEcHBJfFEP+m54gzgyaRjdIzUktnxx63dEluL19IzKAc
/d++vUquq18hFV1XdvGptu1akupQH7G7xS5YB7WNlZqgJhgiOe2yuuq0sIuoLOZBikX+7iV8LhOB
9btM88ONJn0XOSb0E6liCFsnVjYvhFUW1R1ABD+xDdmazophR0UttbkiZx/OsUG8vTe9zl4c6dcz
OVIFTG4ClPlyEOXLDAUYY8HB7yDiu0QbSsPezQEFzkxZClSCseSqgeV0rnXp8emEE2xTiE2WQsZU
e6Fza2NqIOS/F9VvP6RkQQEjfbOouMvWx5t3WA5AeVXYM9BWo0CK6/W8Nv2hJAf6wn50AXeiBBwB
LY4ERntWoupRaNH/hH410VZexh7O3f7jlYy0kDIOdjP4GfqnGe265t0fwBfJX+WQHPGHgU+InYUn
D3N27KlVvTl+WLUEmpR2DvneZJfzSrKzTYS8VZFkJNMLx1E7ZRlB5T/fsOvUszr3d82P0UrAE379
Tx0Sy+ZEupnUP3C9AMDvQCz20VYPBKDi6SbbM7f/2V3dqgT+0xI5fltWkuf5HTdRbdcYTNVFUAEu
4HbxFQVkB5qvCLWedrViMqzYFnFxd+6t2CwYxW7T50+MONtJmmOr863nrXmozafrNeLj+ym/PbSe
uXASZ0zB8NEjsCFp86CS7PLImtTLlw0qD1AfZCORnmUWdJfVVrQMPPdOKgQHyeZMIkPr80+vcdEv
EkGuGQXuR1jJO+XSSj33AFYQS7lSOlqxey/KeArrwzgvtkF5aLIc2RR2Hy35MU2R2bUJRrE76gl6
OtCvhLpj5zmVvJctMLbgDYKfT+MU3egDY6j0J+ILMn8+jgAmqsA3R4YiIQpXB50jBBQrxsYwGxNo
4fa6KT42Ci/ds/y+XA53Z+5rJtoEWJWZiQ1SBetC8liTsEnILK5GaHsM2dFWsTJZNbJjd8NU0aOg
kcIXVSb5OnQYXgJytiMCK5lntWkaGbCnFnbyM4/3KEZYbY1fsbYvcQ/RwHcx14PbLbjxn5O096Qu
NM/LSoCVigc5cG9Oh2Ub77VVicwEzh2r16V+3H2fOWQj/wZeMuWzGSxUwBJWAgA21shH86fn2p5w
qrLO2MrYrhAUrRKIsGnve3eOR7n+NN5Wuk/a/GkcwgaQxwawhYbfHlCNeJKe2Crmj/dVOXYWQcI/
4k2h7d6gZsCk313u2uRQJ0eJvo4boMHxIBA+5cMcUKyttHlEbc2iiZzQ4PnT5UlH8Fs8fnsh6OP2
gO5ibRmiwPk27IuynJfQNhkCrw8PBCnepGF1nn+X7WGswYstqqETCcL6UtaqCDPswbFaNnGUFy/W
9slRS6gT5bPjhoEtxRGrlkm+vTaKbXUeBhxLalHklUa1DPm/JqdoafWFUGPzN9kouFZe9+tDS0Qb
tfEIuuFk5zAMUJuotHBQDKSrv00nvjbeFQxoZDU3h36EpcfziDyyNvdW8OznDrCsYOLp6VCA1trn
Yw4wAkVI6Pb9CjqB10+AyJOSpSN9oxy1rodBIXzoNlchHvMiRBUUx5RZ5ymISXJheztqtWFoV2OQ
LRqlyjgwotb+nYDGpvwXGzghUPIjkdE6TdFbiRDyNh+6ikqMSUeqwiEiJ3bYonxVrZmcEXXUn0A7
1d3zvgeidv2CxjZpmCCGnccAMkh4Hn2RD5Ay9bS+Hle9Qpe3qHQl5CM36tf7YOJ2fyUaWslnQX2B
8YiAsvxgPnWErLQyoB2l9sX6FgF+/hQCgjA95otK6tF0AiMv8LLRyfKqo85M4atfHgd8E9+7+Q+T
NPbm8mDS02pjOH2Z5HemaO0DdG22YCnjv3GdJGUbBT86U9jH+lAHHeIMmOQeYh8x9l55GWWrrn75
GUxsI3XEtRRJadwByWgn5ZGS6sCiNW5E+LAjIWFPMdoEJ9CFG+G2LS79f8M7ACN7WCDHDLBrsGwA
De9PWB9cje4SNTCkiKpQ3ZziETzQVppt40XV6aQ8Y3mTELf/WfCD6sTBTHdvAiVrcPkHfbKHNtvK
jheZDTaGccAJYUAIQFDvUZ7rCmrF51iMCovqSCaa79j13UB5UPkC37np9VrdKp4mNQpiZy742Fgc
nYrob43Gkh1OnSOg7NCYRZPW6gs+N14XQwu3n3UDG7q5KFWGr0qLCFUSP7BDWJSEX+CjSfJPKqgA
4flMiBD2qJeC+GqdZTCbnvStqCUnsUpyWqxojh+IEW0vygEvW7oIV7CNlNmS9IaLizQsZvmlz2KE
QGRxHf3mp/ugqQRTSgzZDma3I9XsFZ6jRwyPSQp96TZ3cs7II4yiS54utWE3JEiH+qo3YCQ27CNi
pimE5eNcqXVS/nogoMA+GVbcK+ex/9Zwt1ME+5tVE2tOhimHVLOywFfL5A4db4sCxWCtAffADc+8
eoBtXAcs6jxyVf4sC0aBzzjF5FB7uLXRatTUrI/eH/JJ4Z0ddB2S31FRXEBn0fdx2CSBo3hicAEb
SLH+xLmTUXXfJnZR0J8itDX8di/gb1AeJ7bwQ8qQ5srwrXXtSkRABjQeNT9Mmb2E5/AlO2Wj0URB
TSiKqXfWZl6/CkiFw2H9Jv6hkXZdlrOJHOX76dYnuWljLbQVVTtePmCrhu08V1beKpbzTx34fMxp
/xGGHbGxQC21rrSY31ijd9sS5h/qA4E5kIAn2BcjxdOtHexwckgp5N/X5w4IJUO6x2ZvMnO/oa3D
aaeoJqu8mzZskjgEWR/AZfWMtq+49PDyu8csdE6jSKW+aKTC0Mi11BuFBqZbIljzUeJNcqjH8Unh
8LKmg0lbnM7e233XPhQZs5WH4EV+dn90RUkE2xaTsCLiqbSZ0hbGw4QkgeZZF+Tg6oZD3css6LjL
qSz4XNCGQqaqgBGm200p/6e39Cq7Y+A9vSksb6chlq2W7Vsl+JurfQF0fratpQNnraKVN7MXkPKD
F2fJqCQET2i637tldeCN1Nm+SwJTK4/Ffs0wERcGNcg+yFR27KiuojnP4Y9S2PXCA+GX4dP6GRip
4W/d+LnZ0OApCezQWC+U1xeVYolR7+8MKHX06QwCYe/xVJT6rw/54rNQLkgFavQKzXjpM/MagMhr
8hTIiuXuM8BmQTJhFvVmliHO6xOR6VavDpVW/OfhtAyIu9axgRCOImYBcO896/lTIRaH8yqnAy6u
+HS9OmTGvHqE5r7Xl8GFcWt4AWR/BYRzN6seVImWNvT4KUbzqaVd4TSMFfXml+VUI3EasEITnHE0
mfSY1poQRyGnLB+ggfFfTqCHjB1T1WzHKDURMN0AehPPizvrATlF9yz+/PH74+szYJck/MIZ64EK
3HEFfmRgt7gNi8n/8Ji5f1GU8OZ1rKuxuJDNjnj/Qk5Xd3/RlxZAH2p4ExM3mKA4Xp5cqw6cB+n0
tC5LcE+K8RHBRdtQ4WvbuUu2urOzLe7KAZgYHc564KByUmDZCqo1b9U/e880QFtHd/xj9fYfEw3y
iFo8xa8FzwBrF7QRv2hlkK6x7GmRJlhbIMoorV5XWg7BE0d33AmGwBIW9bV7olrrpxs8FwV8cIRg
IIXmGGXuJyxx/MbfO8y0uUTZOIf4uz+MBGW1233J7y34ydFnidJPyQ4IMJCdKW9M8o1mlxpy7Efh
YYTy7KM7rPl+AaHfroDpi0j6DZk5zsPOYY7c/AZlYDxUQ3fSvKs1LkX/Ee4p/+j/ALVeWzd4ql5C
8wI5DfpPC3DYyqiVP3eVYzxkESuzcgd+q3+9gEU16o6Gw0Emd9DK0iIf6lFFTbZ76MDfE5wCFZE1
gYB3LoDgakZ7Xp1mrVVMq6etB7EceqMFjsQ44/sdIGCoPaQtVClA+XCi5zCchzeGbaWZltiQ/b7l
MDvQEtdS3cdnkjMg3LxRYB9NQT4DWQ+NHRhwi9M8P4PKFEgslMZH3PheQd82UhPbKWUOquZ306C7
lRLVJiTe7udA4lh7Ie9e8AQBMJPrMOJU9wHR0+aalqfi+XFHffr7zdEWWzrycrkavpkYGaG7/znQ
0wlv3z/cZWYF4Oq4b6oEkCwCfR0BvfymOrlkxV86Fvl7oKlJ1Z/0//L7QBpDwAHZXkbfHh6LaqQQ
hXzm6HAXPZOTfnnIaB3c+TpnOsY12uEpjV95D6HmAnqf1+8OqkmP7PrrzIFMLHyjrDhPcyQKZgOH
WW5pUtsC8QRBU5zX0x29o15JEDFiD596kT+jhRpDcPBuF3Pbw9wE2kkeOOl4NWhI8fS4UPmgtMI6
C6ff/zk6Mw4EwMkOsSgtOEWWnwqajpggONyfzyZXgdr/xju+HlDhLWOSL5ZqHZoiY8mg8hpasTDi
Wu0sYSivxfcaqNeOCEonLv1/2hW1e9UsHATBfSqRnu4Ng603AUCk0M9wEsKDxZRov2b08nz6fvbH
MK27YGicHXl+IcfsDW2de0OfX9DtM4s3tZfBf6cIEazgaLrlmozJPcArsNrs5q6ZzgH5z1SN1F9H
91zgPWyj6Ke0eC0T8EB56UGpvwaVX3HWal/oAeaakUu6d5YI9LXXzDnpfLKmzXeuPdsciug4DsxS
fXbalXPXu8UnsykgCND6/g+mvL5AzbzMNsCmxeIOsCU+qImylCzpIxi8aLofSgIHwcohij8xv5Xd
pQLvxYSkb13cJzvtLrxFTxNkNj84FLjUvJZDJaKJZZzawQmeveFklpNyJsUeaAy+rm0XJuih46Sg
1Rd6zQp4WbCwQWZtkTtEm50+BWeSv8wpzDlA7dH/riH+7BbSVjrewLer5Xg97djhjfUhhoV8LTY/
fnsTXJ6bF+jy3nCsZILqm8Y7y0Qu4OVeotn9nrABOfcOLlmU4iIAAPxb8TLxBaVTev1ZHUk3X26k
FBkD6e/nr5G2cKbzN73HFuvqiIrwuRYqX0MUwvOtKRn6sypKct4enmtf8BbaV4LBfqfPJcG2NUev
GnfBfR+UbXAxcluQ+qWSD8Jr5Ss80SSefHLcTkJwO+GrkT2OwzSFin6z4WWO1ZtjkRKSuNp36PDw
1NSwYgumg//z4Wz7CJJLYHm5yt5n5zUFJz1uXw7qyEyz+zo3jDn3Ozb1ykLMU97vCaYExths+vkG
J3h7a5D9oNVlQeGKF8Yz+gUWyUmtDwMSbrYN6kuhNhhsqFZG6WsVrPilpRrfl77Pq1j69joT9owi
YFlqeZPLnrC5Gakl6BWfIoOK30ZhVXcgNN1+UVi7zoE3OPvbNqupyrOgLDaSpgp5h9Cf/RSHrK7x
EM5c9i8ROOcziEMlflXp8S1p8T2KwngZL2smd0GHGslP3qFnHMlYV+wBl/zy9nbmMYZP+6R1IrdX
OSVvOpIeKZBYp/CNrEfLTy/wnX1773WOp4XsHqPoB4Iy1B1YW2L8aPzc3V/9l3AnezjBq+usG9rR
GYLBj6uTV0J2ICC8h5NL4YBdCctkzgrgvNklOdfNUqocmmnATdT1ktYNLR5mhzz9J8aDMhH18FYR
3jYb4G+RebZwXgfoE5k7SlVSu7Lwgk4ZZh3pwzp8i3dOk2gX+mNpOXSdUup85O2pbHqZxnelyUMu
rg7XNhY6CQWQrbb+d5B2o2H6Vz2rQ+q8EIe+/LWWZ4yvvYJgHO4y8Vy4b1KOOce4PQAEEnQ6gikH
W1gnmLMLi914xJtVJsAMYCNaJ+GVk7bAuDrQ/MnNTqt48FLwNK/YiB4TYjVlsd140B3yFzhggNwJ
hyQ+ZgjO1mLxtjJk+xxUQeMHMlWdqtYY6zzM4AjvTB9Rf8+a1r6AAhdc2+/+5oLBrG2a8L7QCvch
kwChpYTyJvdtY+PdAtPm64P35NzzCv7TOeP0wl0BurtjAIEFUTz4qr10aTSWkCeV1uCXENyNdPcd
NmOilnJprLyaBnXlH0FhbrerjXDdNsLYawduOEtgPD8Qb9K4SOpd3ElvHHyA4GgxRFXoDilbLXJS
VGOaxUqMjT5lTBOHtpWGHyr0VK+UuONgAoHaRFnxd10nxOaBb0cVX2LRAMBblfPc6hGbpLVNK7wP
qIj327YZ2ZXF8Zd4+l0fO1zhIr0GIC5T8qu6j0ERz7D5i6ZQBqJyaojlpV2yg9PYTQDIS4b85JF3
3n5MvcxIgwvewVoLDh4SUM2EqZmLQOmfzlfYt+sKInXl58g/Sq9pBJTOqqQso6FBqjDLLoUGXWvo
yXZYseHGFWSCq0X3DAetreP8TOKq+dMhSPRpKOlJWBJWprlg4lvd+skmlUYU3n3QyRn8Y4fI+x0s
ECD5KQPd7nZhREZcuaplqL3/urhfzNBE4I8NWIb4mtwxtjK7Hwbgeduqk+s0GeV9Gv29jD2fxBaC
7Y2BUehzG8fxNYLFNsb/oMSkuB41btavkLueLzqttcHqQc/TG2Ypm1yJ5S+oj0GGBjJ0i4Bdopxd
PC07LQPS4FMxIVfYy9qGWrTTTeNM971Zad9McLOiocsihl334kV6HImcLkowVHD22zvMiDwaAFE4
sUaV8h3S/NCR68HPjQX1YNRQrLDeVUfriPkMev7FPUmtpT/0Z2YQIxx3/7mSKNWABI8Cttg9veSZ
3y5BwXhvpg3l05YqiZz1kiAKP4s4frqP6EWGT4cGftfYC8uLUWmw+XA/JgukyO+YDQ0Mcd34JLg3
fH9Z6Ghe/TOvUrg7MoDyUG+5XehVk9ubpVAaM+DnSlprlgHZzlGvpmL3whzf+6oVIKgGSsz2lq8a
srM/M7xa0H21TUDH0NZ5fURLoNQN8s9xPBFUeF+YG5Z2KoNHjCb71qfdb2yD/EpsxIKvd+lETtfT
89N43zCIKrMOWwokv/6qRa5SBOhh3M53ezmAx7/CHgNvbaFnRs8dw9cmi1bQW/0ZmWHeXyeRXu3E
ysWG9NOo6xtPprtmId0O66BJ0mfn4SmtRgn3hfdgoR9/HnxrIpJxWxbjDmJco8m/SRHAoen58lbS
FuFrxnC26lKLmmxSOI3NsxTLqCbgKn4z7qLyPpTlrsvlltAQjJ/kuEJW+YQFJhZMUxXFpZzJIuXn
ke10HbQ+VGBtRNoYq0dTUiyObBnUrmS2zVfpuz450Ycjy1ZaI2SCOR60bFN7rQ4Y7RIDWL/RBjvI
WbxMGq/TsYoz7cqbe2Hlz2C+1uvIba+44mN+Slob6W3DQhsu5n5WSNnjn8OHfc0vJpYlfU+XJ6A4
H4fhxLbSxDNmleOudjfGabEQL1FvECx+H/EWf4tRCOGi1aQj3CO2hDrI0f7RQkOduG2WNZ5HtDY5
mjsY+QPICdHKDj/Q4IRWurjmKS5R+q27n3w+zYra5AdTS3SUSszd5ySqHBJ2W8UMF+DeYJsa5zHZ
bwHzIn5Dql6b3bvi6SM1cSQzHCRH3s3xMiWXP7ugysucoeKyt2Uy3BTTYNGFgVZ2bpqNQi2dvkKf
pFY7frGzVi0U8eaxAc8rwoQAd9mK8n6Qpu7cfTgwOgWJXsdDyruko+ul3AxtsOBvq2Q5BPOzvzrO
ew9TM+X4bpbzKgsR+eq/GIg/yOtPMZvDTjezjxh8VRU2ouzIXjh6gvAKJQCi83IWHg1o/nY9+8gO
uX+Knr7lNPj+5Paf94U9FN6oiMCd3vHi8QJmNMA+jg8rOKD02WFpxvJ7ZwHBSDRwFhU5HHxt2JLM
sKT29X7xfFwlbybxlVQxA69FUuUUeCp2flFlEhwRZmgZWyFhjsmf3DawbVyn9CZBkUx0fm8+Io3d
vsU/9iLBrg8L3sxEKwdf/bn4d59gqDRG/oplXB0/OCge4oJaSKpIUmKCQ7c+Cs8q6c8qbjXCznIw
8ydJYPNp0Cj8KaR08V91JOYI19oJe7/aLt/sFq1RVWH5OpEDWbzzDhfMtDgmX2sQWgcN4UbKtifC
fFpOdjUh0g2RMcI5pajE9aSD4fmw77Udsgzf6RBttUJm/D7c/vVaudyVUSvLIVF0gMJvv0/1WFRi
O8oLcIaDHrXsff2IXItvDT189PebGSj2a1tR2qQ93t4x7ub4IyRK8y3IXVqzFoc6in5va48K4ilb
cjca0fPqASpqdd3fJJ3aQb+/lljQeQQU7P0ZnGlk9Mq60W8x0PMRN25U+QZ3Jqqw15b58J6m+V+r
tHR2ahoobSoW8gCyKpphnDX1CaOCGTqkpP1FjLOHDjF2qzPGeWrk+npCZxwXI9mr2gXq/Q/KiPmg
4+cHF2buFSymTclQ1T7ESUJmHXBK+PGqE8fjsNSg09ApSAEtvi1dLZleNhoourej9XSxnRHseE27
hEsbG8AeRL7YlPl+Sg/KMdBn0e+4ckjcax4Y94eT5Dm8bTie/YuHcKRq2Jq2qf063ZfNpJBU0JPL
VvCI6HuyGhbCB7EShTt1HFLb0F8GGg78Fi1PXHDQ4CusdSK5Rfp/7oEE1X3CyDoUrtG2llUbkrBg
2iqwe+AE2Cvrg0akfKeVabe5aQxaD4wFK1V9g7f9mdU0jltQl//Voofam2RMYIaWMxSbpBuAlGE/
K2HOvBdUfvykOqirhYuhLwwSpZNNvgoAD+XElNMqpqRG+Gw/bdpjxX3+0a6M2r9ifUWROaPEQV2L
ezVOuBpwgwcnya8kfLowXidFCcboQUnXUvn7ya/joIJf1FRd6xnU+pXE3bhM6TRsOfpNMxn8ef0G
sO2uZxaIkp+VkAB6Iadqc0m49HA4p6nSZnt4aG7BR28ukh3eDU7vJgR/79H/+wWRIalmrz2L3xLg
MOt5ASQpnTzVRFe5hZ9mEIwf/+hfzb7L/4ag0Raz0JjqcM7RlBcAZPur6AXF1ezq06T/+Y6eX1mL
VP9QuORL+x22JDg/O6eb+cYP/809G1th5P8MnNCtoco1k4SzkDV0sS6VDYJAtF7stmRepSNzuERk
Pl9ZSGAK3kHStHFmw0rR3T4iTQCdjTVmQuQIpv/AzKoc/9n+zekFULq7sPq0xQV0fbMvfIYU5HKm
HjSTN7xE14T+Wawm4xxcgnqFjeQpT8g9+0oE7UaAVngrhEW6zlPOdcPwASd4n/MM4A+Dtoa4tKzM
ZHCSUBuTHswaN4jtLO7nG5wBiILhrMpVYHO0q5+5rSGkKygkSow0eWMyt61KHHRaYOlsawnIYjb2
Gx1OGs8xIppEn8ZuhtuJoOHWUSb1l0OdzXzgVXJbNP9Qi2sCwxouY3WfFRys6Yf0LPNwuqs35roc
AfOfOZhVcoHeXBQ8T2XwK5iLJWXX4mmeJ6pkOZpdp6B4Kbo8p59+cGxzVP7METAfhF8Shn4fqlk7
yk9Uo2OCpm/nKBldHiRMgcZ9VF5ne5F6DabqtgjggWaOgAFeBviYWqXOc56Akm5aEvTOcB1fE6Ap
blSLAIfjXGog47AOGQ4xxlXTO+9k63qH6NnrS5PkodW6JEMjixIK6arX2jn1xUuTvdcY/pjWDOos
EOwAaSQwFB+UExful9Zf85W93wXD7kg+ZpgfGJI2ltN1TQQBoWfcCwlmdAnvUkasoC1gMhqo+/g9
IciFD9FFg765Mxt3Mb9Z3cLll4gELe6/X5oBIuvv56DnI00XPYFeivgT1IAcG/z1LHS8DLE0G3hz
hJdfCYDm1/r3YGCkz4gQX/FXikBq1fp66feHx49q9W60z+7pkG5snXR052XU7L5g5raXCN+tFFty
aBg4S7WSg/ymu46suNbgrPcyDBOH5O4+ucQZuLHtMUogb51t9a1ztoMiAQV0EhXTGGrAYFeUIqFI
6E0z/U+ZDZ1XyjkASlfIufWL78I7TtMi7ULx/pDoZL4L1h/an6Akw8xiVc+VApuj3dmiqbDhC92R
kg5yHqWC/hhRP3TmqRNJN7RY/Eb2Ms694c3MG16NN9x+KMlxrhZSemNHornMyYh0ybSpiAF45f1Q
THyGCyibhjLZiKGZ9Ffz4w/6Fa1l9Oy9LKweSgMZXFCP7VQsAhfUbuleKRZBDPSHQmsk3qQGv3Op
oc57Bx7gGweAAM1l9szkDaQpHmOAVo/R7kZLa+eZ5HJ/LXsekO3u4UJdX76xpQO7MyBOihZZkXq0
lUgghCspXn77IlHXM1YCUZ50CAzlmLG7puJ6tS4Boo70LqiPgLEVMeGr+q3QOBykhTH2rFoLyQeT
1PaolPwHSM45mVitm1zPmp00M7LJIeqtZ1TP1j6dAae3VytxaKW3P/Kpg00r+W4/dOEtSVpnAU18
6q0UMQrHG6ft0r2HH3HJXylHlpqLWftFZNt9zJiaA3gC1TUdfdk7TZ+DG7YZ9OO6QClU54xBkV7o
GMEPQ5EHlBEqTIlrDWWaPCwnIzMtCq+E+LQxuhzbBf9ZHNKVOWVfYNVrMjsFrhnmsNaMXXMpBDlm
+muYB/RvVY60Zy24IwnNMdoutqZ3l+5QN29BTi8PgpViJXiYBRYFgzki4n3QmKlW8trm+JB8qLeS
iYBzBYuzeKCTSHGsYED7wgfES8ZyV8CFj12hw7hC0fNJUmoG6v/GgrSRVFuhVR5M83oxvaM21Meq
N3qAig3tk8LGK038Yo6BDxyaPLAzwfMCASS7U6k3dDs2Dc+98IbRnN5OixbTmPSN5eFZ2gmkslOM
94cjrqGEjamBW3M5jdR1dHz+tIBjs9IUCm7y6KoEfPsq4mofnQpPIlYI2VY00hg0qRMutwMweX3M
7DXf2RwfzaE9I3bRahw1XuqnuhVxv9Uu5sEsV8zRPjet9XVI18ajbrV/zvFXXHwhoShMkPv9xK/G
UpU9mGN+yBsi/8HjgfVxA1anT0sN6dex64qgVuCRHFpE+6PLXc3J+Foo78Uf7gT7etxTUgH8s7Le
lpi4G63lKKFoDxw7qxqh7LQ//JqfNZLTRP26VX39nzdIoWM99efctCIN2ZZmripofaKKZli1sjw+
DahRRermTSiYNn6cG6E43tJlsNPlTOg/yNfvu2KRDc1lAA1JRPIIlBD67Aqvuonva3QhineAPM0j
US4wqkWQYHuzkB3VvRe8hPL+FdXcz4SJVUN8vn9MurhlCQFv8q+l0C1IhUeeUgsrwx9hKjb5nY4J
8mvjhvTtJcFnbUI62mEjARbvlkb2LaJrqBjehoDylu2NnU/JAparxyJ+gNTzvthu4yBSe0nUkD2u
DFTAnIAFj1HyO9TUZ17Oq9z8sZERTuyz5YeC0VH4a9eRfy0tjJCOXfYI0THnRbPY6AxyTZV1Atgz
xK6WbwpNM+s3GnP/DPP6wcNDfqYi/imm6BIsQUG1wA3G87eQYmM7Yol10A59w4BK03TQ7GLvKAcr
woPwggp0bRFL8bWoPCTKIsLu8VOjkIrq7eerwlD4rxVTxc9tdayOXyXdvkBlCAFlYKrCqZckyh87
SIhq6LQvckjJN3oatnFIIDyT5hAj8QpZTw+cdwuZoIRPNNJCrVkqUcm9yKaiZrkv1c5AoE7rTHiI
jEjrSfV/aMYq/tAtW0VJftim2lHYu5Y2txNof9k2vadWp0sz2QTqFPsBZDExMqUKdHElSiA3ec1h
uD533j2VdtuGOOGIRs98Wp9EE0lV1qvb0dVHjygUrjwlgxnaO3BVAZ4948VX4z+TejO9uhRcydH3
ZweoOGwzFnovPNk6GBtEvI88Txsj1b2ZIVV9JUWECq8G5WnlNLt9v1IJfmc1O5urwCQWfmEQjl8z
vchXJdUWtcG2JC0d7bdNSn3hpqCLiceUVHN9LsSOU0wTF1WVYH2mkXIx1MvOOmjtmGMz9dnW9pdY
tZ/KtfFxMjjtMZT6CutYZ6o/GIwSLzeFqlGihqDuZjlYUaNMUFKI4m5Ah8mrY5uNTgsK5AQD1ZXc
h6GeIE/exP26niN+6/R2LMREA0vkwdOZlxNYlQx7cKgIMYTmWozfeUQQQLKIID3QN9YXll8SOOpC
BxL4k7ukCS3BSLkSApCL9rU8eGHxn0UDGZYTvB4wSD83pF5rhp1mlRQ7qrbXk0r6ifXje8/9VO8U
O9uqy/MxF/juq6L0loDiy1715qQR0WcA+rjOBTDYqLNFKuu4vdpFXOVK7gjDH5VHZWyYBrkIs+O2
cUNuVCsHXd9wiSxbvxxjaqrMKukvhQxpBkDlgFQQ1v4+vExj/OTw4baAWxhvWJy3de5BzD14dJga
0PN5bvagTNm8iaiQdIxf4M+ml7v/MKhZfYR4NLqCAmjKVW8hTW2jiA6aplnh0V2LXautN5/yuITC
k9JhQiKPgfmGcYvN8/bGyZvEWFY2aGmCr/6ieYYqzHXEhBzU/8MjFZACgqVZpr+HZcD2S3eqsd4T
df7CFfC+pNMYf6ipn0nGvAsidiZE/gSjMAkRgsinqeeJvR5x6V9pqD8mk2EYfNCXGvdG+Hqksuki
xG/meygL1KEv34tqD43sL2dVFj6gZ/9pzTGdI5p0IDPuhvYx5XlxNciqu0C+MjKhkUzNSsJRckof
txfeTAFBlhJrR+n01kOL6ebVQySLrK5dCUSAsQ5K5jKzMZ0FsHOrYBtzMRrzqPGl9f0quhidVKsv
V+3DSFbG/wPLMbvfbd4c+HAe6JNUTIy3U7TCGKptu9xRq4CZf+kON7kEgsjH0FJSNK344XPevAlk
1jlBaTA/DEmqGV9opf9Z0/Jo5mQIBj33x/FQdP6E5WzDO/VBKLVVvSjbXvQez92bFJKgXwfxlqf0
AWTo5SQQNtbFne0OA/c+P8zfR+DmNkxxheDrWDDMwYUqzPGYFOIybwa/FEjgt4P09luGofnkrzNF
tgh5KdYS1cfoiTasrEyxWn6a42absAlIYnR9RzgxMBl1Zbtha213vh2vg7xrZzkFXxkHjpgI8kTz
itFeK6CcwABTiN54IyijwOP8VcWzBRK3/kAuqkl4WlCgXKmSqbCUVUPZdeAxWX/I+ZqexuxHctNk
RQufAqRkUtIy/KwHUWE6nxNGXBLLZN+9OlYN3LioKqSZxK15wzPH1h4UK6uRCQmRPwf8bOzXOFqz
bg43yMCbZLCFLcsiV2OlRsr4RXqf27MzQDUvmNtUh2w2uEZrkAkdBqZE+mgB2UDUqChTcBVabhe4
1zNERjkpXH6bzqkkpQNXWQgfGxLETboZRPOl/cfwA1HptHhwztsmLa6TCNsB8hI4OGGRimVBqUap
ZSGrENfj0lpRhZ9m0g2cb+Tq72haUo8wVsgEQHUK3xIRnFxRJEyZZq0evfevGyYoVyqUlESn3EXw
kIYkZZb0h4l6UhpH2tMXoFQ9gQVCTZBA68HPFazphxfJXiCeqJ8GIRlrMjKcQdoxPMFubYEetAZ3
ydumYhkphbPcuYQ8dFULKlKMwjbI3ipoqbN4+aLm2qO5edTcMUJPE582hIUJR1gGp2KsirxxfftM
qSpB6r4ci5LteXwJC4OV/EHa8SN14tTbvTxkjcQ5MwOerhPP5lMJRM7gw/PiDu+kz2Ci3z9urY/T
n1nh91Bkg5nrT2/STmQwCp4nn5oHMQK79whJ7FzP+TwKx6emSs6nx+gm9yklIZGwnhi6IM5VXhPN
s75SIrIk44LYBQXcFrZVRfYB1SBW7AAvf0vn4kode78Mp6NnZdARcRuEg2P6NRx2MK6w+3/D8ws4
+EoskuGccvf4QxKlacGkSlk+hUWrFfRz08qd3lmxvAnu55/6q6h9NZSz7bLBnKk6dSMkdU7PCljs
AAn1APTe2axEIYVTg1QjXn+QgIABuDM9Ka4W3S3swfxO0XivzCXULx2WQ4jS74UWZjKJMn10jbCL
Z7LIu717XC00fb0qUbzvIPtaNaLIX9iaqZwuBiEQhMJ6tjanyIboLQU4+MmxqStXxTrhuDqp2qYq
7b4xJCaRqBxEtTKWP/qiTRpvem9QQmPmaEEt5kUTEVG2V8lOO3mD1oRbrkJsXfJKv85oSzWLUg4C
rR6Ank+CIq3vqvyFkU9+IqU+eGmIkK1TNwNsO1mxUQ7lia8ugA/EfjjIIPXt7fP2k2uzK9DKmOPR
Sd9Bcn6B2WT9Ct+JzXPwiUPF5eMTgSWIltpFY0NgPeCFfz+Ms2ZWHnzpLxoLVLmQuG/ZFBVRcNDR
NzmoPNgNfoTEK+8vRV/iF/ZOM1mXkJpV1Lor/lcdjkeZ1CIJN5FicRQWKA/V11in23QE/xDPDclj
UbdrCKgv3rFESo7i5eZJyvhrlcegGWu3qry16Aw5vnneX0kHn2bPK29BwWVWFKstdHjW7SiUPeeP
ZbYp9vT84tvmEmYJrUP8OQpo1pPg9r7JcuBcK+GsduYgMLMm/njBJ61fVAYFqXgdWclUDfBFU5HE
ulyiyf0TwKuLCsmH4XgFeokFJ0uxTQGVc95EL+o9ki+F6E7AfCq5Ev//LiJMst8DLjQ3bDTPZ18r
jYIp4Dkp2ESrFB9udFfiMyIwjCwTeaYdf2/VPLa+rI8qd9QNWZMNmhfG0knMvDY9Gnu28pQI3Vx0
RLykmCyLZL5rXyQbr+YPcULWwKfH30jHHYIZuHRrd186IghA6fQKddi7OBBHYe4gCdrqleMYFEy/
AoGHzb8NNh09o2rosF8KnihvbmSLbbUOiTAxuyoiDou1Eda9L3lG74+7DNdq2MoENfv3WVMJ+tfL
cGlxcScfD0HhuwpTwBUIJZeegzuDi6nhRLapuV1ZDALsfYFKxesIEQ5EiWW1PaoGiNiK1sP1iE6R
iBlP3X3ktHM8LZC3PaYY2BoOBwWwuhVZ70+c+vAsdXg2PNz89CkS1K7u+KKh/4AaMjGP/xqWOPUe
Csez7zLSseWcU+q6WXAhOWovCfdQiZDzR2XFJI3XEWUEejaDE0IIwNwRef364luCEB4gTS95Xbmj
YG6HzRr8DFA9SvAwDJxbDK93Ibar+2T7AVNaVvmHfE1gI6bzT+vSBKrxZLF+5c1JuDW4WEaU+oO3
fAvoyj92QV0+FLZ7gNL+0s61k963By4HuEJ9g2ILwZ7GRKkEUbJDDYMsiL2OBcUMeSSEDbioKbRW
dDp5E+DJk2qKWDb/LBWHVzKfXfBWxmgdYUHPnHG8uHQFnMNi8qOsbPeGEbnXKpb4A9wWsBlh1hTL
AK0ffSXpJJN4OE6jLpQkM8u8KfNx8c9/LkcXuFiyRcL5O7mpolEom6CxBO5KM6tFNHRFu9+pBoDW
uN+SNuwQtt7aniSSZeUj8gAgsSWp3/a0Qt8w1E8Y1NJPEXTt1UM7VCe3X4Fu6/ccrhkxQc2pbBn2
8K3H4ZQmNU3cB7Tas63E1gveaDV7D84aAGMr9lcZoRBc04klryDZ4JKDCZfAXsXBucGpxepF+C4/
YFDWHBSIyKnhYikchAQIFJqcKimTf8ZZ1gyVkG6/7+3/rc7k1y5FXKsiYCaxlT7hdeJTUvilRaX9
z7GgBB6LfDbQ+yLrMaIaLa9BY57TzUWm/alZaImarEGqCXaKqtHGEn3m7sNfZM2cVFXaQZkjnGZR
+tyq4jooEcsR0Qpql1FQzFCb7tC/qAGvvGpR/9q+8T9/7mxHl1NTOIrOMoqmJvFVxfRboc2oETVf
xPbr4NFXsBLuM1bCR/Vz+WHDeSKS78L9T0Kzpq/Vog/D2OoIGm2mDdKy4KnoWkIp3n//2ksyz2BW
sd/4hG88wJriD8V4hrozzndn4rAzIcsZvQnApIR5OD3PQ0NyqqN8lfWAZj/xexGDCYPMcDie6LSp
j85yxkXqUd8NLmhYIWMI5XexW4AvOurgPfYHDgPty1N8IZVqKSFVnBxyNk/3bXHuIxCpZJJh+FIq
y/sLrSW+AA5HqJU4hyA7+562vtJj8n7UjufRGJwu1wVsi2EP7ac8OPt+WEQi/hMbD0abgBjTSZy6
Xq+ei33S3zXLKrifhVL7FDV/pAbntq4DtkKtlnVlCnhQj/u7qjuutKP79KvM+OxRtGPTJdX5Dd5x
yKii+XrNKU2Vgzyh4oqW5QrZhcBERAjpGnU2uK6B9mDGXPVoFrO8v2eO8IhOQ2tyXuzlYR/jCtyB
RCT9fMPt2QM/qt34GRzdSVbgh/CeIHVvh+5Q6slePRvtu++USlDHW/hmHsUSE1TKFCiDo/r8Utsk
AmDfQmpDKWGd4N1NRR/SyvoF0H7h5xPac+EDjXJh5UDDVKcJOUU8WuWaR9Dup7IvBKjzS+hE5iqB
TrywnyntwIkxG90UClL2QRvN8I5RUhzGAh6UZM6fCxyQBriUeI1nnucG6k+FbaI4bNbYETo/hhjZ
3Q1FXfaEh2IDc/xA41zPz4BTd69q6SsB/ic3JeaLgm8B1yaoxFvb94Wi9I6Rp/+i+hA+RdiqGw5w
ZKcaqAKZyZDLvw9l2Q/fu27Mnl5BpmvFfnIZRA2mUggk8OxmVlR0jTxNxgnpSiIh361pCYoKJ1Je
VOpmuM07KSe0VlhSi6e1Hn4HbYAeiDM4NyA/uMLPcyAvAtdeWqMzlVkVkHdu2UYQlkrJlFKOsSJP
oZCtbEIbl/dWNeCRUn4pPofDXgmVlD64CEq/UithatzXV44HDJ2vb0E8dWam8hXFM55OubTZzmG9
9jYMI7+z9OS4xJH1BP2uelDAGA7xwfZoOeVOIBG/lpdgawusUnz2efXkl1/6WpOKa95iwXScMvs4
mzcdMvLX+GY2n0Ckh7MYYXcZN3qXFw2tJ04tMovjNCJmRqay7XbumrpGbs2uDIorhA7JlJowTdg6
Xdr4Iq2Puv/c6keXQ5tE2MIgvjb3Poo6wGN5EXmvsrRasDELrXX5nrNJB85vs9TaXcE9lfaOmqpD
Ul7ho4v9OApPniKdYDHR7y2Wlkn7Ch29ZpZU5vI+OHQaCWyWW3ErZKXrVmxO89vGdoRwPm0TSTHE
ZaF+PomL4wA1VSZI6L3KYEIaUeEMjayAN3lzzc+Ys0mHqFhZ26DiUNl6tctjQldcrAH9lPKBxVKQ
wFedxYMYhkrkTUVv/jpJAN15odcSIEt4uPSunG/Jw4hIvtSo9FW8aSQJgYELfd8kWAs9HkcWAxMX
v2wNNWMlMQnAJlrLEzpSfnWtSHZMddPHGMcINEMYVQxqLffZToKx1xIj32Kqku5Stglfr8ulfz7s
57/DstAeI9185W6Co/xpSPiRJG90VF4J1Q5Fxk4bJNwDbDrv2tqNYNJ28lBeO9fMU8AoQpZdSfbe
iwW1AZtXEs364l0AzAcu07xfJnkEX9RiwzuckmaIPYZ0zpX289waxWveBcsmOZTstD0S+T9cEFYh
VbnV9lb/pHZPYy27UDzUOO+Ij4rvcLetUIC/aKGqkXYvCDndoNTXRxGINeXploOhGq+/JJfmKL75
iZLUk2yIoC8WzJ2/2oZiO2rsNEF1+82GTQ9H3s81ItZ6h7guyWxxNDU1R93vkhc44sNaUOpDBql9
/Rzvwe7aP4uzIM837Xx9nqOxe+nWYwBO0sqlsCPlTNGa7HXWGeZFewdqThSb4oo7AQ9ny0UPbTps
SoTJkwZMPFVzx+vRdxBMhtvJXUv+8QYLY2fRglC/L6SlYwTf9QVjWDbyjuACXYJX8FlrIDWadgE6
dqWRqBLklOYlBa0zS1sU9QrmY3zlg841nv67eMXoQ/XIDeQAtmWndODI8uesbnxWl0gc7J9Af1FO
ZSkyCEaO2sGUWM269oydNHH8WHyBM8Iz6JVTuU3whIgC9AhzWXAO7I3+cUuz4I+YOskKLqEv2U0p
NBpWf4zsxdMEV4WLZ0DOmgZ8FGiTopuOFzxV1bDaIKi85iPskvQCCgGY32ndCyusnploLOF3UqcV
4JHlT2sc7r/92F735mQA51gMAvelECd0d9Xm8BpRxLFgErsX2u+4I2ZkczUEBJ00BHQIyJwYPcgM
b719zjDWrzYpinXzfIlNJv0/yPysrKKnl6uyI5FjbUE7HXL9IfsxEF7n5bae/Vy9U3/VlYle1y+3
zUGMZksffX5z65KVYKesMJrrhqETJX1w6ETMSZnffVAeekY3weTZsjs/owNwMxPY2xHkUMltu69A
Rt3XE127WXW35YlYOA5kPvImZnbVMspGMsnw6R9Kq+mnFt34nRrxR8Q1G+l8PcEY35YY0E5Yqpg5
irBfe81deZEdAGnx0dujHqZALXYJVb/WQZMHN5aT32STIx0X/q7+Tm97LpVsnESrvBxWl9PNkMcF
3mMRnKtQVjZSqHjSTl0gCwRYDAINTZ/eufs+kKEBuegqJg4TWLsg+4ZY/VZUVaVkxhmqhXlE3IML
HGVLmYmj9ZVeP5drSzknPJi4qXOpxbo7NLagLJmAw6diUi1+WdCg4iZXa46SueLq1DIXLJYD4pf2
Ov1GOKWHEdNqa+yhrcmMvZ8OvpioesbbyGgAp2RB+PaqpdszZSbkUHQevggt/6naO8JgliFWa16M
HJZhOAwdSTR2cKK4L7l8YO9NH4ejEvfQDfYpbtbcYsbAN9DE6hNdUdmY98gKhJKep26ZqWTPHve5
Tw2fHmMnC8o9YOngjm45GUXrh6Jv64g4xmZVr9murelcP1wE07Cay6cVy5IE/6rs6qfp2NOrqVdl
jey+VbCNBj8RLV99x8DRvhkxrA/BIoaWuacN8rVHtxiYKvX5IGss+1+1jxuVBOzQveWTzI/g4F0P
0M1rQtaeae6YfYtt9myuFfVDsSltjGEcbSAKiAr2Y/LbURSI59an9OzBE0FlkcMJWNTvRKY0Bq8I
TzA4gXlQq8uE9t2Rm2cSkdNYohnb+2nT4NMf4aRC/Wqu4lEDg/9vucDeeFmfJh5zppSN9IR+92rq
YNhJ5volw4zG7ku4TNZFaKjwqAv/ljOStLsZ7YzFv766QJOxrQ9wcVIf/i0wi4TZdr3qajeswdgT
qLRm1slGkzHJe9E0vetoBpyAIoRkIgpGSLWoiu+olTcKM2K5AAq4gr+U68gt23vwI+2Mi6NjLSyl
hX5RuGfn2KadmV7SVsvTdTmwSDlxaZK0wwTaAZ2ahohb4y0EHEbGbPFDVc63PVY5UVceBf9DgImB
4VsvpNqMPwL3/S3rsGjPAw4XQPf8GTD4LIEsieohSxvWnu/mNs6J+7xCIULs28LqxhG6RPUxvhb1
GxjLHJsyN5JOlrqE/wdJEUfsWDEoKbfTwLLS+3RAtgHY5DMslkvtKlN0YmgQApxLjI3torgsOOxV
Z56muk/g3v6IigO8DYlxiUh14STHWeAv/aGZhp4ZB/wg+LptVi21nvAgUoGp2dzBUr4QaZjGt0G7
TofJVB/xlSuH8XjcTbD5gNmonEU6DVPHJzcoDxaXkVTcQL8LLjo7/0HEkiOXJDqwNs6OAQBs1YgC
NH04uak3N6owcBycdxqGIaVHnxFRxBtWrXdKzWYw/fkeMrn3Fcad1zAGgdYcmj37OCu8w6iMv+21
fgb7SIDohLFpCGKbGqP1pX7gw9V+gIcvapDUuYBWeqZ2IBqLSUf5zhrwcB631VAIGMWwmCE8GOOk
ssfUuEGF5TEeVEXf7/0f4bwOcMkAPg2ODxrRc7AkGUsq0vVC1XHUXYrEJ/KXSmcbyghnuI/nwSaZ
at2peXxLOjVPYIk7VRD4MH5YUJ5dYVviTRDgJnsAS+R89+mn2WidHQu4fWb92jjIdF1Sq3jVTXVs
rrnnNGyRyl7vEca+8dW8+j1QrSPdqRtmCBLuwXYNdcz8lnlnRySJGH2jdkyI5Od6zG8DWgVbtKWL
o7ilbpxazgJ7kvXs9QjCp8xKEJAIaPELYGoWFOjhGI9ORDtsXRuweRXwp5CEOHpr4eXRahj5KfdQ
6RdlKoeWTsFsnHgCGzyLLXNOuxQYtX6XtvzJYqeRC3jXadcuz8H6TjHKZZhnA//yTL+/wO94px6h
Xj/CADa/BmhTIYJuTQXSClISKgDBVgA7T3f28rOTWJJ5J0aqJqUzF2AB2ZHGRAgnkcq+2wZHCmPi
F3SIajp5Hwt3YEHMm1+6Uhk7fN9hBy2B3VeY5WBVL8yGbgqfiey1hA1bXozyRwag15u5zUrnX4id
OZVM6/x/qUeS3Zndl15svSq40QuBmmIgZDU4F99dl2Ke19DTVxCsJqzII2GViUbbgokY+II9RGf4
Ogp9qbR/f69GnKdI2ooKEMu7H4nRqOacdWTikH14Btb4DdlA3rvzXegCUtgdGxOcoF9CoV0svZl0
NVxr1C+xmGau6Ok7HA+QhyLVRaFaUu/CxWnhYnplViMhtOipgrVLW4DQOa8dxjexCWYK9e0TyH9T
OoDe3nah7JdDTymLtYaL3zBso/8TfUPR8gR4ECNFPuArmSuVuGP63NQKoEVjJ3Cvj0AQhJZMrrKY
A3S9tSdcsoj7c43ioGJG7oiPsXel0XFxbzxPNvF3eX96ZOkvFynng0rafeNwjdpxi76f/DFnrnf8
XgEoyywuo//5wu61RcdgU9896Bd1WP7ETlK2yHiB/hwrvHTTawQYOCXppfwEipNvNWXnZ6YR37La
upAaJSOZvJ3qdgu2OQ/0IVlPrqnOH4FqnWERC23DP13V4e4o7jkBdml0fEdGsbRZu7vnaRwGrh3n
tQFMsKmdDPRNiM2yXXEjVHZB2pPioz51S7ZNfO9JZ6eF0Dg37AjIF3KQurgBJxxB+2zfdkmBfU3v
Y/Lt4ty2OfVbNk8uwi0n5f4ZIP3DrxwsJXA5sobsYz7ZlbgmAxwfIT+YcCf3SVERXW4DfyfLGYlu
a8aH4pPLM2RIqYxf7FJW0vhpkZ224aJbFyCsw+R6N4LFZDurGeJr4i8S14QMr8hwxUQbrfhoYuBp
S4L6yJXgLCNzOTNv8MeDp+EnacMn2xOGWBfpmZcwmJjW0V1GnJRYFfSknthQaKxPpRZf2nFMjbW3
suJ6fhpIXjCMp6WmtlUt9qEVo/L4kdRigi6Hi3fDBmL2Fx6Gd55EQKnN4BrZ8jG5A7am/PaJCqd8
ez1fRejOIVcE4gu6SGV3JpOQ28BhvT67tkJNXF+JwzL1lSYuV+Dr3jBR5wcQBcYAQ+4WWPY3ONYZ
ZdhcJS1cx7eW8yuQjl8D4jlXMph3jFnHyFR+N5e3m0ir6HztkMB7oOhS70AnpY67QYqh1EdfCEJQ
2WLpnW/p32FzePQL0v4BogmLwCdK6MgDGSqSdKVsz6QKuko1QIcd56YPHy+SwxD2vLM7Rmb3if/V
YhzcA9rUwLI4nWYiE8C3UMaA16SrN/qI/4iQUxJGnWtK1buYEG/RgxTUBnkkQS7SqNK7/algCWCU
7r6nMf7FnsIR46wX3e3nkkovjMEWGHL5ud8CQZhrXMkDPPbFLp0jhffUyZtvSvbtUrXZZ8yNrs7N
+8gEy1oG5wlk6r805Yh/i3OqOVyyD4nZXtRkKWa4MnJka9Y/So1LaneljlRtUVzYrPvDxqpyrq3j
3cU1tY8aA/PQjuTmsG6KJwrhnlwYkgSzldbr0ujcwZLcjeOXM76XclmWawSPP44OJH9VgwDKopXT
pzJ4QVaqtgalFCjrXqtIdv22MejR47CrQIsonRVckTjvt7BsqteseFJVJYHdkFw1N9qQKpQl15eK
XBIdLx7RxaoXNmej1jx+Pesbw0JkaKt4GH7wlw9RFXgY9om+c/+ebE74AxMVtxnnFfPQhtkKS5/5
MvXwMVNjDH6CAG8rmArmmrjW0a56GF6I7xhs7gyneT1C41Awj6paA9mCCFLl6NROAPyNJxKKGRz5
7dEhKPbhOuqoxhWgO97PFl4L1UDHi8byr5QZpkVqQjBZWr/PFw5NiROS8xm2BUPQVWz5QkjcF8tG
4Z0OP0c+P4dpvygnNyveX/Doh+mLhk3b/IgZF7+J3IjAUO8PlXkZgeLfosazNABB3HufaVsigxgo
RYqpKJl+NV0GZ4lDVD56FGnxOI+CRdEnW3GMr31o/kj/zVaeqi0McW1BxMMjfjRrqxz7ODQPIbnD
BBo9+5qJ6AcgduKwwGu4jqlrP45nUIreZvngbFvMkyMQoXfCs09fbSm6VgFN4rFxmzkvi0Kdy+VB
plncomUjM5JUAC8eORhCWj3nmmkaMGT56LIrnWp6xaCWpPcqho33ME1YeEeEuoz2/ow1t5KATMBM
6JoxiioOdBEhxuWG1Nxl8iKfG0LlsCFU8JJTjBaNvvBmPn+JGJzfqPa/mIiIqkzt4jtWDzYye85R
aGCSEjUnUdfIsAPhMzB5TRYK/CiiqQ0sZTZeyBYaMa9AoTrMBf57gmQuktrK3Lm8TEcKL7aISZUc
7aJS/38uSc4tgze8mhJLNpHRKnjWajdHupSlKu1+W287dRZF6iYGeWRU4e9jbAzS3ECdSSyQR68m
Q/Qx9hciy+h3Uhv6isLVUGJKbCv33yxWFf9AeZujpAyekiEvCyEidiQhGEuPWDfgWFJ186uJHC+t
pfFJKmLjsviYpwD/1pcBzqCfP1Bg3PmGTHx7GgwldgQRjzGabPxWFsAtBys1BeCdRIeffDTv4Ppt
FSzxhR0/oawY6tkUJpkhxZ2lJocOCsb2JcW3RIG/FRUptaRx/FvrSj8SfO3w0x+LG+aGfyXGws5U
prdIgbwz+ylPq3Nof2sw4rUGfqMt5TQe6Nxo2TCW2sOemAJeO/ujcMgPgYOk8GiqNXKoMwCbKszw
uPMt7ywxhzIkUnfecVWSDmX/EB5wmhF6SLyxI3RR7i6vKWgOSef0/jEDHGLi221WxdTinBU40EZ5
H9jH7hVryo/e2ju1/4SfP3+KZ45XsGzPiy/3NB3lSI79Ktdf8rSjWW7hkXuFJAfjnF4M/tZL7zuM
/ULtbNGlJEjT75ZbR0RD+0rawyWaqUwIbadynqe7ZUxnEIhMdoxV04qvGUFvK1gP/OaRhZJ0HIm8
wq5AysKl/VkyazKcH25L18UZyaFeWNFO1DcmeZakHhey4KrZnNwNnGR/q9hl7+lzepLPoXWXpypH
i3wOUV7+sJBnRVTR5BUDS6+pzZXuDHBQYwroOvKyB3/4Ni3/Kp9aZFhjUpwlUaWyNiskjbDBkjPW
0PD38CxD6B2HNJU2bJDJmzRt2hRuPz9GZwOesamb4X/AsgrR3wNzDZHvv/43YFx03KPubCVnNaD8
RywrW4a1EX1/z/vBVGtO0EgjoumfN9K8IvRdShniaStcnzOjRdvYGNT6WT0ge/WiUdYJNMosOcAs
R7ssmEtcG261WxFJpbbXeQhYcLUVavQZ7RqyWXmdV3NO2Mj9TVBPzw4k3DN/yiNZHbA53ZF4lSGb
dmgHRoa38mRn4HKFDBScWYuMTn4VAZlGqQjx2bF4YQV9nHt3L9GGcnbmGGiiCd9s8QVKjnREs1z7
FKufnKb85cKm90hN0deDvitQHae2GkTikgsHRXX1p14uQbsbXs1Zo4/z5ySbql0T3SZ7apP/VzYJ
6oe2AIYkVPcGwlj7Wk9jkeAQbstyQA5OBAQRineQLGhisQ4R95YpzaZv1QA8lzSD0mZ5SRsGMN5m
auCGT3yk2+Gn5T0rAmpo5e9UFnpcp593/eaoF99xRT2yEdEfo02nZlnuaI3Hb6X8XVRwZuM5s8PL
fllcgpCdf3YTLVhRAw98SEgaKz8bAxmNbV7Ezs7ok3gvKl02PVB6O92Hn4ziK0+JMr9Eoj9O51FW
3nti06zs4Ba3/7IFpLTDSo9o/oCRArECZPqcslE7DlaxmqUdFI4tt5HDR09fLn0WaSsQmk4ZreZm
qcvxlKIbw1ztiEFnP2Rl8GxQC7RnPtsLkXM+6kcx4GRKE3RoktHJ+SVT7Qn1Gxh8wE0I7TeGUVgP
N9CoDZzdlnxhnQnbyHdrz3t50k2qrgDdR3+IzrorYtgIRPQ6V74IjXjGm+p0/8qRjW/ys/tA/28s
+j2/gbUJM3dLFfd0E5bawkbQwi6G2Q1YxDR0PCaOI9OD6+MMxzRy0iSjdjgMdD8BiIa1gcfIMxZQ
vUR+/i7J3wHh1oVy9qVHs/V2iVKjbgw34p4n+lEDSo3vXSbwORn70NqU7H0OIe5r628mACd0gWiX
+/B4LnQ7ZDGrDnQ0ZAxzaliwxjqDQbA9o11BjSuw008u3WKYzN7VLrAUFV8tIQrjNiww0TvAjP0b
5InvBc/pHfxPqFSqj7ntEpCibmCUcwO45hSn3KQgbnHeGA/axeHAtafovM9dgkNCdTupedkkrjni
gO1cs6CcqxACXaH7txESggfB3CYZM+MRgMge0kc1uN4TTTVRwiNS74Qm8DLvQw+nigRNW/DuhuwK
7RykFPo401JZIS/ppwIFM++HLeqJ8NvLU4dA068iXgHBOkQVa4kGU+dJrQdTK0VooapuEUYeBdmc
82Bno+9zmH90h+w2aZPsJVLhh/taKO/++e2Jegf/VvW2MAM+7gJwLs1Gn1McPQIIayvgulaQobXQ
M32RALaqOgzM6+zQblrGM1IavRGg72zlW+HouHsFkeIOeafcgM9IEl5JLKXp1cwy0qwLfM/aLZ/Q
ISvlXYjRMR+c269gGaB68xN26uLxgmQjsF3b04ZzRXJqSivVlTp7xxT7/63crdfJykEBdxLOeYkV
UcgpyQN8EFTLFb43tUC85AtzmgKcRjXsbnja2UhmCcrkKxf/lgO6RLgOgoPy8k6aFn46AZfLv6qC
QpGSdUF49VyG13Ef5NUFR5ENz/hdnXxqlaVqMsP+jyfDJxvTQ2Xzs//fixhlxmVbqgCAKOtN35Yx
VyKwUMlPVfMSZgVGWuwjpNeg67wxhWONpgDCMA+BObCFjCDXbFA4fGitXJwsS/nqI7wkAr5pWwDP
XoFysqdke1sMhpmpvbOnhfC14P+gtNrSK4S211QLJtGNqeIQrLfdLzFe6OU+iUOMgmfVEP4nKtQz
UWg3bNFXbFaIYE4BBKAVY32f3UMV8rBikEOGngp+NoXDeiCFalXUBvY2ZE1GMDL4nZl5ezKllA7+
LGVq1Gw6kpwiatJBD4rmKpIWB9qXl+QKm9EYAoRgezNQtWao5HXCpC9zOWIevQGVZT5LoR8zZBSc
Wck6pa0keziBxYgqpUTh3G+jkPPCwsoIMUMsMT0+5un91QrxYyfY1s14vp85Lo6TkW7vzzR3NMdf
Z2oT0Sy2yCO+jxnuelKaalFYnR+AV5YJ3BgfCEA/r8eAgDSn6AUhhXKpu3ahJ7tp0jY1RMrT/4kV
Q6YavtDfFyVEohlwayoRwkDBtGVCJAuFojW6tSBBywVAhk8qlFG0jsGx9cwSMgXtr/neqV9bV2Qj
q2O+dccy7Dbf1elwQCNTCHFJ0iT8Z++fJdf79FAGo1yq23JG85EtXEBBjh15RrSv4XO2AivkCA8a
n47iK7ZT4xsggFbOt6AIFZbZ914lx0v1qUbAJg8/SV0A0z0jUmFDby0dfcgJJagwrg45lggsjlLr
JE4h3OZ7rb//QNFS0tk8z1uMWK60mCKZ2mPwKYjotRA7qiwzdOoxiZ0wCVwrtULlDtTXq+M8qADD
037zLnutakg5Fy6y0BSvtyKGvmwGwRok83GBXOJMsL+OfNaeGdYkBc37wB6z8b0B6o72rj96iGOl
21UORPoAVzvlmLn7Kv5pfoSLVDsvIBt6Haauykk0V0I1A96Uxb5HO8xrSx8SypeSHGxfyeeWFU6P
/vV+H1xGrO0rrcJiljw9edY5q6JEAWkUO10dhSMe0QOUuUE8aGF7jk7nxX91yfjWqgd1zLg5HHBM
ebXCQ3Jgcnv74xUon0Ixvr+hBcF2LYIcuLdzZNqqNkFlxX/BD5ECUr0cdLBHqujZBq3EwFtsFfqi
lfQzSUDnWKlD7orPf2zuRHtasP5djdHS3Z1Gu3FADMH6I8PRe+OyOGZF1PJzaeJjKn3G65CgueQy
yQ8lEC2r1fx7ndCWHzUv6ubLH2UfnBN/rKl+QAdyKnhS8OD0wcsGXwUFPe0jzhByJ47592/MHtGb
T1YrYOpEPaINKBvtNLX8vD9hoPEwi3xWDOWZ5tWwDF0Syo7CzCsV+JoBdQU1raGFiXjMWPsLeNiF
ChJOb+4pzMdFOmEIsOLLbk2J+k5WAhCw7G3MLCUzqNwXTdexL8wfQWGPY8fTarKc1oa8tA17VMLn
6S+UjHwvSgpvnV7yiF8/Ic6HAf7ufXeIS19J5AD+PWvx6HTxY9+4pwBmYd2olvCiRXI1HVolVaug
j7QEPSqtKoEMy6UXu9vUxzL48zMHWzLazPWNAq0GO6kF4V+QWqxW0NYxkRlG1aDcuSewBLUOocIK
FC+SEUdDiwjIjYaSAZvVMENg5EkYPpW4+AH27vwEMbk80/Dd4hlIFAjmHMyac9qSNFZ0c2mfq86H
FhYeLE/HO4rYrvmBoy2fcUfaBiO8AXejgRpP6ZuNOAViCnHhRNzg1BMuwVfARAfQkE4d35GVW07I
Yek3U23rZhWKQoPOdJxQgS/ImDk6BIIC/TtrVcivdD4CcHBClTMn+dET2MapkVIRmT46Kjc07TVH
6DsyXbr61BhRDRgHPajqF4ymzaN6u0LrOjOHhGicB/Q7ASSb03cjmshGyQlVGTcItGthOSzcrP1O
RadH8fYcCU2r3JZWrGnK73AxIpn/LfOtaNcX5z1lQ5Itw4FT17RylyWkr6veG6BZybXf7xsFG+cl
pbO/Ar9DnSOmiTC8MqMMBX0YQ/U+VpL1TD4rmigvksa/VDBrE/AOtDsXB4gHsf65ZJTtGOrmMFEU
/pQ+7cnvCfy1OCLb8n5OVYpLp6Bclu5SG2e8bWm7gqQt9P6EmCiXVIB70Bnyq1Aa6A8kJwNrTEDA
0jDAOtIHrBX0o2K0bwdDX2u12KKdNsRCR/tOxlX94cu/yPGVFx/l9GTj5r8nAN5Zr46fuUEt4YJG
LgPzD0SG0kaXzTPsvAWswLz51bJG/L/Vw/ygdkUewRZpvd14/tWJU1+YdZYvSnqiU5ZcX8/HaA4O
KFXCRA2dboLwtJEpW33xVtYbABT65n8gd01kF8sY/NyZJcJujRG0g4x7VpjgtEaDfwD3GgCIK5iE
9+9vxgyxQVgSIsXHshjnhQZshMhhtLwkWFUdn7t6pHLNgi6l+X1FmwSO7AjvUZ+33bH10u8dLNNX
zbc6moUEH59I5itZaFg8n20Al7y4Htu9/qJGM3gmNQD54OVU/8uTzh8Z/qfdbRjAHSlIatQ/opLG
M0Yp/ofkF8Msvj/hNCc574BS5+MBFC8wj8+AfQerFdkBvN8Q+04Am5fm09PFrIYraqoV9Q/VyoFp
zBPJbaXa5BNRpg9cZqp+my9XDYPtXfLI6eFk0i00KGKzmqtcXS98Pz2U3+G/tRbIsDnpgKwH4WGs
CalRYEfYUz4x83HEcQxUB+oEJvgOu9wuylimIyTg/qpZjqbgPxKeNMlZnhYuheyu7vqsWN8vknET
OWAEWPUoJqcM/D6qUJtRu87yGD89r/kC/dh3bpgDaHQcbVNB/JORbea38TqWYdOI9K8C7KndpTEj
7Wc+L/0/d/jo7N7x784YJlpv63Idw2HHXv7CPC2ycjKUo2W5i+QNLiqk67AwirZp0pOf9YBXSs6Y
XLNKNRqwCycFlq9Wtp9wR9RIh9G5ubXmt+8igwlSmdFEyue6jpVUkEQbUfNPaREwLZUnt2srvHd1
r06CZbjw9bt7j0sRG6SzCVju8DF0jVkEU86OQugSgrnvlfM+FFh1w9hBf+Zf0RnejrdUqLHP4due
eFlBwwJiJ+Kl0qmTju6K0PA98q57SSI8pY7q3F/MkUOiVoLiybBqRGSZQBCeEHFeE1cslg7jnKYI
kDpjYgzvZIWLg1GnbxW1d4A9njozGlWovrhpvBpaTjUlrwpcEKvGYoBYDRR3fiwyMGlIA72rnu7w
BJUOZJy+HhJ/D0x49aBTNV+q276VJc7YHyQDjJ2asiB/vYEcgOiWu25X15JnfnZwKh894oGyJ67U
uYuZyh6sy3czNVPTQ5N9uA4AZX2v816wG/LCmb9SvRfKQSnDjYSosEDDaEC956QFT4Pw678fpXVu
KRAyR6EWU0ySPxDzGaWAuK6XxEkrN1NQe6PA6e4ifwRlc1hZKKoh7GuhlpPnYASWfdevLzr0iGT4
8UDAoSJUmB4ssBqE0q9SiFbdI42IRy5dbLTPLGd9EeU8WIoGpeDuM5IOYLBbLD4lBA6ghmPWR6X2
Djd4f0eAl75xrkndnhSpvI/sLqeuUKk59LgqkikrqMwh6Tebzmfb+97UPZNxE6u/qKxcQPih5rGJ
9pP+gOvyDalvhpiywlJCGG2C6rXuw6E72KjGtFXWht6M4t7gEyEUwKd9PB/3UKT+LCFhTax93e1Z
rQyWqi3gfoW+VKVlQ8/4yr5ZwS4FskoUyC2H616zD5dPpHu8IX5OzpVvpRQxxOMw8sABHLnb8uWB
dyhtems2JuFSKxRcQRRL5LrTObRm8zPeA9Ey8MgfB8AMo5wG5qAp+NwHjtV2aFqTo7WPNQp6ow60
whrDjV9TyWcZKFAW20HPrtddbBKgJVCBlJud6b6JPOFc3UnxQZMc9IpVu75+N1MGI15aPT/5XVzG
T8FFclX8b/fjAvjnejgDB+ZYMpR6YVOLQ8DvAGQw7pKZYJTkQF1+10AnN0MlySiq+mh264RmjCKe
d8WbFEalVVJA9fGcCUd+E/kFjcTRCoajtASX5HbTrS3vvIYTHUkuXa7M1Adj1fZoLFWiROXOQ8nA
HxWbjZsIkkzeObk5+W/ER1c2SiADQjNmQKBiVmwcWFmPqk3dnwFSt1xqAWSUVET7h4gbYOrNyqtt
xitnUTKlL0ECoh4e46JYH6MOuhtElXXgMgVzsob8e4wOso60YmboVw2aF1RSJTwGwrL8H9CueU7l
dqedkEW8FI9gvJq6mW1Pw/zJGRn8eInMi0ZPwgzWot6JuroKnkeYtqUDxQW0Tl9ktGLB52y6nAAB
0We6zR2JXe6BbYcwB/DVMmdyLsCPDraHAOT+rudH+S8yS+Yv30fMnVR8mbbXwdAGll/Y6auowe0c
UqFDm8cm4tw9g3k8z+RrpZHpz/xS2ThXFo8ClQHbiwtmKRnAXRit2cJs2NtnkL6Nq4jRZ1rAYJUd
RLBwmtnmbf+cP9mvMTOi1RbPGv/KyA5xR65JAoB5lKxy70cqXFVgHNvC9Tl9y7ynZfZoVN6r5gEV
FZj6Tbdv3IZzTMqcNOdGYGf3/V0qKQPJTihgZytWhQhXn61cEJhsT6x2BD/OgnW3aRBjL4qpLXOk
s69LZG8s6XpZOwKDj5WwlSeeb20SEhLZMqHvw0P7oojy/zJDDbkrFBYi4FyOAUo5NrFSmWar71zV
jl3IS2ZZJ8rm7m51GoBh+X4gjryHsoRX2RCKNeROzCvnJuNrF/Q5iX+QDLGEm+6/Mkt9ejLC6upL
leGrVEo+WZ2d1OiAAa9/Yh5OOx0S9ELx5EGcA1vX+WF0rsmFbipC3c2QkplTv5WbwRjp2QdNclgK
wTTm/KDUebpssDG28SMoUGR0eSsZCeDTzUwE3OGEpRGTCzJlrW3+Q471kQ91E/FpgPqCIlM0D4XS
6q+mF/42m1veLYxaVIpMr5xE27YlojTRJc1cJ+Qw4iiOe7HkMURx6mZj3Lk7LoPdV++KEP6BGRhw
iJC/y1ID/LSxF1xZG3h6sCMnR3yVDLCWAJKC/j7uuvnTl7N5mqEw1mhL/Eq2SKS3vHUOWTb77ZAk
uIlUAgyuP2QSYOl4W5eqvAwmb3AWCqtUqbDK1iXpmnjejXd3w096hhu3L8Nwiwpuh9znWPDylJsE
5pn1TJDWU1DTbcCYjaBIaVGeyPXXQgvNyCBDLkVbuAmcF7YkRZ+N/B/LEouC3YvB64+i/DCzyE8A
TCcru8P98Ri2IeOv2eKJdnuqdoxlcExHbExdwPaWdsP5e7QhSnRqMKVJjiAWIp13hhpv1S5XebTV
vczBLM84K3yz0yYbe0cYf8aTfaU/bxFYUjAQbeACzY2dDqcdggLsPAdrWTZSn4JImlw+e/l3SFIG
Zro+DVkRZk1iNiO4jkS4opJ0+87UpVfL0CsFbkHNUHrNvsEmYHoE0vSiY9T9TrFKAfe21vrZFLRw
CrfUKXAi9BlyZWgWVTf52vI/VWNzL2zfJ//liimIXPL9tkn6EFjoyS1evzSOd1Ld2roGU+rtXKpM
YNdAitjg4Z+g43cDFWa376eP2Mu9A4eXLLVNtdY5ODeQJr6xX5nm+Jei4gZp5B89JY1VD2LqF/gY
9kycOmWkcwTkn/oXROGaGnZtphrwRUp9TA2khsNe0/LrfF3JwzGDgiychW0gTqIvZHl1jomLbNLS
I4ZpeHwtnXuG8NmWzKYYQPzZm/2sQokhfXPEw+as2HHSZCgYYz92J8MVPnk59/KFHby6rLRz1de0
2IMtLtYRGJWzsBcfzXdxVpm8w93pOdvePVadh2ykdBpcaz6QRh43+VBp9Ss2QtLWWjqr5BFGbKzK
iVa7ezMdSRjnOm8mb0ILmnmojggM/un4oUfbzX/pvgrFWetSk7F0TbhWYlsE7/KLwdS59JerXuJV
zZPVm11WUUwhnH5lcfUJn6qdUxjSxYtMEpB4dvVm+NiKCZ1ZluurDb+3MLJ7ZaI/J/yajSdv6wIC
AgKCJ2vQ6hc2s4w4lAUT+F4gQzgBua781DEoafSSM4Je/+sgvSQdAEcJHwv4iINagChrOPVlb6Mm
qi7mTxacDHr3HWss5AwCdF3rH4BztfF8fO6JFzg+jghp0VCiS1qm4tCt8K3jNBBDqUTkr6QjQNj0
vVy9DfWPw7A7gNF+mel5BPfSoUcjydaCxzJbnYGSJxjGENzLXUkAadL36C30k4sjxuLamNs2VJq3
6J8Er0rK82btYdSwncLkBx4AkaUJ7yBhRbkn1+kWHqJnFuvTpK2I5pDrJro8jh8zg8WFnl8isPJf
TnCZ4vKWWSFb5ywk6TUq9LTb6OHFItcRMMN47fVNyInw0Auq+vzlvUaIi3DiGclnluX/+MOXUNMd
dveiQb81uSH728y6cuJjWrN2uP9RI3lIu79EGaksNE5CJjKVQvC2NVWEtnfkl81Be8HKStR6o1ci
trT5lYiJGXl6of95JAok+uiRdN2MZpUwuAQyu7FAB7cdeEgdCxAGm5CXd9X4wFAvpI9aYwWiO1h8
ZOBzsLZVyfBuER0Y1xg0zBI4gfG1sHQaWaPy3+jBN1DXuxXMeJkRb0gk1e1M+84LIetViNs63IV8
NoetrstE2xJpCj7bhKFOxVuwh9OT9aeELdXk+zGWSIE/XEUlZNsp3SxBoUhPXrBtWGBQqZiSKJAZ
ayVavvyMLpBUU7+WNHrIGQk6arnY5c5/1ddiqG65xEmbI03iqRr10aE+RF8ITNIa+Leo5ZvV5sS9
J22rrWkXIAUg2C4sbOQ7ysAB3XbqbOaWsZta+bSASC4iOcBYMdWAAVwL8HJaOWjvtq0vD8M9ljBO
PfCMnPuZHqMRXqX6AcS/UqFhizmVCU/Nlpd3x8kDBrSpx/IaFbxQtfszYpvCd7cQgcCcIt3QXKac
/K9ofy8Lawo0iqhyqOIiXQ4GlhUilAWBYpZbgdR0P10mmxDE+4SbAXJqAhRrWl/aWp+NfhVbhJJO
pgW38JY9aDhyJlkYSYcEzFjADwhMPtJ2Na5EZYYUrXmIMyqEY8cINkf3XMoLC3/Pj5xt9pbAeZhX
rY6AyGXdLY9A/O5Q99x89ZqX/CJW8UHFfea228RJJWRsHrhKpY3EcGcx2vI7b9/npQABogbS5zRI
dfQWLVePSfwm6+D9k6hhPvW6/udqQ9Evr2A2pPkhbxx4Plqz1B9b5kJS8IdRN4XNKkJDRssbjxJW
z0rVHlb0DPvxRGHH6PRZQofHFNcoq/Pp1ot8IKt00A8pgrTDcHKtbPa5G0oR2QXjgcZRhU8GLS2e
jGb1umP/pds3Pbimzuou90BIKc/xB0uv8xirRbTZG5uGPWeZWQq+6F8YicRHu9F6PlT2py7Gg1pm
b0w706qUC3DCd+gkjxauErNsPzC15O11ZxzEWinDVa3J8WBT9TjsOqxv4Njlw95hWXrPP+jmhBz/
vgZ1FY0F6jV5RTd/Fxz5siv/Axs6ZISUXdoCBAm23G91AAhJT1aH0FPkYB40SvrdElKPzjWDPhOc
TVNL7tOz0qJ6J+SoRmIZdmRBNMQb0JP6oN2kzdcYIgujRVodc5NxzO8YLOXzwpI8mRlfmeyo4h6N
vHieiWPY9LtMiEkRAKnlhhZr6Qq5rxlwwGNTyCpY15IFKWjleD2+3YehzicMXczc8guPiTGcqWRA
FGLP+irsM6YtX0G6nWESlFGyLVLkUPeWhMpXX+mTAQM95HfMC/dEl9XsteEir/ddeSag7g5Drqdg
9vUHkFQ/NFrcyNkvUpIbFuxU4pLTXrGcUFD+hNzwXyy5Y9rQFRZ8ZVjL+eunlDVNvjnOdf/ALVI1
emUyRuOT7fiPLRi7vQZNl6ffFXRRWdtklry46GgoGBCwC4vH9TcnZMqd6a3Mm7j4xuQMM8loKF68
u7EX+Hpemk1MKX1xxtQPV2rWtqypIy2o21pu1E9tyLXkbpCxLYvd/KkGTsciGwH+pGZHf/Q6fHVY
Zth/pTlXH1P/zw5T28rMvRq07sgNA0iwCxS9WBQLioturqfeGlIQGXni1qIvqyXKGfAQOdtXhA/Q
MaHRX0ZAZsXlrI0kLMk8iPLJQsjHaksMABhRhHoUIS5b3AdUxEKPSAXgx7Zue6SjpAjAAHOfiidL
OsG1WV5Uef3ryQv1Zq88bGYaWroO8sidlmvhxCiR2QNAfsH1kvVMAXqQ9sbgIhVbo5lHjD+LjA3V
8y6T+yRSKLusbBtyHT/FmbGghMH1IiYezh50NAj/WPAr8+PhJGIHkZMq/yos2ZVWKd6EqGouHHa1
GhJdyw+LNfqhJgIoc9j04ibMqTLOMmqw6dP2k9jaX6PxktiZldEk72/Z9sX+GD/KTlao7VncJnDz
ADXW6jg6Xg4yy0zjlUttbCIiIid9D/N5s1N+bVN/k2OeDjgbVJVn2zy5SCD5Yh8nWN22S+5YPyFh
KMn3AoP0CrzXVKyXOjBj/PoUe+czCT6yEKhCbVGjDjZQmBToVAzm29wxhHOyR1o4irpnwsMLq24n
xJkqAcp7MCe30FHol7X2Mosm0RkxpYjkAtb0hnef5e4oWu6lWjTFgrvsfTgsh/wCNXE6X187Siq4
xQWWP9GWPa2NFLsvysdsgLiUnfwT/jMrsYu06k6SQiu45kbux0IjShF2hIRb7y5Sp9jdHtTN9YaV
NRH/mLVfLfJ1OHCmRCS3pDhzhRupUnafDNamnC6PQh/y78D5cewhfzrUFbCtuN8uPuGfpP1p7shu
zKdwuld1FUy9ntk2gZDVjfHRjmB2LitaNPAS5MpPfDZz3mtxOFiSc/8ZPSv0r273kqCXZsa++3/Y
rPnDzOXkOnad8s2afpvu7oDwxlNWX1EtP0zTGnl047ZwitfImxoHc4JWH7t5CjHv3/UafCRdOUzT
/fmX5utt1O3Lim28xVZ9UxNCBWj4OsuCXaj+ZvYopDvWvBA3/bTB80xK3xxVHJeROE+O9zOOeSYD
veqY4UZdYWeEgjz0kfJn41F/W2c4xAHE8kuvl/MY+O42raSWHsDr8VsYjd0HL3DP65tzSqaTswzv
rwEaLc5/Mb7NlrlEEH0iXTvbVyTKjksbl2iGYqSQYhFzEYVZtK+EvlP8oTePQM4rYl7n+shIQr1n
i9il+Dn9ZylFtiBG5mWdZI85egWE3Sgp7HqzQg67sWtiFknT6KApxb3ZO0g/Kh/00TYY0boCVvVv
xt3UHj5ll37whv9SMbD6hwYgl4oHsq4iTeeFdhTMKrCa0mSSx0O2NQbvfOg6dbJ01fiuASADxX0A
8k/XDxKFkXCjP2fkDEz1Ll80yz9JfInoMMuaR9bHv5CtA0bnKCn8GVLzRRUM3qYlCujBVDc6FcYD
4cA2UtMe2OqY6Xtyi0jgVbBFeXkHJL54AD/3BWLq3mK0yxFSJvo1IBx1eDr9zpb6ASXLFAm49ifP
4J7nHsDCdtZdorT9/aZUwyihbYduO8GRDfYdgCghMz2OpOyrq40wmQ48LD4KHC0iaeAO9hTpUK8t
nf1gzpe/bYit0mDql+qUGozAbUw8h61F+vopT8iu/iq8lppPjDDTYlu3/aoRidSxAxf3serwvE0t
NY8xSQaK6XPKrJLZ8+1J0d/ADO095Y7sqWHfmb5iMgFXETE95kC6yhNeet5OX8/X4rcZwkTAVMRp
E27QsEwZECR/X4HdrF0o+eVspRglRaSYTDvGmB3BvvfUCnRIAuVNdN5iv70Jlcpf9UHWagyUMaD/
Fb405XgaPOzRcnJWLkQT0fxatHDHd1u18xKqRg6gCsg+WkF4EX2r9DrbPbHi0QW9kWJBhhb3WG7r
EaO483DixRirHZbMGjtgMvpMV3FBIfqK1CoAxA4KZUfEHTpjo/CdrDTlnxZMptVerrX29D8hJ82h
kGWFOXVcMb1uGMNpWn4dCsTeW13qJ+6z02IDxp+pP9mUBw3BB44C0EvgHkvi9wTiNT/+1jZl+F06
0EjOubp3cU6WaS8PHa00rD1ycKDR+75dqDhWYWlmUXhmU1LHBLPolhh0OCXxMcL9Slyd7OpeQk5r
70L4cwrSHa+MK/XKrSdN8vV2aGA5Tw1pMRngmOfQo7RpQFWkCbfKxNu3tsYg6OvUQHgS0+LkFxl+
DaaT+i9zxBAWFs87t8+thTYWwKs94c72y/lKQYuvsp220pDLQzDY3uCE2cKLKMbgKkcWfe56CMFg
RzBDF2hJ6qp2ibdmdQ86oZ+9WMJpUxV6MsLpBr4UsmRPAo39rsXcdJY8m3RV9uBpHblMjDRYwVD5
flUi5sbzdOEGptGBj4cqnNAJ6DqYWbZ0gdkFiXZe5PeCGgm1aOqqYI8XV/5rsRmpqp9Ah4T6qTKJ
kwEvTdMD6Hb+HlmM7537MR+uGnnN62b512nxdnPXsvF0EhVWrt5EztiBaXwkwUHM5zqj2v62y228
Z5d4PF012yqVRHhNgTxR69t4YfAuDcI+KiYCYVjy6aVqzVE74Tu3gLHPnFe1XVGSxfvntsf/N5o/
hGAcYC27C9k0jjlgLiyU0dSVXdsVUu9vkMI7O6Veb7LSg2oxUIMM6e0eM4dbYxxE+QXP1paQPRto
Nb6uVN+X5wFa3T4PK2QYNfjF9Pvk+7uU7imyp0N8Mwd0+Dxxk0qWqwhdhRZFxv23bU1xM2iZOAjj
c0lMTTbEvXHdZX+HqBHnaetoIB1XvxihGA0RCk34XoVxJ3Tpc1qtQfOV15AdIqT9gtM4xw2AAVMi
hsQZziBtXvfTGBrQJbzSA5A67T4V2X53HAosDHmnmrXZvIjMbkTz5PJonz1ELBPEdC6WRnXSL27W
x5p0lCcFniSaTrzwXM8Ef4ve2iVtcY2DcyqLBMVFJeEtnoAdskZ1aYfzX10JLI4HZzUQppz6G2hd
uVoLi/3CZeHNIovcHb74Fe/VmNPekHZ2VJrMhS9xxANvZK8i9/lfxYSMIMSV7IH1hzH4LmLpkufp
26gN53GS9zpmxIXi8kEAqB8d0n2yqA+HPZPtRO/UXkquMbSKIB07yu2wuZeUIIXNCDfamvOMJhit
P2MKek1PhC/Adhb8b4vrVzqBfJpTYo+JB6dQRnrsnwokMhvpt/bGNWyFuqabbRsjwpPztNVZLHPI
N/0axpvL8dGj4waepptDKjYjHE7vKp3V9Sty2jXrhiOXfNd1me+o3gloQoJviMFqVFksrB/8QFpn
0ybul615B6+LL5Y1lnBQFT5wc/b7/icb8agJsYOEeb6gCWBiE+mpYS6KcWWWiA6PKsIaQzdjMql8
1ewu4UxGlj+hAXHdHxhRC/kEFSq64oGj2VvX+wBEdghA1v9oKfVjRhROQRDgPPCm14CKJHZyobzP
iplOxMaRRC5yVVoDQi5ZAbT6p0QiTpgdgFggWOfyMPtugnLAa6rh7+AWkzqUwXw0zLtpMNwxT5NY
AZkAe8rmYWgJ4rY15rlO7OoKNvl18e+9qM1a1EUNcxI7GXtCSTUs2OqmVTx420ZbGtPgYVOw88FX
ZKbYM/9nI4nttQGyrOyVRPlu4DGlosGmuZiY/kMj5O05Vu/lzftEnMbrYa9dDiRuQP2PRcn/xQXe
O0okFLxmST+93Qv1ysjDUz0uZdTB8PWhy2GgnumXHi7CZR8WmH0+ISiKGIwt6CUfZftDVFufJs/G
XU3p5768cihxUa/54jG2JF5Up7kC6l+XPKjqPYIUhHPmfvkQzCb4NN0Z2HdlQ1HTXvwiSWW3p3V/
Emlmtf+39eIMChz8dKLENwaWfgYZKNzSZljhuVGOGSXhF4I9TZV/h+YoMy+FUmJ4P5EwzlRb+P8y
tmM7ghwGA6krZE0/DtmDn9/9a2a2+2iaZuFEKnaKRVv0jFCuOd1hWroTxuA5TKGSJ1KYzGZc2hdi
X/SeEQWfevb/TZMu9s1OSCxpYXairDjnoeTC960n58zj1P5lYoRtdN062PxWQ/uryiLOq9xXpE7S
BFPp65uwyANT+Sie+dLsU9/KKXyW63Qb0sQLJXfxCyRi0JU1H/C9Vc6QKxGMRDY+dh0LvFaV7wDW
n4II5lB8SECg7/2C7f/yhCskiDqNUcPxE1f4ODiXAEMClKCmUGO9S6/oU97TXf2Kt5JtiYf2UBf4
4zjndEzrz0dMkzGAEHlStkObR5UyOyNDByR1qZCP7uxqXJ5h7Mhd3ecPDU63v4Z8ITXdJC9m/WnS
2KFxERciSJUtvusS7gpTjveyZ7R7+KTGvdpph0GZlFllKeqftSCM8p4RwPiy9eKpNTGIPDJoqsxI
JDfkrmgoilzBjpX40m7Q1G9Stdp3J7fFvqI1upznaVU0teLoxbXUrqVmQUNqZPOiPA60iHcUYKo9
wUkRQoTsSnMYZ3I2eP6UWc6EOz6MbqxQZ1wpZGCanKBoT+uu/nCdhAv+IN4eVCFYFxL9Fo7MshfR
tlzgdeCdinHrmtqBWVw4o1CF5DXl9f1KLfMRtqPzErOZhxs7LXhwdG+XXR1EAUrMUkN/gxuMJqlH
6TeUyXaMLEWlriq1Hfs/C91SbfDSh7qOWdfrbgie38TZj1j4uCsPVMLZPB2oFrlDJAKUCVu0BkpM
CEbb7uMmpNW7Mzvy6teT1FrPtBejISEOCWC9a0ctOMMO1fzBI0kEkmOsc3GKVA7T5NaqFgvmKNYf
WBOy/IrH5dYEV0ot+25mVJxku3dUb2v6/jyC07umUw+Z1V2rCrTE2eLt05z/4v8O/lrJSyQ61Lt2
dzuM2qjVHT9nc86MpOL7gRTeQmYPJjBimA0fy9DwteDgscO4ujgbaCdULoCouiNQjvsYNjF0P/H8
QhmxzBzoMr5T0dcsO9anPBktEaEHqZnflo6517Z40dXPLZVTgTDFCKW/vANH9CEvgm2sHoM0d97B
yHDvOKj0BsA3q2QMt1rZz1cz4yxD3jfQI/XasX11UH9sMzrdcvn/fOpY+BGCpwkUrXOAY9R3zFoi
0v37NGyVMO+Jwhf3WV9lZV4FZgfBhmxTt+r9JYMjtPnbO0Jfwmzzn0+JypdA3yfO+ha74yvuC7pP
nuxIvF0Xiqx7t3rbRqeE9NhMQGVonDroyRRjh4r23yhpXXLONPG0TOYoaDidUtNPA+e+bSalZv3V
L1BlYedp7davniBGacSmcTq10OmO1UlqTKgg911JNAKx/tSosh45CdwmdTGwX2ElHIAGsdAfxK1i
pnzRO6th4SlWeFkUcLLfJxcbQ4zMGq20kUEpyBzM3CQ1kEIRG+09PbC41ZCl5025T4ts7h2/BJR7
D8EyLkCRIk1V23l/vh1G1fXINbcl/TYgjKwv1VlXaBD5zNxcOdCS+ytteZJRmlxCFWImNZ3cY1AZ
kBlxxtNjljTO00RdFgHv53+4h0NlHt0xvx+1E27PgdqD4OHve48buwnRwP1gftpRVWQ2H/0/UKot
4zS5IYhQ1Cr+f2ZZ3764zb06K8ryT9WhkHzjwWnVGMQZieodQZpfSpHa62OyudZddjQ7aQ604J07
VckfaRb1eJ4siLe2PRYJNocvL3UJ4GAAgtBZfWx9X5E27oOYQTzou6i6oLYaf56c8COOvkJcjBTj
0UzP9i36wlZo2hLVNSWTcG/sN6gku8/NmdNU3NBCa1QMND2pryCGAwSVVGymSgohXtqGhGqV9qUX
YlaXwaNd6fSnYNtHv8pHcYIdd3pbrhOO+7Tnc0bE/R0PrlrBXN34ZYLzJd2YZjQ05tgNB40na+46
PcOwrslYIx0VHTPnEEqTxeJeRbxr/fUgdrKNs+va0cxhOXX9+JhuAm2MjoF8K5Fao5VJTviRsrtE
CF7RFMXUg80ZR5y27Cy3FADE/l7GC+hi+W9UXeu4kCRb3BzS231WfmX+YZ3AsCyqoBDEe4fEnE6g
rZDiIsRM5q4wLK+K4tBHETuisH8pAn0dXzTmkhrNjG7PTLDawb52TYvl8JHrXMjF3vFvLJJf4dTi
dYyf3xSHm+MAgyz0ascTSVgqU3FiPJP8JNdeFZLvfPwksudzucR71AvpFjY15IJYmuFUZ7ZGxlGd
BkpxtBnveGOxyMZqbQP1IuS93ksXurFDq2R7cfrYGIMhvVXwcMUr4hqDe6zOyqrYaUdHjrN5hY/T
XGMRphdlN3iswIWWDLMgAfWTy28dZ8vKgQvYk6EfJF5WoIHsqAtcmIB/skNfsTn4nXkhTr84D/Dg
Pk9vyJo23SG1aomkbYZ9O/8HWqXzWrXNanpGaxYoBIHwnvKhzdW0v6ewThZlm6oowZx3cfW6Gb50
Hh5Yo+VfLGJ+5eTe+fHVw2sdzn/byIo/gWI6EOdQideYrHTR1/rH5MFPfIlheAVTxsZxxVz92Z8U
4J0HRf7x7vZ4AbuR7QpA5nESUm4Xq9NB8PmCBmWb1om538+h0AEcen2ZmM60CMDhhG2cSNnPyNLx
CkBH9xNh80hQrEkxzmirMRNeHXe08CxBjLFZ7ZIX7O4PHt+jOHsuV9uFgE3qB08f7CMMni9AWq5R
n8om/6BIxgn4MRXS/7ubpBtG9yAVpOeX9zBMm+PcNhgwKIGRmSfvyaSAlnpNx2NmfvVVOgsOEoe0
hRp36rrz7Ai7CGBeaasAKiZygRV8N4DMzoC+4APQn9YzhI4T5Rhvdg1IiaHq53iRtU+Btli+QaAR
Q8RGWRFbMlCNqTjYL/3UdREBF6kMhbwcVNm16B9f0zCDnD4/HCdUnqUl1aKdLGc6fGsw763Gbq5c
O5FYEjINpBIqZEzxYRS13fmh4o9Piv/gRIMsoWQXm5EiRwZimZFm6fXrpIQE7hsHjV2/tyZmc6uQ
VuWBUYam90l6A3eiak+yzHZ7DI5KQfsnWdEOjsN8erx7WWHrXodSJ1jfLGC94fyPAV3FWAYToKZD
kqvMgZvFTSIJhs1rpgkz7bIGpPfveRrE7vuDVoKNwlT25ETxseWB9rRe7K5GgmWqc+b6YUUb+8k9
UZhGFuvXiAkrFvuk2sd1JG+LS1TzBN1YqvtRcWbfIyfzlGkliTIcSIhYm+OMk6c0bezlEGlsf1Kg
OGEAiuvV+LkaNbE9LnHrNLtGA2cKfmR55IAi0EabBIrprgWZVfmUU3y94hsHDUJ3IhMYP3Br6vYP
Y7bK0K6thzVaUhnvpPeIPH0mrZSpToLXSVfEBWdwTxUCPJQ9GoyRkIUvhNMfNV7Xw5/WCMPWYKLK
C9W0nlk3lAYXB+6h2RsE4Rq/eQTBA7uHnHc5KbDZwo0OMnLfqQ33Qh/uvaIqqHJPQ7z8Reo7aDQR
1uJatp8M/uQVt1UJrtDSvF3KrAvWZsWT5jlKWRQUKWlh8jb/LhDM4f+mdrXx9yCNTUggCrESKkoJ
pujKIT3Z+Mm9GPf3gFsp7hrmnqnW14SVoFS2UnKJtmRby5EmSSoVx5l11p8RnwrHrTKhaBzVM3w8
smG2trMZcI1/x1ts7erKWVUfZZHqSWi2TFylXlodvlrftYAJ2bZHUa2Pfb0IGSbfBDIZxQk5QPqU
ZPXm4bVnPAHkJZ2U41wVAUWpfyNSsCitKaijQXLg1HYcgoieCWrcx13IGTgyVWbHxvUjtzSSWtz3
LBWDceHlIxQ2g8h7y/J7e5BTSKdS30Fn+2QF7Hu5s2c1W1bw+jSVm4qLOKtmE+78Fv2LAPE9Opgi
8+65Vt17XCKuWP7jOAozhbhAx8EMkckCHy2If19Aq7B2nzSpPOcPNpsOwuwUZkumU5mV3MXMLgGg
pY0PDGvSKuh8In28KWtfNLRteHosvZpor27JGOt+NwN8hwezTpua9Q3K7aFOlc4jainKSOq37/Hb
K8XIKv9Wqq5omLj0D6UJKV6K7qQTjqBewh5TCs8zNuc8ZhAHu1GAbD7bwNji0/SeW8WgqblcghZL
++iJSrBnDkXx4lZwc7MudfwAuFpcsrLOS1tDk6wrsDpmN39cZq/mBTPc4jW5sD57N+zO8c20aXyb
o7lhlbtNl/r9fKNmXzCRdhEe7viwLylvoxF6LjD2yxeJ0KGgnvF4uESlyVTArSWubjLk8o9NuoUn
e0NjVmxDRB+52N12YAxECZAYrZJil1bhXimPiMSXl/r5c8bg+EXxIMNnTZVxteglDzfhcPmmrgim
D3JkAF+jZpNxvnLHaZYEvXbF4cY+OwizBn2aMaTbVg0S24JIheTyVOXz+bu/QrPSLHAp3/bYz+3E
kaEFrOBxdsmf9vtMCUm5DbdSybIvKVri/ipDjNUd3dj2wAyLw7iUuZ+tm2m7uMVlxeDlOVJph4BD
Q4+NN/rBWFfJVcd4Cvpg75sHRQBC5vlBCEIQT82uEghkfypZ0/z8G6SPlBj4mfx47eOCL04ER9pl
yUoed3m6qqCvmRbj8EOZperK7Z9ZI2mMNCYytPqXin0j/Jxou7tWcT/lg7D1Ijj3FkJohII7JTom
XdD5pw2M6HZgTDCZbSimK/PnpTKvfgJNZvpCDGdxWYwYjRlA3+rBy0zNefO8sMNMHrw7v4LVxLJF
pCWTf7X+pCk/KlujvEdAOocCUFvtDd5iJXrrRawJDF+nB3gRZ5GDEuqwbpYnpWBIe3rqDjoyC2S6
JQUNT7zsvm521vZCuhJMvk/Lff3xrsM+FkrFTDvZeCmt9lpIMRDvMpJWPMJVi1ljxYgJPjIbYda1
Bz2ggj5/QW64f6qK0noUzKuSX3bPFLobRybnUTkepDcZ4Y0l6Or951i0U41Mfjc6Ug9SugqWDp7D
HgJMl9WIpkvi8VU08EcQ4ASLA2OewB3DcC0xFukjbvT4SAaj3MInmAfWDmD3Gtiuv8J0sIr8CMU7
xMm60P7+HwHHObVZs7mcx4F1NLweYGAn7eAH9xwtqOOCQGmJvFesA9SyCXwoB+TaP2iv7q/Y89uB
roL+V0UueSBVItqHu+wLpIlTYGgQcevNz+NBWkBxp78qWNjUNJK3Q3r+s6uU4JD0tOfu7NvSsvYv
HG+XnzsCwWEhvyYQuzokeR35o+mW1r3l+oQOGI5dZYpfPHhr7pvFbP9/YUf4rY7u/Rs6QXOiAo3w
/VHrOIUJrkg2bFtpLfTYUhGM7IWSVWmIwfPklaN0xTSaG1UHPPsivoTNq/2y0rzvALdSXIFeiUyV
P1mJAvax2H9xhODfmOfADDbgyuIguQ8Muyl7gsJAEOJn3iTSFBLm/peXgj4/k9AZ9ahegaeN/x7S
3nOmLKCvZjxTYz8/9qBj1xYEpPKCUHx4JsigJ37YSf7XS0f+sHOfPgpPxsVaNq4X2TmpaJFJh9mY
bSSP1GVqhjtlMoK7hEc2Nh9II6n9npPraCUBs3g2CvryQl5xNkzBc9W7K1WPS45tYssj4ThiQyfs
z3weoCfYLGqwocsV79HIUXka0Og106F+9IkdlzwSQdh6Xbq3YTgFTbQIF/nSiiDMA3U3djJWbq9b
I0A7vfX/5RRXs6IHQ4WvaGtqnH2Exr9lzK56WxpeQ8rczznlGY1vyBPB3ZZ2KbRW/mDCsMd/G6cV
9y7G71EdoNuojPYGDmitw5EOZDBa1WyOdV2WV0GSkeCWoDFbqbEFTKpxABaUeAagawHY4sb6a23e
MZCXq4Yv5kZ5IlTemaclTQKrzC7MQvU3CgwWp4gZshilx3wKvqH7exf/1C8wGF1/f7uS08Oi6Vzr
WWAQbtdvhRtW+ZifsF+PahfGmP5IxT6UppjbbdEBDbiTLD6NfQFgmzHxYN2pxeEMsr2qJwrzWua6
06Q/cDHi8zjXHtCCHFZSW3ALnB33qNiBCHlyQWh9GES5mJzh9+QIf+2JMXn1cD9eNklmIPgDatQU
ARBqJPTBRfvWMfdBCm4/Qlp4ifyScUa9cFTziGAHN9f/Tk3jWX1u+ISUo8CQSprlP7gkTmtSeDyR
i2kbAaes87bY585aVQ4kaPoMzm7pp/h6muQW0MkXIV4Qbq2Aps/KMgswlERlBrdR8iQ6t035CgGv
O8FxU2IcYJ4NUdeqBUwAXm4cfhpJtynwBOz0tDPsW6hxL6j8b4uUMnSpLju0/jAiW1710qMBMCMP
EKq8zd3E0fxGxjQIOJTz5hBDaFpjRN+tA1VmOpIxZSYx9MjBjuM7JMebRPdn5uoocsRPz5aiT9Yc
hfVPDdR3pkgULBhpFNu2/W1ExpQusx6OOCcn0DpkQA5EdBpkiUXYUnH3s4ela+KZg/5cDDDmM/r1
KcGRl0SoE8MvES7Il8alvPs/DpvXgkIcz7W1TmpZ6Esb9gvo94uI/ENTJRXs9ogKuBcHC+3eLe6+
ABpHF3tKVWspdV/tq5oH2ccqpvvQHX5chmJuXtP/Ibn21bX8QpGlQskMLVIfD/N6zgflSHv27QJE
LfqsI4vUuNYbgrCVqet+Fxn2rwykbZGqBKoGwOTpE/U70C6Eu0llbVn+7xOWu9JkreugxaHa90d7
n63wbBue6W60B3qn/PmKsHurZoe9z0RYcoRdKB589eR1iLqBK0ym//LsVY8ZM57JSc9EjKAMjKgI
O5BzfWDcz9TJoxOop/t5av4fRzGnOxX+Ca3ORe/07dTYiRmBW2ULXJel96e8iC41Ovfhodm6/wpY
13HNEyZZhwXthjalm+dbUKdQfmkAI3J29j5jOeirsvrYVl7f/JQ2zlI/RjfDjJQdtz1EI3hKAA5d
SIkWZZt7LQLsrl/XQ5A5BAVyl69/GuxYpyVljS9Ga8XFNS9UhEvhngKPmKw/cBrqa9g2C0j6YnGb
tkqqU/rpjpgLLgnCoquvArw+EHpAaY75bGNvWqZ5E1bGFuzvnf+XCQS8zMLzqZPjYYx3gsIKH9xW
xUKKQLOqVULGcXS8KS35z5MJJbC+NLjLHh/lA+KNRsau1tZ10gmIpyVeh01z41RG3ZD9vZSZ4QGX
N4nF/FWnvyrRW1fC8FnMud0nkT14mtLeJ/qZYL9Huvzjr8ZXTfrUXsCuxNm4pIMttUfJOTkvS8sr
xKj8aYGQNTr27RrAsCo4Pq7ZZNA5R7SRm2fUrMI5mUg4nP3Ud4kP+U8MsfrKlooeuCbJgTzLcNPL
X51I949ptQjNii/e23xBhhAN0q2l4oMoZAdzK7MEd9jnqzOyYA1ymkkLnKrFjMuXdzihFbJ6hKDb
jEKkCIqdtr2FXQQyIX5SZ3pQjURcACL8Sr6m1hk2/MOsHSWOkNp+S8RTJu+b0L9NWG93eMT+ezNa
KsPx2OGm8o8b2xAEEfqZO6nleMiLnrAHEj6kmyax1UPHyF9JOJQV8IiBsEXw3P5K7gr/0+1JAmtr
m2fkCOSgZGiz40hVm+nEcs6T1yzPUCDhbRC3170Rpqrtm1quK3IzkkPiD6xybva3du9mBWMOHjF7
RIWP5MO6+yDcNhsrShnjjBRyyd8ndKNKhoJ0muLHzIIO55ysOI39geUL63bOZIAOA2rYI9RROhkt
OgfddiWZ9x+qIIxO6xMNHoW6SGLMf54PMm6bH34MHgup0KmOg30Htt+AdfcaD/80c0kvql/xya75
9Q7fQnQsH9xvczNYel+pMEUYXzbdH0WdRJsbLNMCSkIN4cUZePFDHvATjrqKYfYFyKEDF4/r/YkX
ZIndakXkBZ8E9U1eH+tKyEtCh60ikDKY/Kw1p4Lnz6/fxMnk1TeeAdKYp6OLnwxLay6CDtyjxWpX
eKvLExH+fKcRw4ZOUpTBLjkB28v1JFlqv04y5PC3ROqM2TUbdeTkLbf3Oc755UnOYnY6M4QApEsL
LL0meY8kn0bwMkfw9AnKweS3mEquoU0kqDAk4kbRJwDDgz1n2gNxR1lSXV2cKE6P+2QZGafzV5uL
ollDMTtYBDLBkyKis7OOurr940dsW7qipP/kEnyQJsAplzm3FsobtctKODD4SmtDUWSN/RrbTaZV
v5QrHnYsjpO9MpSSh3j77jGcev50yEAX/t3N56CLYFmNrEHRlscODLCxBFp3jeWg6CZAW7t24cJ2
FGgGUWI6rpgtPheAIyExx/nN0h8Q1JIfQWOr9fIZhu/QlHgMN3SImVxhFZNPiR23cJdhUH8EEpzN
5y+g58hdEZKT0n6GGcITjZqLAKdbM+Pg9iZVuKlk27wqg4S68CerIsl70Kra4j9sq3K3BAivQj44
6v2WL9elWRgDFPuQ15WX7ImVEE7wFgCU750P9ibKFVvymrEoEwv660nvoKWG0/teau4odHvjrieM
fvVK8FrL5Whp28IaI0R2AJOadKq0B3DwsYL08b5UI+ttqY2sSu/+KKSAJFw0NteZ2mWTZvYY6byl
w1I4Isg55ByhdYAG+cM0ctC8XCOXgYq5Q8yEqAOKOCsVYNH4Ro5jEPovpjZ0gdhiI6lpzOp1ecsP
DbB9S3Xxo9MgfLoc4NqIUPYLwQdQQ8HDM7b2Bvk2O9SCHfvp+6AfVKJEsj6ah9S4LW+oSAaxhdN4
QISjQT2ExPmH8vwdBw9hIwspANmO/h4cNaKhqv51gYLv7Z4bSp1lzjuuM+pVzY3fZcigTUXROBAv
E355HOV17DQgjI9geB2Nxlc8KXPK78VEm5dUaCo78fLmFNs0gkYXEHtdtlV1liC332FFmEz/fHz+
juRXlhuGCGVceZ3K+fUuHeE/B27NUJ0qX+OlujkXR0k+OtUOP7jLuyH53z8CerYZlP4YDKomIEEo
XJKtzp0WquFml325X8RNqX7Cjo2ddxk91xBzuJBoK/x3OCLX17wEF17nLXvOLDuJeDTcE9AHCf+i
r03O8zOOT5IzYvLZJTWjjDuYVOJ5jhDyLLHcjZUo2iTLuOq52qAQ+338yV3fdWytgNfLQjUVOg9n
/ya6awNPmwP16k9Be76Vy8sOlaItQsEq+dRCSnlaTXzkdT5f+YCov45immtx7AWnHvf1FfQJSTBf
fKX+tMTW+g5QqXOygkh+5qKhkV4Zv+J4CgGFpKKSBf2tdkBV/vFv1lVnYtP1N0SmC5s6oHeDs21Q
UMS6MF0/UOyEqv+L22DLNtXCsIU8I8YLo6fYux/2bwUq7V3cFSzlEWUYVytxIcJU2qYNV8kDvlFo
ssBdvF33dqiZp3Eaf52BEUn6FCIGOacy3itbCmqC3eeRsbqek9Joum0HCvctvU66rKlqg3aN8dVz
e7oL533F49UqLy8aksrZTVLtIu/WAikWkibULVvfIlM+Ptygvzv4r+bSE1LmhNj86TAM7wEaL1mh
ktLAd1Ttls2Ec1ai/wr5SI9iHvT9+5mG7yhv02hE5MGgdnWF2luJsse5AkpHAbHq1YaISEOQhwpV
uNAZi+6q/iRl4/7YugecGMWxRl3lbhuNdksGvxWhJasb5jpaaqeNTmdSZiVnSD4nbcF4eer9b6LQ
GdUkkP8wUmH8jp+OppAnvPqp56YPnDqJTbLktsUzKEInc+qqoe+XhbJvW19EiEICv6+gCCZTljaw
gFC3ZE8ASiGNcehuV/egrOCkRGAZ1/tJIUzOd64QES0haknbbvCswppiuBOZG1mPrkBlpm93TO7o
5esYB7f4qUqSniwIaSttWYK7TpXqxn7TbYGxge2HWVVRPQ+QpWFuEbwKvT6So8nogJgQu2jecvTJ
coWYBsCvbEpyixu0AXtTfguCi+/GineMZn56kNMtm6R446t/vMSuxtmI1pzizjP4IOxGUCocbqgg
/vxQVnb070gjhok9PFO/2hH7jhKu90kxVldw4hBoy9jeT5YshUaBFfm/z2OtGEnYZeTqgVp3RvQM
8Yy8vxCJCnvn9PKTMDTgUvms3zXkP7rJXqzR70qifk85P5qTdYld2296sbu6Un4S0QKO0f8pZ9Wq
J/LS3YnPI6/y/5rtPn+scttGzA9aztue1sbl+1z2nMyaZ7C7PcXG9lOBz9U94qID68gehSI6xrgi
YfONTIePbCl3ooCxFgR+AO6+Uu6hpTUxLKITfYCgQOYJd2dR+HaY6FMeJ6uWgOG0SXHOBVWiSWhw
xnJnBVZ6IV4e/khjvDQuTV26q/eLbxSu7Ii2EAXCuSdGZWcfkjIAPYfQA10rK2LeVrI6WX158PLq
P17Cb/E9pfiKMBm9DBGBIrXIKnA/6xC+BmWwCtDUuXj3zyCfWnE01NUhPS93wJ9NUri6kum8y9/T
qMehgzX7wuIkrfHHcCHcs8+McOoeiCP85mvljgaSETLFyNBWpjqlIxXOfdQH2b/o+zdzLDpTMdAi
wgw4JWYjvtVWuy241XpGMKly1OzbknZ8FpyEHXkTrFxrgQccD0mTWKSSgLWGurela1nWPhcdjqXp
bAg8DaE1DJRgs8f2uVst2LQHmpEM0ASRcuqPPmy6or0Q24PScNHHUG7QTKehvtaHNgT4t65yFuWr
fNFa1DpHgMvXEasAuC5nDxvt7pWrmZx9vNx4I8iF9D4sFyTgkf32JaVtpDsKr7jnkEswxVtubuus
xsNz23VUh51HcsOyPEC7za42pFCjmWxJb75ON5dFg82ckJNpOzx0qdJQ6fillS0MBs3octoNsNx+
7ouXdhClXOlyuxHFo4pE8sYMwryPPR5PoQ4NpmH76Qs7VfnbxUAJyaRlmj3GSiC2pLWb/NNvz0Cs
OFOyEE2l9chjhKUcBlAUyO4uVl37A5i+VbYgPjZxdCPqSBg4sk8gcw5puemhOCdreliU4df+V1WC
YB5iLSfqjuG2G4SIYrbbIsiZE/rblbsmBRVo07q/9MO4X67jQzC5HYHqDehk5zs/+chUuInvVEi1
HOfi8Z8uWra5BE43wHdeyDc08RGfAmKdMkdX1pTQ/JPXrJT7EVuySqPzqX/LOC9zTp6zpzYfj2/1
40Ni6U5lHOlwttnow3CI/dWaV5Pm54lMiy6qmL/iTtRoKB+2USRbX2m6YEIvw7qmKd0DlU83UqE6
xBy/YpQrYjMGjMUDFl0O8iF2M/EcHLz6VsbM3Kwexdo6kTDaqGpovChkUWqzKd1/Vr1sFJk+pLZ1
OXDjK+4YwcLa4Tc0BCtpqNL5YBp1/CGqCcjfmQfgiIuZ2bK1rCp7fGNa+wQN1IQ++ROecvf1oeO2
a3f/Lg6k/lGoReoiM73qyfMxLqQDWr7UwOOaM0fSor0+iwJdsOfKF5059eNy+ZmFjoDbT8V1QAf3
xz44aWsgksQBjph1C6zM4xA+60eUWIads/laLrbecmuhoc8Se0QU+nU+wCU1vIYogSw+e8EC2Kc0
TOF9cQ7K59ivYmIo31ljIUkdhAHj69s6n8MO+GrlmzHASJM3h4852fbaZBCx+Z8auPi/KBleFuVY
54TCSKbaL6P+tZG2zYfZgvvBZntF8mTXNMK29QoBJ2WVOdSuyUClR21y68bvrzGD7mVjewr+PRCo
SKoZocApgLW/Gu8g8aQ/NXps7QbKUkPhA1z7fqPrJM0kGE5lxwywmAventxc5pV8BXnhYcmcGqcy
2dJuceJOS0l5DPnDfk8yg4m5s04gmJWY5tbo2rTLkAaJwvcVP+fFcNSSSmypp9REH+f/zPWgF/lV
XUetAxNRqvluPIWvBleZE1azkASHy30ufdVvUdxwgCRaNYz1B3wzAE3k1tepIKQRSJ3GWppZ842U
bxuvrHODItbqybw+WajswaBszfn7M9hp15XAlivVkehU5qxOG5TwBHmfaPdPtKFHWk3JYLRuI+6T
AvqT/iWmcVUzWGo7z9TJ+JyFrMb6tpvlCqjHsgHnBOfYutU2k19dax6t24tbOQzZF2MsyD8tv1a2
MARxu6Who0x4yYUp568AtrzoVldG6RwWoGZGinGS7UQzkakCxxmh3Hwipru7i8PNqQmjr2kCe0o7
1kkiQcuv+vG5x8yJMs18ye2ijDCt7YnKORoZiEGYoZISECl5y6pI0rIH6Al4S2RzyK8Jlf8399EW
LGmSXmWnljM6tD7pHZRxKCJGqL8dUCZXX4twcRdpupNyqqmgnySnhUOsiwM74e8JP9m5JbDVz3BD
N2INZCzU6B/hy1pP7PpHhNEg97a7iODPABiHXaCtjiD6M2AX6/B/gvaVgnuo4YlFrrQ86lii/Z2T
dbkmdo4wV+oSRjep1byEKT/cnlqlk0od14WLjKr4GDzoM5jgJaiDK7t0cCyrUQgjW1W+mQUII9O5
dOwARPkZLiaz7iEomIybV4evvYHB7XkLcHZWF3AAMcSDDSdmLmevaP0V+KG5IiEj6KuIb0vZ5Moy
7gBow8wyOmxLrKz2tZdkhC9jHg1uMGSi3Maj00AV2bzI82+bBYzk2+U7yJgkWEuAMJSPFX+HMM95
YvrRyj2l8RUBzSpsXxl44jfB4tt1K4hU+W5YRmwSCcY/XKz9P6t3lmDJH3qxGngTHt/t5BSZ3wWJ
O2L/LGXlJP/Px1vtwqog/n5bO9wv4Q3+SxPyE02Y+Mdd6Hq9TEX8T+XxIvMIsWcC+6YNwGkeRSle
vNncXIvltvFFhmhOc1znJJYWptkAl8O6pmHT5XLi2vocsucmXzSRgJirV2lE41UqBoxXnEipFoXR
TTbXA/to2075G73TwhzcTMHU2oOhD3orllfoCJhWS9vfpYRPoL9SpegKHhof9VrPKBX43Nns15/k
QLMNyk2LnNtSnu8PB+jKPSjwcUqEBTkbGOBktmnuMXWMo+1hUKSA0WFY9GWRLkOF3+k42QPQ7N4J
skC2uN7tVUMfeaaKyTIzNsGiNlrwk+0lLNZvZTPq5TEYnCqMIUCZRx1mBOiW6OBTsA+CgOovEYoO
vLIkydLsrh00QeGm4y6DRuJk1CbeIsMx+iOsdDEHMYX3oyx5tDXNxacu4tXcwIA4a9jAPdnKPNO6
SnwFRtRNblFyU9/U73aQHzXaReP4AlK7o+Tp0X0CE1+AgVSdquWRNJub97XkH7EgsNElkKAHszXT
n+pyjfii4V4TuYiJhglS90c3C1QxczktI8f9t3NU54x782CRo0CTcJxUsl+cnyq6rev39JRQDCEX
iSfKOrFUJWP0nW2X+cdtTEFaG2G6s145uEgwLtpTwIXQNgwZRc6p9c3h32/AnphtCP7gRCHx5B8e
xpmuJ3QVSVh6SMxFCoAEQ7XSGWbxD2VIBXq3jaKRmcnarRmzMDxkcclwVDJCK5XtTyqRqSXsyo3M
xHTOOSe3kTUw1rg7T7nZDkJ544ChFC0YEQEJlHgNIiNqTd3/VpHOcgOJDcpW9xiLEp9fanUgOmxx
hOcQmCHDjHnxAjcX65g6y5WPHLCRXDuNCX95/ZV1+oWetliB1o9WPAsQt6CyaTNJ8IEEhFrMRE4q
lFjpwkqtyyLiX4wlJoUPlMrpxKtRSrB+2bS5aXfJZk+qWUJrDGyZ/uPzueMvZO7hfiCAmo8+p7G5
Cjl1+ucdP4jd+x2O9i4HIRFztZILo41olL0qxWZkPl6lcDJBjSvZDv7/OAqIXNo4uxNA9zKDfXkx
Dl74JvMnh4CftdAa8THNDt1TlGtz97Sy/WmwY2DPS3jYtGWa57sceVodJApp6swHOIaeMioTDlTG
ruJXw1+cu65mKbbenhiPTdUUx1fM0dhE+EL/mmivNrEfub2HuBokZcbaSVR0mEgdRxmNEwJX5GgL
BF/SCJyTf7ln2SmzQ2boSQAsgxNsfhm0lyCT+xeaD++obilPY5Jqzj7Z93zHEomJjrdeQy5iJ9MU
WyynAbGMxVOKHk3VGcn+hrUVgrDbteHujHSdOvZFcFg820Uh/tt6jx5cR/4/ME2U8dFupOkkSShl
Rh8rY5Vjxv/v606ItJpnB4Ye3QL3dULtJWENKu62l1r75mWZhJDWRyz61ae5T9rMxccOvC4WZB6g
rBBySDcaXjpMGhlyvowlxk7bQrndOH37g1ELS+esTQTWndTNOoA1bZ/uGcWrJbbMyKScCfMKkxNB
AiXkU44M4NNLKiCZcdbAstXPQjdcsTmDBvIEzcVvBDvp2q6Vg8uAgFeu5zGXFnWUaUZequ/i5++N
wd3mLCm6aLaVWBoG7Aw+e4VgYXezYTvCVF1ZqraKSAS+hEuYVtkYUxpKSec1HNbIN5LNsdvD9Lgd
NFv1SSFOIjcwli+uRp78kgbdNne/F3jbl0yUg6/yPXdEPGjQ2SVXRX56Wjn7FqX2mdyfac5I/dqY
+VUNE82JMhvsRPsKVHlnXI1al8ImdKqknALZ+NksExQ5xnAo0VHgLlG9QwvJYFpbvWGAgqOMPFVP
QDB8uKT1IlFwzunWMD9Br8xFLWpK4rHFhH4WEgDTedzDzAGBqoJhcaPh58WzWJNDcGno8yUOYlh+
GoyxMo4lTfy3dx6tuSqdtJ73FvlHDjNlZ95zy1p3RY+8Z8wwzBZbRytAy2Fcji4rj8MOw2Jca3nn
nS/WqLbF7ITwDsc681UOkWT91/xbi4FGNeYiKZdIrN0Rum6CX9To1jp2LcbheQS6ut4g+EAm84pI
mTqmETV3H90b27XKNdRg2yZCNV1+IHpul2pD20NqT1GxvHgMJ3jCUkTzKQJY3SL9U92uNR/DloKW
MLwXsEq0VmkompSNCu1B7se71dLAqV4ztDBsRVmP3jTElViDoY3XZtx0rddNVwXXJpZ/BdrEryRK
5pLKJSiLP6DOdKhoKzC8ZNcQizu0nq5WneOV3UFYTf4he/Z7Vo0gMJbXBKr7NmxdSYCTxBphrtub
cAhSAa1G1SWqh/WJNraSCaQuiz0rFuqPTwtVEC48C0bgq2Zh/95bVu1RRJphzwFfg8jJJoQcfcUk
ed4osHAQ1lwtoyas2rhOXIdTIkYQry6x54SU50we9V8KlTkkdvYOj4qaWp34HSic80nl+W32N2tM
UUPus+CnPGNKywl6flTkkhOI6nm63Q8uLfsJIv89uCbFOwZqkrpbI8IEE/Md5u1IJemfd7Th3T24
49qouFGJC53Z/S4yc3js7A2wXi6l3W9eQHkH9oJqhMVEmpI0wFtLY/rAKPnSVDF6xSvjR7qj56vf
FRuqvqck+y23OW6/kCkEj2/oO4I/yN5ZZt0viyQEBqlUS19+GBI3sjJCtHDpS95gDIl9f/AaKylK
Twi+M0jwvnCllTQYGt+d8vUD+wWittVDx/jovl9l25XyfREsz3B9TM8+U4Ui4gk4EdsKNuMMk8kc
2CS3Z7Q1Y7zNLvVHNp8I7PUcFuegMRImsZlm6QYxKi74yCq3hEi2ehuDGDa6NVkjKt/M/sV/fzb5
qDjBx9oyGCoe556Kn7/ZNUs7eaMTOaPV9JbisDlS7owUBv516GNIHIullEs4eXa0FeCNEJ3qq2On
KtQfQU5MSPyhpCtNmKwjCNo1DRlIeEvWZHMMy3xcdp8ZIbQTAGxigiJPvZTrR2spL+FX3u79voFO
qqIAjSbSKh+jRaSMqd7bFMHBOBtWET5XPwv8CRRRI8JL/yplQfzOyLwHdd7f1urBkHGOtXQaUP4g
10WkogTYp6UbVKMXBYA/+WVI7syyVtDBpfv5XTPO6gVHZWJPNi0p34xe2NEk2qFTJDVJGX25h2zY
x0y1eSZ2UD7vi4kgxzqaQLXcKpsWDBloOb467cvTi+fDonT2D87+Nd/vEJjqjKE+IjJz632gbjTh
0QGZKUSSmDRvOvr2TBpqjWRBrJhZ87O6ZKcFp8Myv032TZ3cr2oSegRgaWWM/ew1uuhLFMVXUzbl
yCPFFLUzmQF9pax1tSq1TN9Z7/DaBWbhvMp9T4W7EW6nsIUJF08jx0L6eXKTiePwkmoXBCdmg6wR
dLZP5HvRTm8D34cTF/d3IlLRE7uOnCN32YsQ5SQMB19p7s2slhFrck6/8/nj0SFKdxflEIzWXZwk
RRK8bc2akktTHPKglYYCc9mvmMtV9gGZwGuuBs7GxUZ6xIx5AVrgVmFVAIcR+Lt3858efPW7eppo
YvGnLhlju0hILxb/e3+FFePE6pTScu9cr2ADS7M+K+vhrURgWzEL9VJFKxu0mNwMuSVRgzOaDaJA
itCbu2Cbk1f7U7FfGQPoxVFGQkUWoac/gDJnq6PcZoBdl3Z6kwUC+AmLqwBQMd5daHVyeQRCLbRm
l4U9alnkEFZ7fCOM/0fJnmlmOqtowl3I25ZSVGRI8YhIfu7tuIUPADXAumgSzkXamGnZZxEO4RIo
6/tSt0nngL/viylZnFERIm9Q4wV7i9pfGzaADKr31xvIKCmMKJpk4hQ8wS/skUD9ObhZ7nOJ+AYp
aQE6bqFOKHLhUXvPYhKLMBGqE6iHyqdfZ6RMaQurd8Stmr2+F4t+TL/0n3vyr9/2zKE5hdtLy5OT
vBFkeSPVnb328O6feUQSlIHbAsiTCk1Ew22TyHQpz3ja7L5ByjvOAOM3f/v6x3PtW4VYzPFIKyrY
d3mwBPXmGD2rlt+hKqQVJUfMhuzfddZkqogQjrzpC94ORHsT/17iskZbb6mQgxINdUiSUtleEdit
/Di/V1Chvr9RzGYCQw0IyTNEekhjHsIEeo83aPmsl4WF9fzP5RmBbG1+0prPW+nMF8jiWGG0y1y9
jE3Qj6UXkEBl2IeSv2PVsgak3ZRwkXjMso1kDW9XnFAVmrjdR+qddnk0D+YVzRrfcGSMp38Y50xz
PV7cqPuB8Uvp254el/itC1OCn+i2qE8iDFSHYO7hLxOUbM+e25KQZDUNdzfqLThy6Z6w5CHYHa+b
H359Ksf8RZUyVpjLuPjrgEdTnlTXiVoEiNedewRKZKvB/YxxvaiWeQ9+T8LxraSMZdNbLp2bruU3
7X8YvyI7EMaeATxdqfaYLUu+ELYkBgYkxDKaEtJ9o7UKXVL+TeQja9/esIYvg++bwezgrlIzCYC0
EcCJkwbM9DOPQz5MOpW//ZfHRVpRJb+oLR01IV1RxGQ9GkMG9TDvsrOhcR2ZBAIkg4qG84YJ8a38
MRnzMCCW4tguBOndFkheSBvIzaL3YGSNoT5jkz+Fhs3MA//nfcfs6bNxF+j48s27kxUjKvbiTMJJ
dREiZFORTpZaf+sCATn9Q6QmrQzyVv+Qn5aN/0+j/lb9Etgssw4EiE2c3UM0b3i9ZarpfEPGMNpJ
e67KLSvgqbiQ4o8tNmgeGdv6XqFNCHbeqwkP2B+KTWfeDuqUpU8RLk+2Y47HxkSG8IgFrlxf1GWq
ndooohXllIUWKFnOW4sHN3CP95lBZVv6+WMC4lBCiITBmPQcBlU9Qyj40k4B2JKDaM721l6Fp8CK
eGBzruwDXKL0M8BnRS62bvdwj5rVHbbCfixt8dG3I0vA+6bg+Il8/9CIta7ev8z51WDx+iHjQNa4
0SFFkYmFY/WPA/ScwFoqoMTAW1f70NXt6JYcslYv52Teik0hmYEltbFEVF3ryfuWudeO6Cyy2ScS
uJDuR8mBZZCeU5nDr9zyuKwTnS+4BI2XgDL52jvYqj58X6vmkujF3GdHrbsFBHSLBsog1vjOdEwO
PMs+pyHE/GTeGsOk52w7vZfOZTIq54YFYrDQ1piOM5QjSNbJ+kUplSvM1vztwSjwk/Yo3dRsBcRV
Qesg+AvqvoLxgbqJTTLyg0qJOQ9ZqXQn2R7XsZHZQj7ZdGWjt74132GkllO1nho2ch9U9Qo8pO8/
v6ZIO8IpGLcStNOnzC0mxDbvy5llI1qyLkdvItQChP6hMA5znih7gqPeurFi3C0UraCZGvUu0FKq
gF4K7wHIeJPNTOcwcLGvC5UXS6Fn3BaRBqtlByuX628uiV/nSq2tktoOo4F7dbdm3CmUPxqSkBpk
KHN8VYGY8DavmGsPGOcUQKIWz52De+4dqlQyzhcl5Ddvi+Y54Nq+jockzgYm8kvv3FgdbqUyq2K2
3znKs/BLksL1cyn2HGmZINn8JlJ5RpJ4U+KLnF9SgUx4SWnqINsygMjbHz7jYj1jVyU4MvsiMlKv
rFt94tYKtR6cDMjcBLPEq+IoVDWiTv/lSuExv8qGynfooXFdZFiR7fRiJWeJ+N97WCDCa5cGD1di
QX5ua2XMcSrNrRecAeEJqCqjXrtdRo+OnwrcDNJzY2ZwYBSUBZVQhoMh3czimJcY21HaDzkr4aYc
LWzaMWehiAMpUyL5osf1LVQwSpAVskKLLZH1xQ6FQl5c4KPI3O0IS7C6lAB8cdONAnV++5BNO4cI
09wpXdS3hZncpPQEYjkkWxfdLqc83qzb+EMpt4FFuddVLiT+f5AA1nGPe5BDtscuF3VFa+k/tyrF
95qD9tmY/YflTS2hzuRCioabWPShTBLJ646sOMkd9nB7Dp7es0vVAWD1vi1gA14PY8KkvD4+sshj
e8g7fg7Pe5cGh906CDVPfxt0mgWm4nnkqJBH4qKvHCzbpY2pqJnMTa8o84gEH5SQkQueHVoJYgXq
B85KUZ9OWWCJX7ZegAucEHdQzPNUKUuAw7IwEymoTHvCXbLzzL23hs5NeSMIo0vTubmQbJkRZQdT
/riYtrvcuCZXHF4dafJpBBVNe8yym+smLPTQo5fKppPn8m8v/wvkpzFN7qwvG8DOB34bCbFYtsgw
l+BIYe8jEu6lm3iAH6GrJ6cl2vopeZWDj2AYlQA0Yh3gNTSd0RwmxKNuAmGuEF3g++Jj6ODRRx5K
4Z+019O0ATZL4YMaaEo8C9FYTc/4VxHrx7xWm4U8H+UxKW1ovX0yohlMqObfmaS9/U+G7FdOG5Uc
C1gTG9xWDlgglKgapk/Ng0se/qEnx6TduEpeSerQOjRM6RpUGhNkSpEFp0HDu4Lt4bUN5ryicbvY
1Kp4nIFEhQNaHyC4F5hr9GHSzYFDLOaVBGVS1sSD6NNSA3+UKEopMoTvQp0Sftk3wIKde3n6Vauq
1JWEwkDOKi8ReW6hR2LqyNuWls7KGj7td/tJBLXAFk9F1XBnpgkWlwnJn0HbrtZtzzJfrdLQCE2J
V1/YExU05ud898jppyXbvpAGxBhQ9cbycwBomtRsDLEmCHmAiQCvcC8IJlbWndYrbiEVuuxb1LUX
BZdaqnhkol/Gyn8ANLVmTkAruYj8sJhhZBiO4WfvbxMc3DxySF5Wboemj2Gq2ETt+ErvYloJIhKm
6q0XbBk3rTn06UM7qz7yd3JPSCszuOYRr4Y7jA8YPFijzfF58rzbqgDCVEpp4uhN3qpBZqHQ7V5l
GIgGeYbry1VvhHGLuarXbHlyflDK8JCv2ZhUa25oIeBQLK0jcBsjIqys0ITsMl893doL4/301Gih
nGo0DUXuawJx7ZbY3l1NM1+1dOpuWar8A4AoWajT7EHdnF17EJIKkSa73yqSIIxzYgHs1PIYoEEp
SImxBvU3TN3dNbPrPe7tF7dWrsWSPaNTSFRJPCbUJf5ISRcGoj4LFL8rTm+wOncBct2tqOhpJXrG
lIDanTbGu5l0vC2DYelif5O6LC96A1UuIhiBv4I2AE4ADJ5uPTAelH/VMUFjwIwi4pUuPqgo6aRj
2ICC9Za8bTH77bO0aAOCbEN3GPsCYF8XcEsenSLqVHb6OKLzNgarFTu21NkRjTPD1okU+kMe/4dT
vNQ3MJyLIVctY2Rh8xgbYd69SjpvfAFe3etvrOMJLP/zBpQ9fOUPqCPZ5l0iKp4fidif39V1ROTh
aqo5VDRAd7T0g9MhMT0e3ooa8lgh12f1zvdFtWu36liCIZV2gNpmIM+/LlxBrEAz6NF/HnkKQFxA
sUJ4kMP6W/3Pp8lQhIiWOUlcj9z/4Sf9UDSyJP+TX/gn827I13rEJ1ECO6g/Ic/Vn9mDRIHQFy78
m/aFn95FLrrxpAjYP5hKOskE4YVQdMTG3BvyS2Hr6zYrZ/+Aq8F+NAk4FPX0FXJzQv96YwIaucN0
vaDfVBD7zyyrq5MX8nuxGGOxqPHV+9Ym+4Sz+bUibxrZ2iuhwIccFBWN//R83Jeb1ztt3t0PtHGL
ajrFSChTfsTF7+Xhy652F4tptfEKKfgAGi3RuYO4rW92gQY0Q0IfW9zD0Fn29k7rSAybW2bjfK89
z73ML5MW8e2vKWYWMxF1301fh1oalu4U0yBR+HGGVHkv5HcdXT5f2PojZS49NXITED4GeUW6h4TM
uCdFGrDUomwz0U9H4IYzZf++OlQoy95IP6cAliSJVDpaP+iY7EjgNEz59NhizdCn2XGJyAlC7igE
r8MwDCB3SEvy2GmVovgSgzn2502YiXtCeiAAPNnQFyCpHc0EjhEpjdZQ5kt7vL0mHt55NocrGC71
NJ5HJVc7JOsd8YSvgKfZ3qGMcyrYiHPQdDa2fGLV0nXP9Piw/4fijQhJMCpyJa3BuZhbAby4V97V
BHPEWyJ++3/Fi9KH63pzKxUf0KQ5ht1NBQ5nwsdYK1F/FandBErJx1kjFw3v9lhbeYA2jepdvbl7
xP7lciqEJTUl5dUWfVVY5cXbOaoUqVtW3SIPs99zkQjfB0xSkhz8+VjnstriTon5wQMbuDRRcr6i
Q0UwFNzicmsvz0ml/+qJro4sVCUiMS6s2eZ+2zuHaQ8MJGyvuxmrTvg5DS4U49ZghaLij8zMC9Cb
sajVRyIheKdU6z58oXDNy2nbsGAq0xz4Xqd8tuAVhhbM3oxonOWU33F5zXRnJ3eMk3giD+h2sDlu
22eahpfuiV5iXt7Ssr3ah8RWYfODqh3MXu8CVoUtrsyXBrZAwDocTHG2bfnAcX8Io95jIg59SmOn
ztSDfFTrE9C8CXf0wyj/w06kl/cHd/u9bk1nSzL6E4JCrnnWCpZonrD5TkG+D6l/2Q0AmhwxDU0f
3AWpNmrf4+nbK1l+BV66RduAKym6b1KoRIzcvwDHoEx3iRNi5btWCD0kQlwIYWclya+wzyjJJmj0
wwFqPCNLB8l8dmHXFY6B4OSUMZ10oplgSjJTNd7j0QI3PJv2K7j8eoFRUFC4qGLglRUv2RtAANZ3
Fb37EWjJbjMJodll7YvETL32liEUaUSRLIzFyIkDWmvqamipG+9trjfBPwjVLgsKR/rzmRIgkbZA
a3eh7gSIp0dyXAbtQLtJzO7aWN1kCPyfFmBcXSFZcmKZMJdZ7McQJw8bxmwWwU2TlhJnaf+KuIMd
qfU1XpAFNQorWu1YprPmQZiN+AIs/rwNF4UOuhhZSKn0Z6DVaSh78k56aGiX582dmZ55YkvGEP94
ow4cjYeEr0MoMTX7OEu2Tn6Kk55weqCT4YPrxDy2YEM/SZ+2AqKTBqdX0tNvMaBUAR1zyhdYKFkY
T2pVipAU2AXpNFb4XCIPjt61LT8ykl3l0QUtQbfdBQczSvm595W2kDYXhkfGmlLUbh+6W8fDY8kz
cgNsxA5W4jGEihYo7PqjrBuZP+vSYrdoUZmNIxjGmPQ3mWlx9brZop0pueUrrXexHm+UqUmYelTU
/+XhYLNXqwnaRi0PEbPTCIbOxVW2KkXCH0+zJsx2VFQKfLz55s4AdBF51WLEzr+/8tDA5Ni1Kfx0
zHMBoG2PO0SKpwada9PAfWhkaMbN0k9MzpXjHezagr+RuaTLS47sQ71ln4nPb5PTi+QKQxK9Xd3W
D2Ifd37aycj+Kazw9M5eY6gZMWBf5hjfdOuUL6Ju9gz6mBgHE52x92yFO5Dbf5jMZor4R53sWRAb
8cRRKXKzVKc+qchJ4bmP+SLtzrxYz4TDIxNIebhDtovM4Kf0oKzEXiUPT4lM4RVNEfG5qls7DV0t
wBHxCShZRpXAR0CG6E1u9IOKL1Queky4NuUW9UULf6E8vjsaNcZ810+F9wnx4Sex7NpMuewP1bZi
k7aVDWBGFpzqs0xjSPmcsimMjXkj2nUtPPeiiQCTGkPSAEiV4s+6WmIecwxmlWIzXduyE/0YSSyZ
DKNPmCKf7cnXKoV3GbnX9CGWxPIPwk+QuNTqv0CBhsyCFoRZySViJawQGd/4j5QWDDbXhv+Fcaog
ZOQ3LSk2woNzFoprijlHOPSA0F+dyNFi9xIgKiBhISGh+dWCLScQXv+s+d3Nm5gNZtKMgrJT2SwL
uexe+t/74cap2VCnS/abc1KUwZbjp62gOcd8DYGJBN2pzsrp1c9zxLQ/FLA1KMY/bunNy4Nq24Yv
ZkIDlGtNxEZw0SXO1gg6pcXkXk6fQX1Y70xdefYxiYmBeRU9D0BFbpGjIvf4bCB9/H69VHFQbUUf
FYezF1Npy/2/28mad/vBDURmmwVEPvgOEb0xgo0Pdt9dsPG7SBhr61XKvBqpevGx+4xRHfZUhl3M
mOK0I2GkYPpacXlvRbEjLi2Qh8x/naDg3K3O2FhsNZIWSslklzXDzB73jn3Ag8efKKLDSLl90gwg
h4wJ+2PnXw5vMHFGeOpqfQzfgAXrcfunwrfe2X9ZVa5Tjs4kT+R7JRYa1vZzioQUNbdxr07sPjup
SR/WoIsfPMB//3zPQEBb8vF3OE2ZLBayUz3LsXWnTh6YVABIFDIyBtebjK2M675EtVyEiJELmAsE
wYLHBATqTECr3cIfS4ri4QIIeSkI7kb7dF3AfMmUEf1vMa4dMZl2JRsNq21x0R2h4E82vo/EkddQ
dyYkjXNZHRrOPUNm1sIGghAaRn3QuKZeL4tVpVjqga+ZfSdvMz8qIoDNXB6CVcZ4TeP3IpFtGpCR
cOV+0I6pUg8QauJYQVzt/m7cyWQ0pxoA7WwHX8HJ2EoFL0ybGImyVCrjP4qkgJ6NkQZCNg0C9RvH
yD6GP85mt/ww/+ToqqtmPrtBk0IGLZUTjoPD1zfGXLpedTtVMKZHxSQwN/4ziO/4GmDh/9S9HRf6
P4ZCHSeGhOIv0CF4iD2xFiyHavDcojaIooZHplZAnTuNong8SwpjVttiZ4En9H9foK56LzCj9h35
4UbW3UfDwpyRO6Rrdja6LQm5E05K4GiiQt9sZlTgbKbyuxxWVwZjZsC+0MFroC3oUud0wFVcL+jU
UKAqIjSpHCEX6hWti7qSg3DYLeB1b1bTwr8pvqHnBmcVvAKDI+L8998sTuNp6FYCMwkfkwpG9Gr7
JcHAFqOCgykhJpDzwqcqxmMoFkaLYCXbTNniNLejChxiI5UzUfQkMh1Aaezv7PF7oUufvpvtWums
vLXJUy0P4H9Zfl881NhBXNu8Z6LZ1ZhsqNpq7b3kCHuvCJZjSwoMdwCuyxJcP1Ty5z2hYRuWecr1
mACu0klnYtmHiv4V2qne1FQhwuQANlCQkK+sXL76Go1DdkpmHcRIagPPdcwbe9E2Y6o2QR3oUJuE
AnSWrVRBOwhim1y8hYe0r59ZTFI5/w6VUpjlzalAUodBJRy6fBCuYyyAhsnmg1oWCy+mIIJijZ5e
4r1Enc2V3udLCRzfxTvfhQ1ButtpqIVFfpkxKluY2rmH0SQQUMiWFb6d/7d9LVzGctbp1l0hWVs6
QTJ1zEw+L3ZhlRruEYYomTsIaTUXTcAlviqeSt5VYhv9bu0DQJIor67CLZD1U0GgDTOWDusevdO+
3JQSXShV8HVLSw+F0krhtHr8aVGFp1FqSnlfgqugKPX87SGehd66UjXllmP024DMKaRGmwpbJXWq
swLWKhYFEe81QZ/StqJ/LjeJffrknu8Irubf0imf2farwEAzkKlAsBTSVQW10VYk9tmC4lDmbKZJ
32/IW6HYlUf4aL46e56/71wBzfFjqBk4M50M+GEndt4VA/A9BIWkO3YNbCoqBp+YxZsNuGNqY4vC
fMpa3u495ZwYsLBlog05ElxBpsYYPZo5+qAz7yo6j/7DTeUSvtNm1OhPDLx0ia+aLw42fhCA0j+s
9bW5R84scnIJNGLzaQVXNTtxsC/+Y6Kqg0nD6Sc9g9P4qAqDPRrzCFnRfn/dKR3dFKwNY7CpZrWa
Fi6JEUIUI66heD9nOLPgM2850oPCyi3oxq2hP56ka0fnReBhdOLvx5W6hpvkqsMVHdVKtES/1U9p
7TP1GUASeVJHkFxLY0sQKx7lX+kJmTvhmla1i279GJPXBL1CtYmBwYz+kXoPXMAiA2RUtVakSU/6
QDnAwrpGaGKK5uv4l4f4O3bC1MOUKmhisMN9mMfREU9nQDR9X8OeYBb8zjNFIt6dRED6lxfjqknV
1Ef1wWA4NapnRKSOTIVGiS5JgCwU86YN2Hq2tojEQMto82lP0Ss1AknFjvAINGcYBmxEF4BOb5CA
ybT94ROkBUipZbJTvSD3wonPXfplh5ZtCKIOp/fo/kD2ddwbp58dgzMV0NPcT8iD/qNTU2AlDwVR
F5LeL5fEnKzcquLBF8KNlzBQKKo64Jrrhx1jIHMxa+f9I/hDYff0NZduAbTw8XydvJhg5+aSZbqw
Z5+Z4jGgZSVPsyXoucCrJwHa9qH4UeLS2QsAUpZCL2Pk7vjJ3w+BFc3ovfENrqOzMjF6JHMTHFCB
41Eu1IbjQ+kZoPXSSG9HSmqWVyrep1TVtPGtJNjZYGS8F8Zku9Qkb/O0soeTaqnjuplIDpTQcGHl
Z8SnHRGGYLH6bwK7pidyQsCC39RxyFDATcmHq4HeAbN6stRhwQb2NncF6gIr5WzMD/xxYO7PSxNW
QedCBjAxOiFMuA4KyjAWLe3qbS9xsfaCWQcA3HETR51s2lKpykFLVNJvlECUCVnFNkt7JmRRkSQf
p19/k17wRAostXOnrCrsqemBjWcvBDvyX9HDsuiFGCk9C7q8i+yUJvFEX2Ul902CBj5VL2RdEmqc
lOzZcABAbLD03tqaYOXsWSS9vM5nJ5pntHjtfTu+AvQ3r2VysUmx7TcQ8WoqlxBr/3PwH3ppzwDZ
Q3tK7v2Q+3TBZlW4xKJFCSDvDeTFsGYFSZfYFJ0JoVbp5hxznR5FeonP22VD6D6I1yA4VKXetgW2
KGE6b4vqXFnkBjs/8CmgYTlBm8X4rjRdxeQMLub9krbQbSqk5i0Rkx4Vk6bdM4HuyCiHq6qeXi//
qBQTEZxggeIzQ+EzPxIEp9gAzCFQVE0ztVV+AuqUJ1EQ1yDzW3ojzG2sabdDgFcIPfR43rNBn4+6
GSftsZkzO9p4R6OH0F7wK8xGpk6MliwJ5mC0TODmqKRA1zZ5387WuvW2qcC4FQcYBgFPHNb9ZH7L
yYk8VKvAvRvMycgYE/ZaOsMZlFPwSf2XdSgWIV8lVitByBB2PkAzz0+YjQ9kp1ng4CZZyYjDP4rl
ZlN1tf9fEOyZsD4wLtGB+DtxaGYbe9PubvKRsi58sk0dhfUgQqbwoMRFSUrxnqkyEoIlB/0hJWeH
CZiy2xjz7iznxDMmA8vgoRwbApb65BssfjvuAHY5I8zw/MVRNhexB5APsGIdkgfxDeVcZ1f5CqZs
kKYThpl7UUHG8uvhsfmCroj51eVjuaUD9f7Ou4TJGawUgXwy/MBhtnxCn0pQ15uZjyXtfCWdMLnk
bVEanry6RBenhvLXt+TcCn5IPldhDMzgu+DheWoUwpMhBlaqncUuUiIRVx7ddN46S6xMul6jK4MK
H7I+NbAUw2xG5Sy/jTcM0HiE9NOxTOXHutkEMKRmpmSUCGS8XiG1PwZIYPftXq/g0rlzeY9wPRQV
1latSZyBtI9UgH/Z2ohlBbPvxTyMOJSyOrhOSiAtEKgENBC31G28F20RfwqaahWLOL5VzhbgGqvt
lwvWqrh4Yl/TV2yX/+jNqHKxCR7O10IzFddzG9xDP+kTtniPnGiOaxM4B/NKZKAVBlvUQwMesQ5e
tdDABExl6GrH45sjjPahgS0yo6CYep6RhcDFXcrl90Kem0EtINFeKLmv1dvmDpuz4U/igcsOnENu
5tSnhG5dwT7bZmU2ZF6tzB5ZUOXAmwtrHWgD8B9X2/z860SjC476R5WI/w633PncMn0/EjlbT8iC
eSF4aa97QHeZoV3I3Wu6fGZOkJc+7EzZ0IZJQ3pg9VAeTds2J/R7Zr2xD4eDJvTgtk+NilZh3Gvq
6p/vl7Q0aSgti5bNyxucUnqVH6XgQnuUqQWFCY4YwFSDTe0ejX41i5fzfRsx96PSkow7q88+zFIh
kPTHlk8covjKtpiskra1wtJQkh3TI/7U1pX/6a5EAIJgNnDpWZp/T2fqH/rkpYbuqea4fNsc9k9x
va4uBtm/j16fTOcrYH4oZJb9g9pdmONwFEQBKub7B/p7e3vumNDF6oNaIgyCUqdzNvj2cJx533j+
RUe25ffWEH2lTZ8P+ZzR9Ew2kQ6kfz61tpl5T+ObVWsVRq/XV1okkTIAp+PMEVyXQDIKDZZdNQu3
2YptOJZjFPt4O/OGRlSuGeDoxF4O36qlesFLX6IzHkUijLe024jpa8g5Abz+S5ofSjiyr5/lLP4P
naKOEtkhabX0b8UoynjRsL3yL5P+rEXkBEwN8mfj+ckeAI4eOQLWAX3ftjyXrP2sERb90PT76IG1
1YHA3GrKRpVysyJary/FCqmBbguvVyYxVHkzj89dC6itUq7iSvv2F20l2W2awRFqqtwcBYUpod56
g1vnAGA6GstntFetSuuhPDePvizje6OnY1duR4djiLZUajJcmpm57S/MtPsWo26VUScjiSIdJeYd
GYsebPauK9jOkyMw5LKw4n8YaPoh9lmScXdXO6i7ZnzQdihJqGcE0XuUqlP1xjK3uUq2wSoxYgKP
0Kn48k+sR0zSgkuxVIJ2AsZvW95tGKIWImVOxji+t/rHSoj1HuUG678R8r3naBDbM5gofPwr8TbI
Rpr0kPvg8RIF+PBkDEA5ayLzIkyJYeCxJVrXn1lxWItPffLgjLW6IA12pBHMS5vrQyDKc++n0CIB
Mr6tcICqGqZTm40qqN9xhYzbpL/uH3bTyvLgMab++lwVLnEQikqnzHzLhjxLeKaJviaznPmuOQ7p
dRMiGWx+URockHVLS11UyaKULI8BgSP0wzEBJxs+ct5I0hC5chM6/nmpt8794EIPhGn6cBl9EY0R
nAT9QP/Wf8WEUpquuXR+7+kTPSsDn7z8mu/0lVbPoEuVn1H4HJdWKuZeox7HkYAV2YJJieLUInHj
2ukk9Cno06baoveaCVSJAqDdo2BUmGx+auyCEr1UMqRSbF9dDGAngBSuuXSF06rShY8DRp/YG3VS
grSJ15Di2Z3ltO3BLhXKkSv2H3tw6nDudPwJ+iBTj3/BcODjCkOiH7F0RrKOzDM/WOQiG+RGrfne
yG29hJY3KWuKvGhlAcFfNzoqpDs5jc2D0oasyB5PSgldW+1gTAeutsyuXW+GsqZZcvQCNr7JDuKy
ZVUg7xIj7JC1HcijHkVyO+6I2XzuQgnyZ/7zGVSonr76NJcMZIcfeyxo/e1C7R8qhK691UT974f1
C4qcLwDEqH/wXa4sQzTutY2A8W7szeLQac3C26jM70fG9Im9H0PsguAJanWVKGFfI5uupBi0lqNj
XXhfdff2bGpmdyrdSziesfNXTjJKKiDBDiTwKbcyLhuFEqQ2GWL+7Z1W2ZcKdlTRo8dnaE44yzsh
P+S7CmGZmFv1zUW7J3+nnKrqy+mESlTvt3MBa354NxSbQ5U/nFTfwgb9/LbsnJHJEKg1Cm5RPMgy
kgkA2OzyDUPbKnDs36byXgldiEMEaoqG6t6if6uNPkvQto9mMpPmikuWI02AlBLq37RSI9JWMaON
VImmCOSKUaJ1kUgan2yiU1bBadZSqBL3snuPS8mrSr9MYkgmsqcY1QpcBjZLXZszs73O5dculVyE
hMticf70M3bJr3jib4BAiOSuLpd+nWxN7gHGNdp8BAf0+swgzvViZukOfJ4+J6R3MiD03FKZ366d
xQbm/cPU1Ok8wGWrWo1/e7xggcoID1ZfY2ZZXwIkARiZqozJdGDrX6MS5QTg+BoAOw7a5MTbZM3D
kaAGdjn0JTmf/nDYHlIkIee6SC4aBMp1TB01Oi5Ny/HTaRur9cM9a/su7IkW7zJLV9DngvwDxAWJ
BGglcJse5RUhu1T8RNdqN/uevQPcnPPyOgd+Wpc/WjDE923Ypsor/S1F6ldVKNLCxwUJfxpzyD3v
2+eS62CZrO3XtjBP1Y/LS1von8ci8zRk/pPMaPHSd/6z4SCX42olkFk4kt/LxFO0dFm3WUOHraTP
4Pg5MkSzwJnLj14yj7p9+EEu5uueqA0QmJfA6wnF4st07tyy4cdD4KTLL0ioijrxFCIW6WO9gBJt
v/z9Pq4PZ5jrw0DcwYHgshIAM1lBRORezOoqaPl3AuUuErncBo/3QDd3M19dZn/vMbRaGjOJFkHd
km3pvOjqXoy3G4GnNAszbsNmPWBdi9OgmfE+c/DFv0G4IWX4d2tPfh0r38pN11DVk2r0m4KyDcFS
ujk6BbZPRl41hvRyvyqv5IrMCD9GhIa2ET2Q47hmuUzDhlvTdeRyR43Lf2Tnn1E9EZXUS/TkqbLG
xzTzaFOCObANdQFS/dVG3uBhCnVGZofEQXJhLTYiqhqoJUNhb6+5HyaHF561zcKTTfQNS21w6RnZ
siOogSgQmYZmo1vuzcGGk0c3G/NCDrpBfa2C6kEeHnz4kamBPBclKJkUbnA3T9/RweJxPGHqnGkH
s/le9m983aiXSMetkW+2SnaQjPBS/Tj+JalYWC1dsAJh1V8eT1j+tj4zRX70cexr8wOHu/bXn8T3
XohC2YlFx4i6Nmfn1eTuoliHFrrlBPd1e331c7GfMnIryjCIm2vy777yKMbQoYA6nB75/rRAAkTK
xbObZkT+vJ0QHIEqGX3R8prgTcMPCAS5LtbGbqdJDATPbOsiSf1qwk1c6n/SsN+aOC2zmT1PeTdB
QAauMzfsL4XIQuGJYfaZ0ug2h9tTdv4ryAYS/CJRlK6Y5fWkzUOVfLBQC9e3LtIi95rvL3hkkpMM
oLR8vqMnsY8Ktn+PCSsRe+FH0jmjXHkHnVB4XSh2JJsQdqVWTdakd68jOi0hfdxlkcPlNvB0I96y
dXlxmLuxU4rVeKdFOcqQMOKuWyeXfUs1ai0JrYb8A3X16nOU5NNNQnf2BOBkK2oUrSVkBdeA7fKG
H7PhoCz48V6ViXj8etbVBNeZ3/tfEbIT07rhcd2EYwJmpv+NuAvxZn0rr9dYj+i5gGyUp3GIoYdp
5n/oqaA5lQVVOGK409VRgv8XE5BwWouHWPC1BdQcpyywknmbka+mJRJyBDu0NOL8oipTO15zg/xT
hdZTKLiWDIY/3Cpq+2/KcL//eoEwJpwy3JAvkp+QfMPs62nS5O6IimsBMGeovwsbqp+nTXYunpOv
O7s8tCBIeDJ22QbEIKm56hcsdyZXBwpIUQYyqVXAdrRSa0n7oxSodUgP0j/W9NQ8iaN0eMuKTzRT
NqqAetdhx3/6Z1u0NXttCnUqpyccko4W0vloeeocXENp7Tw1wLUL0jdMBdofFP57WbvB0dUIUGvd
HgbghOYNGG6p5SUzLy5Sl50tLXd4ayyI3AL6RTKvjGBNG3TvpE2Holj0uhvhLPu6wwoLqwEQo9zK
5L8NX6Mcd2y+lbXNAECuG9ZSrTtnCdrDTr8rNE7kIHbZlD9XD93vddfLqtjiJ3lcVyotVsEfsdmU
ZIN/pNSWVu46xCe7nCL3s07UszNf5HWmiV0yNvhLm/6xFawVJap6DmalMkvXoZ7969aGEF3AKBOM
HYY2LCCLMTGm1uMBQIr1P13w5Ee9ryRo/51fdfGqlm0SPPnuT06BNPswoYwZpEgKA/5g8Pf5XTpu
DZtWG00F4P9N10N2VdMcwmmjub3CkfH/mylRhbjZHMm110oQ6ywIH6ldWDcrXQiK6b4WWX6NlSab
eOWkb/pHajLLva1qZNpFq26MOggOqlBRO3nN6z2uscrzwQjvJTLeWe9TPjc15126s4q8vCgwcPTH
ivuQpRsGhlao7gCB5+Vh4hdY4hWtO9AzfUEbtfiFA1FxAyXD7uDwFZQdhdaahP6dJJMJj7M6hxf2
xF5bX5gaMyA6tJlE6DBYee15/Q/CC2ctzD1Z9Kqy6S+pyw746c2P93nUeUiwH7I0qmBuGGI1ovmD
i/Skft1i/x9SOw6Al/WB6S+TYraKBmK37WKpx3CoMtS4C5ND1eSUp81z4++PkUAdP26soedhstVs
Cs7yto/6JqD9Vqqe5AgsQTc7IFRF6Pr7CzFS83t0zovE8CSkq+SdWGjjwPgBL63UIYyIHJ1EL3dc
ow8dPN/kI8zHKQILCnT44/99E3GIpX2nmPeQixGhf0wk0BSa3/C3BUm1A4b96gLods6vSURxL41R
unv5vfRukw+6N3gKaoEa09e11h3QGAtbNPgFrN2R0wpmarJvWnAOyNZzf9QBuJZixCGue+tdZqm1
AcGqz2wgcXmaAPV0qfcXUzPgHpKWqqF5F8AQovUj3+vnmxACLQL+nvulYDIz7SWs5z6m3+qLmG0y
7+q9E/t22t8gt7HTQxqPA8ZXAzRE8sY2VqLXK0AizgBEasLM3lmBN3Uu4efGBk8vYHeegTfx3Yq6
gwLfVtD/kDUYnyO0uNk4OO+kDV1gAH1gA9N2BBL6pPtJgi1VvOBJV+rA4x/aXap9mlF/GbJXuUvM
nPCudY6MZ8c5iZChfZlS5CUJgN4+fPsTQgpFzLA/GxBeo8834re6ZpWUMBxVzJ2bINb/4EuYW40B
Bq/+y9H5/RvFSVD9DQ1/WSehH7zk/U80+ks8VzlvMlkYB92d3hOrufChWI8zjGQu46aNG8i4fKLC
tnGG9/KpQgjlgGCSpTjbLAFNSIoNQkFO/1QJZMA6DCLl/P+2zaMmuyGuJarvNV7U84iSegIe4WPI
E1wbHoUoM9NIp+EU3KHn7SjUS6wxNwrecFboBHH8DlbItt327+WwaiyebhkerpZ12fGyGgGvO4ro
2CkUDzaP2b8pzhGwHFSnLXXcDYx4YMSf460mOWXbUIshX86Y/I62JXLvCkNnlAgfRPPX/HYWQwk1
vYTtpP5OoYeo4V7PAiXKerlrvziCkJUVxq3pIiRUfDTMGickag3NSo4mVi0Zz5uYH6Cj5RNYmAQ+
fP76B1QYr7Uxhry7GAQ9RgB/QUbJueyQy2iJ+JRxtI/XkEmTVPWd5M6BEpRfyZ/2FgZoEoPTV2dV
DuO+qo5JkEfUwVRg+PvYDEZK8K0t0W5gNLnXjCo0J/HgX8rr/f3r6djiIlA+iI5+91AG5zbpt2Ev
3bH5rhh7gMUGIwBCw8Tddi7TPzXsGvJhPw1Mwdct/XmKH1yX3TJgQw8G7vTpN3JhOcfsyBvnVzXa
jWhJnnvAFxijD+aeUIXTmzItLMXw6toQB7nv6RtZLoeBn6xdF83Hw1LN/e8Mr0c66UwtnEuUm3dP
xSz0rUR7bB3w1WC4f5E8if/X+HkDutzPyGwE6mN7qv23nkO0AEsoPD5cHcCWXcuqMjLIBVjP9hxy
n58S0BxAdBAQf9j6AlkMTp7aIU3Be7KNE22CmLovyyfgEGRNQkvjsWzDomH4z0HoCNR3+7GEhs9L
l0lvPjsEh8TdEz6Dgbf0SqUYszICQajwruSvzTsYGd/Q/kN0qPdktoTeKZFv7qNg2j8XMLwhvszQ
/5sltWJM67p9tTi+UIGChhr8NJwpE7GtPx9VGSWQCxHRHKxfm20aO/DVwPGqBJBUnJYZsg2e5Uwd
JMDMJvafTxzK7828xfGtkpq8bTiXO+0s+MZSuyCYqSvVAu7xeL3bGKdGVSKuXqWOeADxypjC7gGV
sLSlvJXkcQqOnISu/fgSHoqS/ciCZT1mJGIiV59OKZv6c4N9uTBYkbx+DP0Y2A/AzKI0MIfv7VNj
1cX1Jk9GA3CMTeFfs+wA6tSUq7E8WWETZxYNMkCEsPPzYjwOO5b/ql206QIT1QtPqqoWUZDvkit0
3RPtQGP1xuV60lzbzTgncOPUTtNwvEOq6utbjPn4V3PuVeejXZhtqUTZZ+/Eh+sXOzWPlBEylpAl
PzzS8ApfOg+qImhEOW2391Tw0uI2aPR+V/pwTlv2GSUEZQ11hAsTeCYukcxhKgUXzSYsLRheyMNe
uzHl/MSVKSAnpWUYuhE22dQw2nNm5oan1a8J2r+br8LuwL619tpexXn8I5/Pf8X713pF5JQS952E
64XLugHmbp92QnSITJRh2roFyXjpTKPpdEpVvTcAuLWYIS+KSHx2dxKC6NfE/6vmz0QzIl/173bt
ycMQHlgBLlxd9utugjmENDo5aBqx4/HbUX47rtvTGvSsrqkYrfWdlO/Fe+sWP3SppGZD0KnjMw3Q
kFOgR6Ho1YzehmSkl2ObVoyIsViHG1L9vc2R3iZ39QRZ+kMghITk5U5Cb2KUe6c7+w/GdFZiy0nB
fDsWfpmdqXZ3Y8FS/80qc7Na5h8VWZmv1BHXGRyCWoG92FREMQ/Q/TOMWrO3qQOj8y1lIyan5hQl
XGzBEQtofvY0JONpIBTlMkFaedytoP//H2wy7bPW1MGsZEr8PWE8v7nFAks0O4DmuTTi60l9ppW9
q+99u7P0D8IQlNnqSaKjijaE/aKvdxMwQG+nB4WI/TJxXc7idc5Dhx05rwcHPuorAbx1jqMMBxvK
2NeUwL3Zc2MAK2BPbuURz+dcd5vocch5IQqyzt04a5rwnwioOGdqX3/v5rpvXCmq3P9ZYgDkScEJ
0MDRmvNdZwJBa0BoNSbyyGGIWVTy3kfB3w4fNF6iCHqWMqbMUb5giSyzqxGdFPlVNjObosFnDSkl
oP+PhxQtiXwWwGA7enPO2OS5JWY/3r/hqIo5NXzA10icr9jRcCotSLh4EgPZ8U3URotR5NkX/KN1
PMgyeZY15wd16Hsg5wSBvTRSK2E9qRRH/WSwFDi9GGC67r/afOWDCvjmJVLJPdDhhVHhs2Zwz5Pe
3b+pf1r+tUyY98qxYOxZvBmJEqIGOiwVc8pr7AlmoFzKjF2hSHqOixNcZDbUbBQJJhVMqCr4P4mc
RoMj/5pj5YvQLsI+Py8VMz9z+d1bw8ilfVEH5f1HlAp9YshK0aYVHjfoYxc8oh8X1zvBA2A8Oa+h
gCbZQg2RVBVJEbl1hYEi6UXmzaK1WyTbVK+6FVkme7UVZYNOuwn580ujHf1OGrR/VUbiZ3MZHvFm
EzRvft5jJs+DI4v8iTMJDbQtxJsfbsYbFYgor9u4K0NoLsDqoZpkYKdzV4U00hvFe8Mu5HwhuYwu
hUBz1ZvPi6ku9DlaCjKPp7hdoDPlOS6ax220jBWne0ZcV9lbu7coiPYho9efMxplD7/6ZeLMN15O
l/HPpwTvaU3ZGIGAdJiqej8M9p6zE7SAh3eI9oyIgPT7d7Js6w+6GvpyNK6jxuCY/oyfMN5qRs7X
JPgeibGh8+2k8Xh4aYr6GqFqMQFdPllNXnH1qwaXa4dXe5rL4GfVwrjFMrnnVho4uH1Gdn6qnjBR
r2s73BNrYo8qjFfrPqHtAlDhYDQ3WC3U8ntSW49GODfJzuFcJtWxDKx+xWKBfC+a6mlOBm3GfnjC
R3HSg+QHjAbFSZVaer16z6A89RqooSV/B2xRAopjvooi6xqPq73AB1E4vbF8aHn8HXB/pDoFsRTM
ur2HNxMdJNLUL4a/KO/H9N16eOBb9Uv4FXTYDxC/GUvOb2SXa8AJSsQq0aGAdGaPtlTfUBt8+Hx8
we6DA99Rrw2IH04ply1qQuYv+20O0L+gjon0uJSzEND9Bi6JOp4G4EjTNbmoLDv/wq12KrksR5QZ
uMS0KpOtyJ90hxUI4qcAUkmuPIgTbKefmG1iIaGtzXQ1p3I/pt+3fQlkkgwDSR33tZnZV0aWvHLk
J6rO/Vacw7yL/cAV6aMzNrcPVt+j3mqj12OnW4ScB1DWOJrZEosdHX5PRMSg5Vm0K4l7/LEzXH/z
5FP4NnI/ovA59+XTYc9qJsUc8Dbo8MxcWaH0XWOV76dvC2sj1TRTZ4z+ojpdOJZnEGzcOERiiinF
QBdWKiC5SHmcUygoOiCPiqFWEnfixIbm4DbZNFSVb6s4x6mJEUbfqwmBDYznmVy4S66kFiJhyKZD
pU7f5pwhnpsQrSfNYflBZhToGisxwCasrUYOEy+MbaQUBilegb4nu8hNAYgOLEPSlmc0xtjcdYsm
t7rKY3r5m09mljmHQMfWVsKfs2LgIQOyJ9t7E/mNpa65de7CnlbrEDQ8BTSzhHYHdj9/m/ej6XT7
vF+4mrjDpJ6bzEyJKJdClcWCaL9+4fom12OHscZHwk1pBvCk75d3yGvH3ORDd8eQ6H9BLDfiYVhY
/AYhRHPfeTsSbLdZHILN9k5j0SOQ+7OndzjVOCwRj+Ik56GUnfxhQ/fbEGVJ8Q8hUAfEyG7EMVi5
kJA/tm6jS5iUAutWNs9+bswMBtmjC25t685fxQEImLdk/m9Qpzm7aaFGBINDI/yIy3K70To6Xswo
+BpnPRaLRtQwk1CIB1ct5InpHXiedFfbdFClIzvCBpeXZp/DcVcMlx7CrhqIIG0qnz6UacVe4FWT
TnumRIzBmGm9IPW845qfMw14cx/h5o5L07F5f/dThOlLlhj5Xp9pDhbM/u7nSCl5MFcCw0kZwn9A
P2I22a+1tG4xcYDdhpp4SnEe9984GcS2V97iDWWCIfi/394sQ2HtjzQBzSal5uY1iq9yqdz1dh2M
0t0WQZE+OSYVLikuap16AlfpmAY/xBkruZMcNV06a4nLMtI43PJkCepfLA6lbV/LTRwlbXidAqyk
n4yaPKRU+XInmnR8cz27GqVbt+YBP1eT993Mk/bb8tE1CEE48QLriFsEoCratYCuhZ9fVQ/CbOSS
Y9TUnSTsIqAv1ILDHbTilanIgMfxq3hxE6cPV8F28mRMoQUr7+j3Ps08J8acGgXo4XYmTUwn36Xt
56yxsF7bIXD2/Bpkhi05GwDmiac3YmSX7r9M7bKsGcSDhce80+TXGWAK4ySbTd6rc2AbexmWpS6l
0HQaV4qKyHt4UNHFgxYqmvj3o/ASWMdp/EMngPVEFO24PRBKTuqTpyRFLAzZHXmNiViZHpSlT6JA
selVqFV/KEyv8g4A1L4aSPmcyg7WQdWhTlaUOUFx5Hfy6Vj5oypR3PufcPazdZptSYhsOhO208Li
bsyfHQp8RYpU6sxwbkZSHER124TFPeg6oLjDFGGGRSqWGMXm22pFjjCElAuVOsDrWWdZdrqX94J7
A5yDLfsOeOzJX/Cp+nBbAFzJ+FWPitUEFOHT0sAUExkwx86t3VnKJ2iYPBxm9u/Z+YxLeNp/ipt0
Kwa/+sslukoriCsIbdOF9u8lCjfNZN18NG0ylmIE6XA2P7gYl6HzkTEUd85+Pzg6z4L46S8bEfyG
mgPMHE+jrtc7Okf3L3dhgzKwCbBlMN5tV+e0qTa3c4lxik5Ew3yIabytcVE+p+ZrzZpc/CR8xDKT
ua82GjG3GfPA45mzk1BqVS2VWpWrYTBeebNJ2CzKNkv/i7rCdnx1wJHjKqq+MRReTI0mTU0ba5ss
EmLZhuk2Yu/nJMzgl05/J7UMRk9cj1gqe++TuqlsCmJ5DJfBI2wMuP7TV4h/3P6ehbVkBwNr2nzS
X81iY5vYrKF5qblt+UyzeKP6yQ6j1DOcNScmFueo/taK1U2DaAFFjEXnuf5gbz8HB1WesSMgx5j+
oMjO+kp0EG873lxkmzFGu2LDST3/QYzJ6lYgwVJpzshQdn3MlkshNp4n44TK9Fsk2aogMYVhJV8+
rUHt4Vm/faq9FrGDi2QiQd7H/FTFg5Zm/D1z0uwzsEDoZdtjSHFYY7q9C1NdaR/FwdxGqIdf1tmU
yahDlhQ+IrAm2QbeJL1aib+Z4RoNxZbA7+Q5WX/Rz6anfwOoN/O4tvuYFb7Pf0TJnsLVG3CGVJc5
aJbS4v7a0+PAyN5h4z4ABTWOE89cnxf9yTCMoHMSkzkSkAAMenZsAlKsQRk0mhmC/y53MhP/Upeq
M0fV55qWcFbDuoQqbSafPk4Pw4Z1ISua/4mqtDas4OJEa7cwkF15GgMCzjzu6MsAAkcWyi97f7VD
xBciu6CGSVzIGA4ASJpuSzn0p98YXuWnDTy47eBSCsifWuRxfq8uGLbYV9FZ4s1AeMfch8R0bFwM
iBvzMOfP1rIuI5VOetBdi0l8u/RukwU78KgBjeVfCnyCx4cFD2lAH6Dw2u2tNv8mA17X6Ur/4gNt
YCxpKCZFB1pmeo9tJ95amMf8Q+/nQ7upMw5DzNRLES3LhhF0WA1GBAS/j6v/IjLb36o5XhkL/wm7
vhsXI73frIBR25hB17C6VPYX2M85HqLKXPknDD4tZLDFJFBaS3WI54vUh26YKushpsTrbxcEaE59
IfE1YKFUhDIoY0RVYNUvhTsyeEHy/6LMt5Y7hlm1w7eITDg/pC+yZmSE+G+IPwfYN/IgbjFawkY5
2C7h7TJknKfBORVT2lHj2QNUf/DTRXEJRepaFb5fZtKVY8aeibHzx1Zpg6TMSd6ZFr/NM46eiIli
NztvF3W1J96qwWRCzp62QCa2qoPecq1gJaSFAlZY0F6K9jTZ79WZeHpAKnx9iMYThMaED70Tzut1
LRPOu3jlkOtF2XMNjyFdizoqr1EPZ2SZsIPahsVXPySsy038y2MnemLXP2WzinhyDJM0yk07lM/s
09v4mbMnGEyCLGt1ah53MlbpsF6DId5a0SnSC6/2kz898S4HwH+4w6yAvM4f3O+S+nYVNkB4Cdmd
+wZjPOB9A4HTg9pUOXSS+a31mXFNrrWUGPFn4k+oHl98nJX5rOoamhMv1886AdicKcCWWiT6F9Iu
k9B1OPCFHFzMlVZ04fYWSnys6GJStqsu0BgUghCRoj7znMI16SpCAuT1oDvRSBiSGiJHwQT32g/4
YsGLfdGzPymgWaPkPpMN1r4XHK8D41E90Qcvzthi2rz84lSTDF3ClfSV+OWqP+71UUg4+bEVcWGw
JNZl5kr37S3egNyib1fbtfe/ri8tp8e2d1LT1b+2KRcJ2drGYxGgEMoVHglyNUJ7XDXD7isbZMv5
EfnH1/4YL6sr3zyA8hGT92ZIcRBiS83XJbmemCDhIckgo7aIFWCnvcuuxivevJ3YiTPZtNWPGqDO
qXgei487YgWnXMBsjyjj1FT3ul4ex9HoazYY03FQ3auyYt5/sysl4x80EMoCMoFBqKD3FeNczgTd
xyaKkpiUV6kIIa+wie2ykA7JsqIfRfEJZxRx34gkj+UQ+OHsTPG/MHcDq8fFgevEF7CmVeDKSiNL
MG3RrYURlENdi5hK5/H6PX3wS9gX+oPuFd0J+3kIiQ5UsItv9p1R5zvWZ7qHUSk5lHy/0R8jMOM0
rLXz3mwZMpx3CoBA3GU+UOUWRwsnV0lCVmnRvXOfUpwtC22rnZT1srtAQ/rrzRu+QdeSHPFEpwoL
gqxAcpjWZbJE9Yxa5aAlcDynxaj0dDXNjzVZV/Gr55Hxy8FtONbhRHjI55zJ7BNJ1adqHK56oqL+
uLp8hok3f79Tf96TxxX1ArQ7RtxoQsghxaAv5MpzrvS5EiSUSc4NMFXI3jAt9YeRDmNNCxavGoNd
RrxukwqT23cgbyatZ7c/jLpacKdYkj0aZyTm80vz3g2hOzQkiG0C6BEsVCNr5YoSzkoUa9yvMjgy
WVhm/MV57de78eGsTspqNNgwPujqRh2nM+6OHM0m3Sn+qAuC60ZzcQrNAtSGH9sVLMTjULuDglGb
Z4tiBCn2r2HMQ4B252/wmTIIhaWkVoPpXgOJwmdhMmSxFMQXcJoc/QqZWnzQ3dE+7hyDKw5Tnqf9
6nL5+iVkRP0muyqi8o7ZDevFwl2tQnn0D5pRyMePKkucEcf3rj3jVEl7WF99xDjpUXDJvzujGxMu
lVuLAjydGO02iRrC2aJSgzdPYpsjnrmoGFSvR7Euys4898ui9akNoTzZ1zHcrZ4di2GyA3C75fMT
eIPv3VxvVBJpIQ0yHu8rgP3OMcAfGD1n1C3ITfA9e4NVM4UJ7ltPR0T/rKGcUat5WRhTclGxsNqG
zQG6zxRBvLIjTLsLPRoji/EJJUl8Y+5ay0mdZtb2Du318lj/4c85dRJ08vy0ysVC3Cz7Ei4BFDSW
k/JIF02dcpYuAByk74nn4P1pDuSX9B0294uW2MvC+0qSd8+bHHWLC7V3ARFU//nqbVgvqDW9x7m9
A3L2J1pRZYQMhZL8223bD4iZw4jHutJU3J0ymYE8xSZe9ku/3O+pQidJVOAInloljkesbjtKz3yh
IT+T2hQzX3/4FdhlOTaYLnSkn1r+QDCy6LGDE5L5ytnKX2jAmT70O5zEIVDzl3xOu0ucsKTS+ym8
kGGrjacbW26pk5mQ8zCH2DRN8JKcSvuhAjXB6fKffIRn4gQC6TRx4o4txrBYTGOMOxVff2+D+ciP
iggDloLdVUsoMR7S58LLtLHqHdJO/R5fjByp5V7oVqxgbnyD9WzNOvuxL1dTww80eBjtqMwV5yl2
aiYFZpEY7Bc8iADyQ/9XsJFWQRS1YpZEzF8HJLvZu8wxqQ8tFr1Vv75r41tRsy6xPFyMsV2rSXhv
zX61+VWYFvK1Q0c048nGv9JTxkT1fZkUPecfEvFvet3nAHJjD41Q8Qbw/JurhjT2ilyv3+r9lj/C
2Y78WyRViWOK0fbRfj26KGEyaVQVey1U1xrG3Ae3cxBOVsONNqyZJ+9d/LCU3u2mQ4gb1dUap1Iq
sKc/w/BMyBzUorMdMFExf/j/qNrEpCi6yFBpdJCy1NDEm7STbMzUQWvbG1QWS7+1w9tK4pzftxVT
VDMjPW+FJkCcouFH1p6SJYQgBM91ZpYbdvyWljh+CSN7boYCzkM4gNaQ2NI61topGyAWySseredj
diQrXpg2dDb+cUbGTDp0tOQzBIBjEIEv16mI8TjDpEX4qb/KRbW0qhc0W46KJcwNaTfRWBPh+Fx5
mgGdY73TmFpOdJoe1tPcnMcOO9U2b5tmL9I++mTKzdRv9FelHT9IwFEuhefwm08kaBEEWX5pA4T4
W1rLCouc0jn8pVTGQ1BllIAyv1i3k87eMD44G8G6hiMwXzAjZK5Y7Oh3cPpycshTRAqqTAb1oFf0
MFZZhOkbZWe28wX1bEbjO8aB/7Nh9baAIASeZzwC7diJANxrneX5YkCXT3D/LztQs572VTadzvuy
FUpdKNMh59fy8u3U3Dvp4UgF/CLMH8iD94rNkVVWNHNGPM9/CHLu+1X+jSmGVk9Shz3X9qZ03Hap
XDst4MY9oeMefUsgsUVUzErC9rgkaWiY6COOt9CmLijHnpGa1rL+rroRah9BOpmf5g8MI/ugmfqD
SQUN63I8aZqGsNNcemLGr0Nar7eVutaqvsH5GAhZvl7E1NLCkulLmsVRCJe6TRQlPV5HWVmLXmVG
B/kkZ7ygf4QSm1OKIEu4gUimLiy38of0pzI+vjvuFo2d4GPlrD9SlO/VzT1jibz7kdAcyVn0mhuJ
rGy4c/SOUfvGuyY/kp/5Z1iBvq4wqLhoKosKSUuIogl+ea5p+4vZwDw/aodZcfP6GTQWkew3qqjU
Sxg3kIBbzatx6BXCFTKND8ylYLnEO/uS8uV/m2lazGrZDEu5QjM5DuJ2ZonyTr30irixea1dUMGt
zsE9YUdMNOW1u+RvUryh0OJdIuX645lLZpDcS01GJjD9JhSxncddkj3piclg6/JesfHRkQb/HQ0T
Au9onClXUrHcMcyZT4jlnkOSuLYeKB9hq287CovgFSK9/hCTSwgO5rFREDxlxgVekSswIBcw/ZLk
+hW0jtsQHvKPdHwXe1GIaNKlGCOOTMJGkUuUtBqS+0Gc00v3eDKiMO8pia8AaXaj+RTFzn+yxpxE
Rp74lo0ERMIrBcanUdAWAEPm+5257c2SHIZxf8gu0puHD2i0m2M4foHAD9+FEvj8ujSTVzELm4li
U9nWV7QyeX45DR5sy/nXffHOmJVwFsyoSBnV2nOY0xOZ3Yu4Gn+eU1WWa3Lbm60YIPuAwl4PIpIf
pIsNtVIA0SEMg1hKcqArbpBfpyRFGyFk5HskW5hzwiHLAZOL3L86hLNkbq6o2oe1FNuwzVXYv2MG
F6qmorjGhRdMBoGGgfChQeUop27e+30a1W5upnz8RMGS0FxJ9ZplHhr8rPaLhy4OQkWklgyxnQ+H
nLizGY7gHAxkG/ovuvV75DKUjl8Id6i0C8Iydkgf1JBBRNVBOhxeYFaB7inYhbFEv8NwhXd5GDQ2
q0XxwkhwMXqEq3l4n4t4Q7IEaxDDWClTzngVcPTEBB7nbVfvd8hlWcq91YihVrIIth0n7UU7Ove8
+YfoFTv29CtraA1pn0rJV7qsY6IV3uVKnNVgZzeE1eueF9tcTmIh+cSZlKNE5JzgtgQTYgsM/6AE
hY/86g2yf8YuzA40iOINFE5bpsw7OuJ58cnd+Fjzdd7SjV2K8dVbZurdVH0CXjrgJaqflL2tipGI
wbUVAAzdPBp2nV63PJChmoKrbmgEorxEiTAtaam2H50jgLreUCeCDODURbzrdhYv4z7yOLWEPGKL
0DKZxIxhtBIbcKhK51wfic4Cmq4WhtBhMKnGoBLBRNnuNy80SaTzWPZ/3UZ07/4CV4I7jZGyXfoQ
CaBD0ITKHpOgsb4C5iyX5VYrpk7WnmBNtJCFvyqWll6EAGMcnxQSOkgQ4yYzP6AFWoPz3dWgMcXZ
0G4TUVFsf2MfIq5lwwKRTMcjhA50sRrZ/65XTX7EXCwEQ3bDoTzpNaycfoIFGoiqBWmxOKc1Favn
EHa/CP1BAOEIuyd+jdFmNZa8BXiyTcqEnGRwOf3y3kWVjS1R9WbdjJ6gKQq6n74XTNgLHng76uG3
aYvIWWMvNTYgxjh4jSNRzUXnCo00W+QxE71EiEuhkI5NaWFqO9LMW1q/2Oh8TL6oQU1QxsDD7Kqm
z8TZTAt0wltBxrtx87JqR2cTEHFCiSNBmEu27Ff6yo/GhkZnhNVPD3LCB7BXBfFmU3VzwjaWl8F6
XH/mU3QmAG6BpearUJbgZZLmQUFbiPEuAXJ2PD1qD9FK1JoO03wKGwxz/3FfFKk5VNtdNDPI6NpT
xI0T93nKvUeUelurSgO/v22lLtVIDUniSg7cfQnNRDyv6kmpGGVdIOWPRtSnthxi9rMGZHBhRymL
cuNfnvxxXScIvFwK6LCz+9UJpebr56eP3AkZARLt56DKYvDJfd0zEzSFSZ9PsF2WbZvPqWS2c/1L
tlTHyZuOJbDLTFRtWDtVtUdV+HJt7qQsKEcuWYjubGQINmx2B4ZwJdFA7pAltntwowWIC2ABw1WH
NAbvNO1vyqhSHP68vGouEL7KAvuWM7V2EneTCdEsefa+HQIVrXV3hHHhaWzE22w3Ro3FvA/9lFPo
zv5KvuQg4jvC8JbTStgTGuHuyMs6NGwufVWmVCbPKmeyOHT02G7qYNKR2Zn2MvfHOBATDgRLzJFT
rX1IigqiBsXPXsL1hzOSenOoCFDgklwi5xAvwnELJFpXx5yrHhTcCzmYrxltKuCPxhWdVdznmaeR
tglI3ncB2hjXBrbjn3YF6latUX6UlnFIo8H6y4zQk7pSwSgaE+hj1AyzBpOPQdchNWwRyEuWoO6N
yYawnl0P5kUh3xdeko7KeIAYvumZZWgK/QGE0rWyn/ozmOzz0A0fdYOvbjdktVdtax1E+Yau4NMN
YoBcKdBPMS6VQ15Cksz0LMXBcwmYMVl9BH4gDDskI5J64kGVg58vLS4gcqTtzKZZh5C0YZnilmK3
X1OFxbA0dVVPFZ/tQQF8iO4TlWjj8dkIIKfkHmaJuQe3xHoy0vgWiEcNQ8PKc6sXn3jrXLKJAZJA
Xh4pes1vDR8JM2HzFW3pP/uq9PdOmSKXp/HgY0ek92HIpBkZ9mSqmzfSjp+kdb7vaXNDTNZUWNc/
jaGGEw4BX3XEQGNKqihJFrGU8yRjaiz5ykddInhjBgjFLFbCdaMuOKVmoEpJN1zKqle5SUl3NMa3
wZSs+3QTdMwPawd/PXsT2kuNCCD24w55/7cIskKWQ7DwOpZWkznJgDrN61ytkseC+5osSDPtZGJK
8+yqJ+8MiZJQDNhrJGw7Gue57tyFTNzHkuuhMnVUwbsfm0GqJfBAkUjfw4+9f/RmVo49T0+3nKKx
HTJlrFC8wt8J8ChCDpDe/OgqWRMpR4rleS3Cxh19K3QXXAOshGNf8Dn+cseGm15md108+5Vc6TTi
WaVebeOpiMHVKsUV7bAhP31OwKtxE/tT4X74C2CJilfWNDQ97jYsz8nD5CkR40ajpvpDByu1501d
MX9oiFGBi6KwwgUUkYDg27959vjwIJ9VJZJ3llEyHwmgNW0ZCF4I2D/LHhFARWKRgaOrVOYnnFPS
7Lc0pahto41Iwe2Q+ynF3W54Ew35ojRh9qOcbWkkqTB9+sNr33AiBQRqXWJlxEGB1NY28OQMfHLr
hCwfOIzZvwxa2Q6m0e6+6wLFr7g/PyWOSN2wl/2GgegX3tDr19/0ImtaoHoQGYwvTcCNWd9LUrfG
2jcydX3ZjYJShQBap87Bh0jN9ahAjHFmldrp6rYtHROEHs7C7Nq2UVsl2RXy+JprtcYpc+p3a7lM
Fd8eu+b88VHDGoegD8uS1LbcvW/d4rXFFEYEgtSajGE/8w0rB+akrEbwJwDaTCHjBYq2KaddI9U7
QnonpabUvNo5CxTab3w2hXozWFzw1LQzeRHMppH/q3yOjaKBh+zUpNpYHxwK59fujk98znjpMdY7
V+NFbBmZA0SGKMIifyIEBLX5tKuf3BVSlzcdGW22o80QcIjPqJUjCwNVt8bCmnpnQV1rN+p4b5Ul
e0uOIYNA+K9l/NidZFIKMhfZpAS5SicMYdCDDLPJp3cLnOvYT+w3hfuqFiFkfd/KnX6Xc5GhooYY
xHA7N8slbczflqbtytn7MBMaVhCmEo1fDVeb+PxQfQE7B+qMNqsu3ieHzi0qHt29ggJ5bgTTbY0K
1ivsllFwjkExIv7ijPUO5KutnDkuLxhinXNCUThYkLLyCMlNQQi4RttHP4l1NGlSCXFeQ3qMZeNx
tIXoaytX3jz+arsTxxUWdMIjrSmSrBhgcKj3aIlv0CL/bPntZcMsOtw8+jb73iVx0gzoeKW5ZONg
Npa0UnY/he1CzkxXViaNTU6LCeJyela1xtMRHi7CR9RDK5d1XTqgReZS/EcbfBvWVZCorvRFg6UB
dnnhLhNEj9C5MIGHsOeMWbrDl3h2GU4KqvorB40jeAJh+W9KUUPYlZNdr/+7lFEzmbGJcrXUbqnM
XzsZbfVMRCvjqwFrWMWzuB1aYlDtp8USX3KpGG/GtYaWun2GTKXbJtZgDQBPDxLtJhMmNfQnx0rD
U72hi22cEkafQic3zkUSwY5576r0jpU5IcvT9EnSk8vFJI38ZUHBPoCNphGC8nlf2fv9X2EB/mHw
bgQ4ZLv1FxxYO2frtlqz3Ln8qwYVG2uT+/QcIsUNvKPaFOeXVsDNxAOgJAMZ2+e3029AsllOgD9F
Oqn5NkJtMqTdtGFUuZ9uHvkiLIyAa7F+1oWL2bktM+x5YSEu4YfNqWNc66jju5KRn85DzqvAgzVO
HeA319GTxye1lmPEU+HklNa5b0h3k4sDRlnV1j6x5VUdNOTBaUYwpiHp2wV/t0UdpDfBVMQuERWx
/+lNcJ6dzZJv+NBiaJYrzepTYFF/SROjAP9GSETNMmcHHfVEiDCdn9FV8j7riC45iUKeZWMY2SZF
IUNeWLFNhJVECwVNc9n294I2TuSdf8VGsWc2pvop2Xe69VgCS9GyB8JGK8dVqsx4eG24d4lLSfx9
VCv0xNZMamFqnxrAR6+YkBp9R7Bp+ahNBWtW0+i0ANV75vtEso5dikqFWADUWLu92W6CWD7uE8+5
cEgHlj4/gd22sJKlZYdxFxVR85KnFTEX9pX+1UzL1rJuFeoSRsS7/JS9I0gkUAnV8iXkVUW/tNJF
tXSBBv5BYC4okZHWUblkNIQUwTVvX8+mnUIMYeo5WizWIck7uWO7jefJur+oAzPCHsBQPxhtbMH8
IJgZJ6+v43ycIc6A7iiuLUrc+t+vHSeWkWKP9ymQLlVY7P8N57yOpYZiW/oB/22J0ERu87E1nBBj
6sw2TS+E2wfKBGTHYpnEhE4XdzwqMIb/OOAbiEzvStwXv8vNHoK1mWbvfONlDJFnTMarlDK0JYbm
dPvWpc5hHNdXGyPS05WuMHPjJ9Usiry0XeMgpv++Y1scs51S4ZNd8pvpcxDMLJrqETejRUnycGax
3IqiMNN0AbRWfKbX5MD62xtRY03NABwVedAlnT3gTT0rwZYpnTO40POD3I1WRaSvPStn0bDjcdy4
L++9UorsIEIgHVP/mxf6SzCI4d5oHVwIqHOzs0E6YpvXeRYJC8JIwGexWjN/o/dnJXZTEGdekdTE
wBPLusU7TyI+vsN86TB0k1ydG6dUjlGgYJ20jFd56983kZRKSWSz8RfBVOIAmnqfjIvDf4WkHQ37
yLGE4D1P5JNPrKQJf1vTkB8s5UtcJ+5MeqELdL3FjBhELuAIvRpnZrDFCDyjJUeCrA4qgIFlsN++
mgy/3iZXO4UqvMa9ZTC5BnBkXSGh8a79SbBCFChTgLbeN1M1zq7L4UqEkUrIDIss1BojrqVBKs1k
zW2CYNNbkvlAfAGWt0DZ75BTpw9mi2qMFfAMRzPOk8atBy19xWkRUF7vTiliwLWqAckjyFkydE2c
ev1pa2QdALKDsiq4QNl6cPjS+/VAumEV+wtH46vRcu+kDywNK9cOI8QZCyyBPQcwRjpqeSqmKsla
mkCjcjO4t8Zef11JCot456I12TUPeNDUqKSBxAtfCn+wc8I97C8/oaj/+ylL6v9gY045mxSSOP9B
avhFqiweRbbDGOA749I/pfIiRAB+McBqm0Pq4edHfGrHuqB2kWRwo++7NL2lPKEef50QFcR4PMNa
ClDvssLeWspxdG49OEgRoklaR0UbrePxXDdbN2ATtKLP3+3vHDDSm91LmaQlCzM+AWDyUbdbgl2w
B0+mOZUECKc0bETGvSL92QVz4670kBbK+RKCeebgsKkm2YuhlfkHu5uBnzFNkQYuybXuHMbaEcms
MqAOZeSm7ukLjevyAt89tjCt22RED5wkGzDoYV0+bcN6apuifJInRy6ahZeq/EHBuqqWTmzaX9a6
S/dVmXMaWDvdMJBMJ4vMO0vV0OSoObB+vVNnfTE13Ku2aWN1xBO0/2u63zFpnG8KtKWx/JmPiKu8
DELGXnnSY2Wwd2b5n+eWnHYKJCbU7T8ZBA+qPBRFL974cNtjGm9QIwMNw380qsOWEYi0eBrFMwuq
3wS1R+yaJL5VmpiprUv9OZbYrdkBK1qN/z+N0KT2AkJNXGaMLIzTFet68VSlkgfUZaB5gKiCpRKx
5q/Lis/Fu2B5jqdmzSnHrpHVePMQYdiLJZ3z2JlK+KNxiU/v37nFu3sDaxChIpJU+P3wffaPB+Hv
FnPpzKLQ5ZnzVet1km5Lep9YvPbq/kKG6ZG61uOKX7/9NYkLZQnlgFV8yf5Ejj+zjSgrElBQ2cpB
NisueX1lg1n2rODwjuv33TGT1jlWCpwkzEGOBlE2ZdkrKIY3dVNHXJ39ZUfuzirut2DG8Lh8FItL
9Uy5IttUYYiIzuwyLGYbvyo7PbztmefL2Kr/ngk182WpMRc+OHoGRYR9dDRHfFB6PXL9Q6YbPyn6
JnuedGcgEB+dJNEquldBqIr9aZN0dVhvXj0yH1nf+4xg3v55nyCY0Oh4d0Fxt3uwQZBCXVv0FG7D
PieOgQ9G2DefwwRerDCYaZ2EILvCVORwDXxPMlD4p03Hb46ffQQJj2cxJeeos+3xsTU8fNg9TO0/
mK1GOOk/qU92a1jIrz6X6O5nG1JTGUB4z3gOzUnqnc9qa5ZMrvX4/R0XjECuYvXs5PBvwAt5GDFO
4LY5u8fBGwfkXANfvysNFzZhtHkjSfAqhJm+QmNhwsM84Ii275me36VYU2AxLNjm00i2JJJxJqDG
LKrqTXT2AcPdt+CtIZcmV2Fh1cZY4eNRxCH9A2teS2EhDJZnyCXHZAPBGyhf3dK5+kjiKq7E0NIw
sMqV/12+iYbtbo9aLUkn6qBXiiPk1QYXj5dCBCxs9AY1beCQDW4nMMX6SxbHISVWRVE0QOG8C5C+
IGldfolIxGzCXHqK0GVZt8jfJ/ZhgiJqWxE4rEatSP2IgeBkr522Lq8BqrH/5XIlxGYbMcAzbQXh
c5PmR2b6aWDA3C6MEb3QY46cJ48etNYoS94S4HEEl0bnznkN6SNfY5CTEFK994X/DgdddK5qSSDN
9IELI1g7lhWvRTdwXYmzDIA8DfLb8Y6N/QVldG913aA+eThaffinOHcUZ/hmIbClLx5cVkW3GLg0
ULtb9f8MOdd66zmaZW+3jhBERiwijU4CmxsPABaPpQa9Xd5QID/Bm1p6lZMnikNwG3duoMPWpnvi
IT65Td6J2FdIAEC3z4CmrDR1lDXtFxOdC3qEqo6jDBrTUMo2NZECyemEPDT+1uaD/BlSaTMn9xT6
V2JRM5v3P2iPdaHmEy/9iir8JCQ8brGYjfs5ziaI7acupJwVhUbKJT/EmCOC/2oGWNuH4lf+B9/M
yerHCXhWJ9HG1Mq9W+0Roevx+A1DFvVFv259uhn+hKNRCKWfAI1t+jh4FLZhBnV8XbPTdtvpPGGL
bk8W/OL+jWpo1b0XcPGZG2n8q1tZhIYXaL5dVaMub6RnKo388LxG38mbcj9icmUbaNo0C2NmyUYP
5ZUcUhk4C3sZ2zgk+G5fKaE2lzQet8+HRCBB01GpznLgFxuyyaa+T5erY+CwOT7NDKgLwrOJ6Ohg
oKUStqHemwf64am2dDTZSYUfyfJfWyl0yPx3aZVS4FVqAoXoRqVKHreKA8YFVz2EJ/ImzKD8M9hG
lgi8yWh5MyPUaya/M9M3gRH7BjnL/odtidoXBJwT8M3RGiBQ/lNDYT2S+XhqZMhj3rHDmDtSQYmF
dybOZ0njINABPordBdGOEhYhTntpxtgsTRq7+Nd9Iww4CUXWHuUeqtGLvpsprmPgxFXgHnsRlPUI
fTz9zQixcEpbDLe0Ey4P1H1riNUiWRKFF3ZosVtqefPe8tn78itKpQ5ZNmtIp9+12bTKGjPZhzve
AzyEuyIYwKmCDnViL0AYQh2pQR7OjRf5CMXVF2DLrQ96Ae/BfDIQpKOd22onRbP+/2sWnMZ6NM6c
y/WxfNE2+jeG7ZTvvLDFR8Ax1ixfeTy5sgnr9376C71jwNYdHsWVH/5KmrXE1RjQ9SxxcbAFrumD
uBYd5Nt/8YZFFzmqqTSupiWGOaM0F4+G/aNGDEV/P2wJWOe/1I359cv8qCUA+cQhF53Tuq6nCxYF
zath0QYMkw76BLmEQH7nBZUO13w3I0zYScQqQBDwVfxx1IUeGN1rID8XDYe3GsQqHHpDHFYzpTfP
d3i5yCm6lnZ1p4jzluAAQ9AZpge1qKq351hzEkBWn0sWEcmaPeBC8heJwIENy4/J8we3C+OfXHGn
1a1vFPfg6DATrpjDk+2EkqZ/lKbdtf9eL/6fInjofC4rdQ+XdJKKJPB4bVIkd6A83lMI3jJfV1+r
/7tKZ0tZvksrfg2z/oOIAcwR25CZ1W0m5rFmS9Rjd93BTBQJxQKp4HzkgsCSjhRKoGolPYTJkpsk
BQhLhUZJAiwzRf7XHtFs1KhY1+plmOVkGXtYPUuZhj016unBWyZoGVUtWsa1fS6+4RyUjqrzwyww
IZKq9iiKWh9x4BUDvcXe0tenqfFn32XkMytm9wxXYHVrUx2BBTdb7pCMM2sGjUyHPgBs6b0H/d3R
JHT94aw+p1OjY0Lc4FM7s96BkBA2AC2ZAzHb1/kZidtK3PySW0x0m7j2T44DcbTSXKBDNPX4qPeV
TNCGMnRrOsz7uLASYNJavF9poGdUMrmJbt1H/8mt+GGkOp8bLHcwk47HcbtW5PhQ03e3xVEsYqhd
pgKv0Z7JWdJ/Nu7M84KTYqvfnTt5BvvwPROgpNqk64slCGd87vo49ttHzq4yus+remI7/NDLbwkQ
cxt1bHjiUqxKDXnMaOrhlvkW89xvcHSs33xf73oVs4cQk2LkPm7eEkNeP78Q2m6cNvKmb4pS+umM
uHFi9Xd0nnnjwOKdizFJG6rHk6/vxigOfoOOINiATUNKzrS+eRJ1todenBc/ntWc0Ae1dlYcOetA
RVLIYQa+8HfwjEOrn6ij1a5oIzZ3WaX7MfPwkjU7Y9Tilt+2T0xu2YZfeG65En8NMN1OfGBHuzJp
+GdK228ob7kUVb9CcZEGcrMWvRVnFkB19PF9gqclou5BAM+a9V60LTlYaKZm8iLfgb9Y2IuYNmJj
8LwuB82s9Tu85FRmKi7fumJbqfBFB0A/WGPLowy4u5sBajyDKKfQIvu6nWGv4LoOd0QrwT1hzwIl
vsx+3yCPmlHMJNVGzLXopKaMy0cCkOMttGya/xsqZ8qNBQ819ajzknbeXF3KgCFvw9s1g840Y+cg
bp6SHRL53U72EP1KEPbLND1sfV/BWSHyDPjKhweVoH1h6/nTii1erruVtEPBefnaeV9ToiLUNjkw
k+5uz/NwfZ0V9W1zNZutgjcrAWVfwt4jUQz/6q3JJl9va7UGI4wpwDryA3ibM4MwuIyWbXfxVhgh
Dy82p2LZvkO6dLxOtijtigQRE0j/wSDl6V8Vjz0xDI//oVUVEK+eko+hzgWfj6V9qf/6qiC++Ca3
TUaQ1sbBJHmGszFZ6DN+jY+F12mtTNUJvTD4ulJ9T4iHzaN/j7RBoOPsOzg82oZ2Fdy6cvnuuHm+
L3NM2WTPhgSreM6HVmwuh0BNgyp+t8azegJMAU/IZOXDWa2dyQOJHFXE2lJUQQNNe76fLu8v6JxU
iRBERbLb1twQySWIIFGoVGug+L5OvWyGh1G2ZFJSB9+U95/7YSuzPWGQz8iQGQCxiiRkwdl1m9FZ
7ZBqHgNYH47fuPB4lWXuvToti6/fcWMwI3gpswZD83eRSRvQZMckZKG9PSq0CWkmdPu14uvc3pvh
ZbElgFVtGNw9yqk7lKO3c2jMC/0haxuelQCsZRk8m7wwqZTaTWcwCTkh9RLCvECLXZt5LiYCmJ2v
9sp4oetyfuX/vQ6KWWfTQZQ2IKyuZZTUqbEjDFFPCdUwjZ3FD3Ey0Pnq3mt3I6Goat7XA5kEXv1W
CWmVajcLn7Zaan+juahZttheauVQm1cFm+fTpKdOve1MyOIiCyHnMs0O5k7I7+fMt7Fa4BJrt/rK
Hh65JWNPaBnWxUGFk8RXttHHlJF7ygbVLua5pD8es64ODAVKQUYO+MC1GERp6yP87zHnhWojhyYK
SniC9l99O//sjzE4ejGXjbL1WdSY/QOHuVvvMU8a4yCHM9V3ww0HjfH+v9fErHjOjgHVHeALunMs
/qBoPnPAC+VzRp1TJz/R85QCwmdgqVNhgYA136tkksRlIJSx3RlC+qzTgShIx4dNObwS1fjn1kSs
BK+mDUXHj5j/AuUPb+Oz4aaRvltjdGV5nEfi3Yb/mcFrqc5ICBMzxmvORhQz1+ax3eKqBcAWO3Ma
9tDJSwf41saTqdn+9ZQE4/cfPpt9FYuDhVSrdar+rxpL592Ew4XO7AzNieE8qEymAkCPHrGLRWv4
YETm5nQq+evZEDPGleUoZjl6qiXR7z1IMJuz0TLucukX3pPZB0rGsPVMJMF5m0oWpbE+qleO1KDY
1CkrZi4K4pd+xAuAEnK/HMgGhVv/VKVMVVjt0y+nSsC10RGKS0+m8rIFP1qpEBkOsIKnl4SHy/gl
1icmO9oAfwkBeCFCSOsL9DaAoKluU0EU+Jo25hvIky6JS5c/eLx1/pxczucJCmuHbIHHtuAZclhV
T6QJVLS7sB4ZLXARLymkk23inf0vQrhR8ooXwuoW/8BITKbw9AHckavTynk43T9xO60dr8J38gF4
8Pc3akSAAe9vAhIQTm4Hp64uv411Ttk6D4ZjtKrtWvTdg41gyFdcO/N4HmKob9KQi054YsRnl2qr
DGkEyz9CwOP3t0WujSFC1YVS7LWn4qz47YpPC2JBkdqKFK7/w3OUx54lBTQuux+AIB+CJ5qcBToz
mJIjpZAeb8sfMHw1dw315HwCmIp3l9HvJCJrpfNIW3ljI3F9/S2dbApOoMvgrPua5Uq7jwok2Us9
Mh5/SoxI6zDBJqyF3W6Ddxfi0W40LGuLnZ4HeUohBL/9R9Ko+szd1k9HrXphYC+zROlkbSrOwn7C
e24jzb0ezeXgZqYlatSkipEd4B4wqJL65YUgXifrlN92OaPHnMew+o6tmnA82vNwW5tppt1oV/hI
C3Toai506rvWHCGRVelTT4lccA9TveU/34fm0YaEeCPtOS8wNwb7TTjOdSZtyNGHw60Z2VbdNilL
0+5G99kZMtzn0v1J2mrMNXdccn6wxUlyQfmS9DcXmYGfPDAp8xwB4aVuKKSOTvq84gK+ehJJskMZ
EFvA2/ZNFU6G36LArw9d55N6J33wEcH+os0bV4N9Lv7JD0vxhhAb7D28jx3BZd8QiXhs9edcruwQ
EZzKMgxQbazqdwiDxy2iMtOI96mG2bEF81mjCJJF6s2jzB/+2YPgWyl6lBQnrPmNV929IfLewVGP
6/tAFbhfNDHPKweenscgBiM792NzC0vXdPdBlTfGF5lsDUdi4BxbkyjsBGlUgyvu/jh9hscUl78m
ynUtXKn0z7mA4/iylXL4ldL4/Lyfbk7keNQg/frflMJ9yib8TBAUVk3MvLH5HeNrwF4+Zf1nir3F
e8snh54ZlXniWN8mTLA7M/21aQBz7bVeOID1LaszR7OJruj1CpoR5ItlfPzC3D+qu24yldA1fEyb
+m+4fp+SyE4ppHfSRxCDOyBO2CGL5DaodaG8wddf901qjFcSjE4FDFfaa5DOLpb1JIVzifd6PMfR
ST+xYvhcXbzsrNI2Edt3yAXblQ7huIkEBCV8bBKl/XeECBpRE1FSt8jpk15NU4J2UXCtzJzLo0Pa
5hjwo/IdRIGQgSr9CSmibU9oUevBLXwymVuZWWqk8/pFp2FGDrZQS8vjTIEGYx1mTkyaNTUnzsAL
Nigg5tLVmO6J4d0VrN3NF0aOuQMs3R0gqXKVCvFBqYwnNvMZYmKjTKtSc42+sZvZsROIJZQFxvEg
pHuqyKDlZpZprsKcx/B867I/6nTII2cHHJhxQLpY80EzekDeOf3HzPiO7NLUq2EM57oaJ7FLCXhW
Gi+6d3p2yej09fi3IAN7TQQBIzgjfq6L9l3aJRfiwtj4bWLEMQuUZfFwbg5Vzg94gM9AE2l25/qS
eN0QQuDOFp6INyic4gf1J0QidbCGZcdYU/b2YCh3p+KI3KMIVlgi2/9WBVDYUtg+T8MgcTSsTvIB
xusLJqvBQFHrJeArY2/FIIfu2k6/lC/c2LIGWZZyFdvrnjxzRzTP/p9yi7GbGlKclKIMUVwCieWj
Mh+OujEwQm11vGprsJTx1wq+STQ6rr15VCL/P6Ib+vWiMCAOKpvTzFuquVfHqAwDC4psvv1idws7
G2yEt5s+HNQTD+Ag0AFjCRqeeGEp97GFYPlje0JyeW7TGwpuyHbcya+xKGATsFrpEB3H1EB45pJu
MctNlw5k1LH7tAkLygvZ0s9HUSxNHDzrYTI8AhwQOytxucGR7/ph2W42llboOxgp3zNkPArdzjnB
hi/WmrWpQLo7VXRrxNPaBYcVR9lo/1d8h7r8vr9AHSvPOle9uKT2tSiahecRGMg649KqSDEoG7Vg
mqWT23dYwQW0WycVOiMqiwZljddyIX7B8pg5tBf0NDDAa1niZuLTinwXzsgcQraKXZryA65v3bQo
XVQwwfVYRlyEtvpaclPBVK5pyAZGF47eqfftRcE+z03fm7s/nWztADWDCAc2DfbkdNzYpFPHvJ4w
52YKS1w2nTtVinKmmJyoODGBvm0j0S1hvrFuNd9iAGlo48SdGDBOo6gVhBKYaL15UbhgCg/6bveB
89MzZFRGRlYT09wFKsS5dHAetEMlGT0a4kwjng5YAkrYR/fTq4b6RE7HbpfrDtoxXUtgJGzL2V1l
gf3eHTavkQ2I7aQ0c4r9XjS1WL+ng0mi3iRrJ0Mb1unzcKmiFRmcRva6Ey4+84lA/SDB2prK60yk
OmWCtpiM3ECPKHcTjGFnvGE5NFd3S6vpnqH9PuvpAdBP6nOUdHMIafEEBoOXzoB3ADKs3Mee2fNw
3DFLWwuAMfT86bKX6Y+Vw869E+UJG7fv9INO5mE61GBsYy9eRKkgY9AO3dVzMnUFVDGHbz2ctPBL
52F5Hoq0GzVL5D5L3t4PirEMzuPt2mlt9FJ0vpnEC4oXcO8ilcEQfOjIhGICxvTkAn2yCX5Rlc9l
vOCnIKeUVKYHYAwJt9LYRxHYI2eNYbJxUri9Gd5dMrYbgJ7hTzfJo1WBXMrwLaDP5VjLtEpVAJ+0
jdXn7sL0TgqSQr2dszYXuJf+HMSSpY0rGm7tuGX5Bi0HCDPd3SsfO3E9WgGOD7n4gFfuuBi6Nkhh
+37Pt1wLd0sLyyhOgc8cnvFn6t1AApQFVSas+Zsw3Q2q0ZgQGJpmOrJzej6iGVEF6XiqEOj6iJUm
DhsQjlCxIE92LS7GmXyVna10a0UHtiMwO3rTL3t4kIRqt7A+3vpDWK2Ephshp65wrMgF2/QMm/7H
vNEXB4/3YTR9xn9vy9dl8KUpNHZbp9a4sHP9BTGOS05zJhUhzzfyAtcocqz9GaWgaeu8sj4/N9DN
3hr3zqgkPNG/ZqyWi7yKiKvZDURqfeEGMXGMobyBEgxipyXUMIAZKK061mm4cphAsAbt4JPoDN4i
gy96F3K1GridqCebJE9XNuvSa8EMwis1H6JOlgbCkt+H2/63/CFb13eMpcDToyowPD7VrNc+bLqO
RAdJ5pMthyd+uQGwsZU7llTnXXo41RY8gHiLW8GpwBUX+CVt8THWLJYhmgQJmXG+lb3GnTZzKNuH
RLDfntNGH7or23xDWq6kLv4XPkbLJXrwlbwS62CTd39XUdoydwhyYV16I1oUkdBNnN7z3bfXxTe8
nvj7vBKEuqQ3lgP4qXs6UF0jYL7q7eAI9tPnkvup9MJoLJHpxApY8TLNu7TnBNT3GAIIo20mGgLi
e2SCMXDqi14v3yci1TMH5m4Kix9yUcXou4IzJdRmJcTCQeV+IcV2Eo67jvvCRVkHr5viyYuLYOSm
OaBQxD/iA82+fAkcSZa0oL9412seCbMT79AE/B/0uipvIAeIA6zpfcDlvZmiUcjoZ5t5jxnVE3Y1
pPVKqMTlGJtiaj3Dw1xvPGIhefNnFg60b4oso38JODYlFF4/+tPJxoOwo/KCn4exQMWmCG0ELzEK
YAnKpWGGtSYRdQ4EDdjEwC8Dz9wqzs3fKW7VW22ewgDR/zgZSG4SnVcxtCbSMl3zDddbwdE1cHam
5hRq2zTjDGp1WGkjmyGQzWLzsmWWrwbAxu0oM639x7P1oZihBZ0FrjaDQLJx5W8iogPaQBGkKm2T
GOKmI4kBWDlemi15AtITilJyzGKno7AR6M1dvO1rB29KdNanIoD22lM3ULWrRG5LrSh9hUUkLBzY
AFaj3pvHJXOSgW8Ws8PrQ6D4RpHCcA0sseLZfe79GRUhkAsPdJXVRGPsv2xOSSPzS1hWxW6RJ1g5
xO+/8YptM9xD90PvjLuBiRBMzFIkLq/IevUxwEL5gJpN8QOihmlGLZNYqYNOKPPZSG+DGEmeftj1
BeJ20IzODBZaZW+SxAi3MYUQp5c6mIobn+iAAtRGBuIEOgkwkcm9JxhRwL3wWUNMY3ZdwE9QSu7n
C7xpnLJGJ4k6M+FQ4Pl+JSjmqZ8VAhBeRq72eOq+sYJG0OvB9d4vi3Czg1Z0MseWfvTQK6YhRsco
VUD3p0XFUwA1fwO28EidhzobodHB13xWDjHgYX69htQ7Ur4HnMHyxf3yd0WFpXe6WZaloYQtWO95
gGSr2x9xKr8uLH7MUgogyQhG0vJsCnowPbx5D9cUi1enVp3for26bfmdkkYIrmgLquztpej51Ogu
kzSY80r3AtbEAiXH02QYeacQ78yFlwu+tO6vU3/vb5+iXA301BOOsbHquTII8EY/pYSoR3ox/chA
So7Tno2budUKKM8iF14J74mVKubWk27HzADFNqBiHvHQ2YxyYY5sCIDHjp37pKIXqqpEd3Mp9aR2
ju4N1H5ks/DBgQJtukIq3fSQKtV9OfJb264smVoAI85iTCflWVZ5rgZ7pX3bL8/sJt+qiSeE2HaG
tyiqHFmnv9P/MbRsmsDhpD40/ZO6wmlAG0FAhLBrpaLWVMkMAWXS4srxYyLdfkvK3yiqup+47wwV
kESmutx9q8R0dEVbObknMUzq7cou+05kG/xO3H61rFZzR4rNLaA+3xlLD5RPvPwBRWxGr9l/9Ime
lWqxpvjaIseCjyos2yuE1a210zQiQv99qZDjE/1UczEss+DxrgalstvDmvdSPAbj0PrC1P0GiBCa
oM9fILpOSTpclBE4MafLPUZlkZTBOvRk7CrD5g8E3yX5SNdSuFt6Jjj3HHQKVdkrJufxAkLhXO9f
ix2fVmbRAGzxA9Z6UL4CTRPsrvbCN6cJo2Ur5NmmDFJsQVgPhipVkl4Ur2u0Sn1B5cH+qUm+YWZx
ghUuIZHj5fhUUbD6Jm4ZWPrja8RjWFTWqqO0cEudET6n4JK058vt55ePmIG8W4L9AS1GZMHkkx+t
bFM38/qab1LYVrmN0Ebt2BNRFchX3w43+JA1m0WNfHgYeB426oGOVFVw5y8c/s93MiFlYe2BvQKM
cREn4ldSB8a7ayAlTzTnO+yYSZ6tuqtVk0aQnyUEfECHRE3qRwhOBG0GWRQQpCy4egM47F7yetzW
xdF2vu2GTpAeHouwhivLVNkx9jEAza+8q0Lc/YHIkP2I1xapX0V78MT1lrBuE9Nmg7LZwARvdQOu
QXBqScUPXxTYVue2ygkYap2F8R/wGCb5AM/yaVcqjM+b3gxgnJCyBoE3Wfgza04E4MeOKg70535B
G8Ox4g7yPrm/u0J+0AAbIXkm23MCWFxP2B3szOnMKKTkeNp65aOQN7xODrfTZE8Uq8opchVYAw5R
54QY2iOwFU/gSD/Aep5eif4evuYYcSBomJgQVJfWW4BgTnKiYSsdw0QiNadd3y9sYOv+NtjkTDne
oIfoZojA3dmBT/mCZu9sYeawQaZUlv/m1IwkGwT+hnWjCUPDbVLQPbdGqH4l61AS7kG+i5MddFYV
pu3H31jGmkwI9Et1rtOn9dxE5xWnNbnNQ7LcMJ9TNlRaCkUOJEC1lBUODqw9yk322VSUg7Nrpi3e
ofE8lClOslDUHpMZ3YCdCfp8hS1y+2HnsckhWa5oVBi5FNeDYLwOp7jiF6b3gLasnmSY2KlrIEa+
XsU9jc9woEb2sangzhu26ZcootZtQ++ss1y0EqmjH8ddVD5Zy2l1AewfUHwpXo117EBL+hrox/PI
2IxdodT2A/Umvf8qFWzn5rARy/05jvbkEI3oKEYzJIrJX8PIyjBu4Rv0BaXPMKrNFdkN3mdWqAo9
cXpuAFeTMNQmyIfgCza4toRqswjLNizbU83veYeQo1LAr0S+ustNhjSsewvtxMdqDQ/LJqQJeKpB
m/vrOujNCWcXB7Gh6QHoSkjci+ZWBuS6wzl5RHsp0Tg9puSBCzKrotljxAiKKe6RNYEfsfEsEvmh
VRUgxiE0DBpNDwkY8nd41vXCj2XL5BfH1ifcIfxRbXY10/8sOCpEBRf0wwh1kAJbfO9RqbUgmBZQ
zBozqUK7tOPmmBodc6TB6A8g3B+Kbh7uN5mi3JOFGqXlTk2uWOUnFvj9/Cj5KebOOiznjABCZJ7o
ZxnWvw3xfTGrF6oojxqBVTYh5rkQb5XWiNlsIIs/X+uTvwAwHn2kRDfIcHHS/vDzcu51MGpddFgr
GbtoEydgBLsZvbe/0bL3zwE5/4XrG5eQjM7j9rbR08fwBa+/KH2kCrJ1pw8m3bc14Tb553kO2MC3
RfTEV9chS1YP5cBuTJeGqMEyHVPIcHkttKz/rcOIDu81E5iR2M2H9yrMrjL3DUeaotcQCyj/bUSJ
nvxPSmSLd1Oe2QYAI0Yue4slx+MOYg1AheqmwwdCuCxakMshpCwxbK2h4xC+svewcJrPXiSjJD0A
m3Q5LCtTauwe4S24f8umD1LnslL8FAy024SqkugKslU1oEbnlIVNSMr/iB3AesWe5PvxfWO8w+LL
flYvWNAzm0bu1Rivf/LyyRSBGwAcxMlbeV1oUEYys2vGGp5Lan0wF9e4AwhFtUlCFwsr85KDnY/N
9SyOgC+WmH8nOpH52sFcexFYVRM/OiYe3QLh3KAsSxeVRPovQ1g6L0GKvEB9P/DpNL0dtPfX15jR
gZLyyx3YBu8UmGPzmJArF/CqPY6Ib5x+ABYS8XODiVj5VlyKMomAfKClYUM2LG0XIQle+Ct9xj0w
dSaOwPvtfmcNziMXP1nv7hQlozZNmO0XbNJX9saPBySQFvAUgJIyOEdGOYs/441z1ObtMv1qWrEh
TWzH41zLbE4JDTz+SXYi37ZutrVvIGEjm7oN9jWa2wPmLYnoMeD0lvhhulyiZHj842pXbzxNl+n0
U1VahVc97b/5t1PssQ771Dl/uF0vv0aqbJvJAugMOosmOx17WEi4LGnTJOYPXK3Kxbd0FqzpOGT5
BqzwLdWxpKIBC2E+DA9yVwLKzVtr5wIFSsHoA92LWKtD+5d3g/qjDQ/PY704cQeqni8u6DLBe5yv
lOZZLro3cwM2NYe/fSY54KNYVGthwH5sYS5BrbiRnx1QMrw/Y7AYVzoZh0Nah8WLffqpn7VOia00
HpT/wHWm/zFFmCBG1JvqrI2r/vnHPYpGlcEABwhohJOCkJZ2NMD4AiSK2woeP2juH2q8S2EbZMId
Qy9I+sCTW4BwA3a1huA70GraoCj4jvXCeH5+1UsM/jSnFoaC2L0w+MJuLQ30/eoZvjSJKUEzuG7E
7yGurPbV0VBhttGJZlx1T4YRS2ciUO43Nh2e3umPG8N6N1/T5PYy95rsLj+htYS1XvOx4bTrSQHq
9uzblOVFrf7ruj3R1VsnkaCweCYKB1Diph+Z6hRW1MVjuDPdM8cVXjcLNuuPyHqaLJmWfd0zGpND
HEMMKbjZkQF4d/g5XQ4+Rnk64Dt0MA++mkCR9cYZLfGzM1OB7rwAmHAvmZcYULBeIgYEednGaPML
fMY5Ttu8b2DKfH5UR/gPTee9pGjBT+lNABpwTeHnQLF6DuQdOE1w2zIFNMAk1lDwpruWFJhsNdyj
sCcSorC1uEnMglgg1qCs/7LCqBLgX28Rx76+F9bgCeb/TfNXnxUulMAJY5+BlPi4RItIBAaXyXyE
BSIordMxRYxOJFhNkuOF1S2Aea0iyW3LPtWyc3Vp1vblwn99zXtBvZUNfKhJDkgYJbefPFKfz8mP
W+WDw1psly0OlZMVnsmtBa7OSCNxS29/5mqSOpRkXHRAzYCywAdQHsN+AORooMnWxLTLi4dJLl4d
+MElaE7/iP4EkTdyZDyv+F8QelQidac+jicxIPuemMzv1x1cHY0BESC8jOl1V3jT3Gqi5K9a7DgD
Dcp3xwQAUY501r4idqAbgzFC+vRm3quSK9z1tCFxF1K7Om+L/sKtcwb5d5PKRr1TVWdLhcT6deQL
YsIpkYYuE53BpmR+kxrbrDSOdBSNZVJpfFlaGYuZjVARXYtfbZxNr3s134Xj9Oc+V1/yl1cSnhvd
rX5kGe2q+p7Jq/9P1z7troGSkx7ss00QSZ8ZP3FLcMiSPI0x6lbPpJt3p9fyorK/X0ek6la7q2Sc
0sBn1Z+nHv7MB86sPOXJaWOZlvTisInc0R4FbhcU+0eKyRdmtLpNFuYzHoMP9uk7iq5IVQq5xRuZ
n+PllGtSYImlKWynt5oS/tLuK+Vl75HKMZZIHJ4XhHCb4ralzn/LkEqdvfINkMwL5MGCGyUS4YB9
a37bEEH2+cZbXS53tJFKSHmuZ2ykOH8IPmRIuAbrPDDLkH48O8oBF5tCNI27ZJwQidFlBSYGoKZh
V/kSLGEBP2MDV/fYfOPqQ49uDvr7ivhdYiRakVC73G5G38Z8lIjPkRW4PavokFxc4s/PUNHwNvnJ
gP9CuxisUbWXENcyENWlWLgxqdQvJdDYIoakeWdvJn/HLdg2znBIZvVOirIVoOt/6Sy4StrRr0OQ
2TRneXqruEjV4D2Y9/pDWr6X3l+MxJcWTgkxa8CYCR87+OccqAV/TjvEHZ0RePKPevEpa/gYZzH3
BvYynNscJHraRR/lo8eDiqcC9MC37sPcXwfiWcVjcPY1xbsgivyZrt38mb8mITsPn9h1B/87g3cS
K2gMiH5zbmqMxR4VHpd+OvP4lmj8mYy8H8YzN6JtwppdBsSWymCF78jCLHh7F0kExoaSfMu1U0qG
luBCWdnCkqout6zmwcyJe0lkVDAbY9dtVVDIED/wyMFEWsLDSXmSQf9HkfgpgQ+eUNNipafsMXQX
o1PYQpM2kiJZEooRV0UMY0ln5fb49tNDMyT4HY+O8KTNPaS904o5aXTQIMMOiBY9ymN5SJ4JUNYV
tgBNj8EQvL+0tCL03sDGFatIh4tOOxIrA4Hiu2OFUUUzhc/rARCo3k3zjDA7V8DRa6LxnOPQdQkh
sSjivzMpl4oSgfBw+WSj2LvR9PWLne7Jc6NOS4N9UwmCctsab8niNWFTJdTo1dEU9SZr9xTB8n7A
53agQT387ptKYbxpEYcLIdYDa0KxnkwdMK60zgAGjcQw9KELIms3jbqddG/DDvWtDvkIFp0SRZ6T
beDmWDty+dLlLni12UJKtb49YaNnZVyaqeyEMn6yjl7qWxmGFdiGad1rpq9uJ9CP8F4xQcMkZ8Kh
xubUR8LAQyfmIjNmtqn8tacfMgFkS1MJBAF/e1U4/JGry9ctGm5DKkXyKIXP6N0YSQ46FRGPs+4d
Cd/W5LZoJHlCkOIidntTnFBoYf3mvcUkW29Xk847IXxVaxL1WpuJAjWm9NWJOmRmKciocXGdw0dO
sn3N2ZHJgYXovgju8PqLrJJP/+rignrUlDDGWH/+PjuHQ4tDTwn9QvgdzWMHXs5KgK1BGzqGoHFr
Lnm4XSYEZexFKIpR4319sseJQmgCjy9oUqeJYdKMrABh4yBNqKsb+WXdGGmi1UKB/ltaVrCiMeoL
i2HyMRTHOgCXDXmGL84jYWQwkaXCZALZc8jHphS+rrcK4lk0FOMzpOb/RWEUop3qeCoSXg/n+jmb
b5EA6GcRQTzyuPXlIdHBYTkXfNY8UOUfJlorO4pVXCsJryUgcqX5ABZw/aOioE6iAzFiuidcSHd0
DdQzMfyGYf9O+2LtWrkepcBQ3EXyS9xuR4sjcZE+gWWbVc3PW+1NXfmm7xe/uvs7pzsldMj28i16
Ftmpg4D9MQIZfL885EcsWvLAJFtXW99cy/4ALF+Qu1AIZOHfTWPMlQ3AxPV9Wf8ItFaNLR/UheZB
0oQLuRIOe//tqD2HYTx052Z8tsSJ6YIJpRO4EThbb9Eb6AJJMNIgYzhN8uvn9SmRj0rFSyu0cgCj
LeV1s0Ey0i59OY1HNLo87Kjy9LVyjLk1NTSEvEBjpRMWwqi7lDb+KUzLUxk6VDY305FEv909gujT
mHahM46RlFzIJGR7+5FifVaUBkq875p0MvN34OwzEOzyfDFMDJEJQi+DrKFBi1EAeowOa7hMydsj
5Qt4cPUBgDX+ByamnAxQLtbM/rJCJXW0PiKycOf6a4XNh/aOgAFsFrtBAIHQ5Klgy4J4nze+EvkA
LNwVNb2CMU0yv0ISsaKRel/uBmIQMWNgp4NKL8dd0vSMe4OokSC82S0bdclqgh5mnWkttVqJZ8rk
P82IhGT/K0q7ZrZFdzi5ZlIfYMdqJw104QRjI+x0XzOPRRBz+4rzQALNo8q72+qboEW7Wy8QnSgZ
YvPURZgC/BNgkDkMl+AA3yefHsGrRhD+j2UvQIE8OYDiBywcwWoV8pF5Ei9US7C6urecGceupb71
MbRagNhhTFfoauXQnKAtNqMcZlVpbYRh4b39Q5Zm0kCh811rD/30V0vqgJ4RBbXifLN7kF0qBy9H
va1iLG8NoAH07+0yA1Opi23z94Zy0qJWBLcgPif1VxcONvCHtsHnxcgHxTcxAIxRIuSsFB6e2ahT
fSqVRzezVF83oT9HvFJ/M2nPL5EhbvE9A5N1ACE6ABebQGdu9r4I3shopu+yHzo8OYmg9S9GSHBb
G/MWbtt5KBVHAwnsim8xnZRYFn9dc458r+KLZBPFw1L5bD9SQpwLtBbBgVNIRq3qz2sjzGAjkDMk
X2ofTf9YIZtbBKmuxbYQ40yFqCEQBSJVYgL/FL5dc+tPkAqbO76j9G6TkQAwbWUzpWR3aIEiCv1L
u1whzmvgsbx9X3W14K7GvdId8mL0fyEb6a8at/m5HYQ9PSmV5d7p84jccrfQg/SainKjSxou+pkO
2IWdwrm9qZfl+REIuGEuet/DH6WTIbBTHO4orLQVpyBzBgpLKosMyl+VijZWoijnWxeU0a2Ztvr5
j/yUL1SG0MIF0/2e+ZJHbxZiXn6Ocgd0wJuPHBrPW9f0AWcYoLiw/OoUP95NgnPnO4GV8y2mGEw1
5rYAUC6nXJ1jMijJdnvg4h2ZSZTC0Nk6P+hZNY7C2cSYFv6jy4MedsILbL6PM32zkwL78n2WvBYc
ZO1GpLJfXH0SBT3fxK7VWwdNNww6Wt/ZK1O7h2ZQGL3lTuctjrh4VbmB09FqgM07NN5Psgrj/Cal
zK9xWcGzokStjU1L9s7noPEUGssGQ/3nKk/uG75p7jVQ4D+u4buZK2U2mALr5PBtFVuTtx26cLZq
dN/bJ4uqQmI7d51+Fa6G67NXekPwwEZ1P7IdNaVQYW6hlg03y8wKnJTUCIYbHJTJ6/dxJW86l8lz
968UdW/Ft2Acr8CoYNEl1rtYppHH6FafrD5+IU44d8AGowIahZhI72SSE8YATppdHPPoxXAlZK0i
QYYUFnTIyw76z/R5GV1evXHB1ZRPpP9DElHsTx8UNN1QCLYatRWMI+UQf/z9BUpnYZduh3GRGnK/
ITJaPG9UIZwTHXth0chiTsCVEZIgeNB4kMXGEQp/YQ8DPUfR+TUy/ukl5e1yU1DxZOs+8EV9EMau
SOie6QWCN634LoYNyU8c7GulgGWyDg3EYtBd19sLn2Cqh5VcqCFAOsBLuzmZv+vuUKVP5ho4Ih1m
nOnn63jc6zCcepU4oW6lpABORUQ4XvyEHRbbfcwvkQ+byukQ4hUBtcdec3ap1AR1G06Zzq0tR6aa
zMUNzSudmYl6UoG7n6xaghnJAWqOo17XwicTLzVv0XJhfJ8Igssv4XSr+d9ZE72zyOJmcaIHN6HO
5BaoI6Y5yuyqubwQTmUBRzO5WzKxQgqTMvZYjj4Dw+eXGnJDfM4Z4wd3sCwYuJAOaqEP14RzZh6I
hSCo7Q9i3yLz0KHK/Jkfdme3wmv7siNFqciEvUWFxH/5oc55bsU3SkAEkcOMIeDgOzVrVnW91khu
uBW97m84CtYSuElBzw4sgRiCM4KtaajdyJFXU4otfCi12Sm7HgUPH34yAtlyWq3cymi9WPfZxW4L
4bGDtIJPsI0EUkXMLLdQXJga1mTeJZVxl4zjAj4fw8Sy68wGg/kjy8oh0knb4vxI229fntY3snJX
HWjlUCHeG0jce/RdmLwVPOOGYk7utehJ/ndREOxg0z99dmMWmLTPxoQ8hKkVu0cK22nMzyReZROE
y77nZBKC0P5fLu4lFZ/UamzYG/bb74WwdE9dWv8t2rPHihmeFa5pjD3bKg+FerKWUeRbK/RUBdPi
zsa9yt1Us9Fk8ysjzxR0r0Ce/rGmCLzW+59UUIh/6vLIKlD40iCBYXBCtHft9P7PGmZq1EjFWTaH
3SdnOuviiyoumvJVnP/BnutZykWhbOqXnAAVM5z5sVTgdrStFVFhUB9FW5zz3NNBhWaMIl/f4C7r
2OTXHaMAKzbiV2ZVEZE7a22WG3fGltZ/5nHErsody+HCU0zKXlevyckZQ2vQCKot6NGQxD0QuFB7
Hy+ekIrmb1VahboknilaG1IeHvTH6fBH8RgKZKqmUJeCz27hAEQaI2LZfmOVqRgQnHFdTa7waG7L
AYZN//+IRKu4WKnJi+7Xr70PIjTXq8gTjkZ73LmTwXaLQ1Iy+yQ1c67Ixjswd/UCfsPcOouqWbNO
nh7GDV2OjhJvKhfdUw4E9trbNdXoMRPTqgOasxw6UmE4GoLpbNRsiMFdklHtpMPnOTDYjEi1r1e6
QkL1qVTkLCdhzsO5ROnNF7l9N9eThvNgk9r3Q/u/oEjcfRxC4XUnuvBopGX+jDOiLRdmorZVtd76
LUnnCSHguYvYweVClAoluPEHYoTvhf6T0vYOaDFSwe33w0VDiJV5yIDn9kn/CzCP62dXebrF/OQv
dx9BEDIoceDXb3wLOub6kzPrrU9m+S3NIKHr4WD5yjfX50NL/qjvtQcX0jvbaT1vsXQcPFM4Arjt
2Yv97R6JyGcBOjU7fJT5ZmIfG8Qa5+UnsIzDg35+LPGslIJ7FMzfcEXwXUG+7QX37Tkin1eOOsSo
Z7fgYRElxh5DySpaMFOodJCddhih5GqV4EoTPAKEkwwAzMj3iz6iKwlkz1yKtHK5Pa6nbzaDc24S
dSMtrLiTr1YZeSWzZn0vv6dV6qA0ccifOWmBp2JiULR4IouR+exuxkSr6HsgCoFfEB/D9gNHJxGF
wtsIgJHUGZXkNIB4ytkR/hqnN62S36/lzp1dm3FFYSslh7hKg8RBxTSKVCjl15MsvvsFD7141PPK
QnfC9/a4f4Jiu4yVAZGttu6PDDjHGlHjWaKEY89nmVy2NnGwPrXjPQzSBy74MpsvKgpK9CUxnWnG
We4sTmvcQQPmfm8fCKF+tXunlWQntdM+aNepW4AlWcrmUUuijsqQwG08tuey3G6K2Nx2YQs16fI9
b3d6OKArO0CdWYJWEjygM0PP/+s5mymiWLnnXuXJ+pb30SDygS5UlOt1ufCoKvHReJlRpP1/CSok
54vf/cSKkVvJ0bNP8b155big/FghjI1QXjZDuHy6UViR+pF20FX/iDu1Uc4udGkj53b0ytSVCYKs
EOf5U4wLFCKTZBthVxCFaVsYjK5adLoieTIITxCIZDK6YLFnf5TIcyd+qRfQbB31+RYF6B0lYMwF
1Uc2SQWsMR7X15fi92Euyw4VXjYGVsiyRpytN53s3Vvr7Q2oswg5aNbs3HjzsxwosSGsI0ZtchYr
4xW9xTHs/O8UZf+Xi4rvEHVKUE4clTNzq5dBvtf07kHWI8o2DC9i9cB929gyjtu2ztGCWI6v9yNk
GUdOpM46hKsDQS0BT/EHhN9aNu4Y2K/XMSNLYgtBtCt5soKDALHKoHHdRg44nZ2bow02impsIvML
YChKD3k+jF0Co2lHA4DMIkhcTBzP9pmVz/pxI3oJGaqwuLTSOd87Fbg7W2R8ErGsFlrt/WrwjzPI
BESF4VMl2x+R4hsX4k1O6Shj/FCxkSRbwy4gBfb4o6utkuqLdbPqF5B833sXNeeC/o2kfHQZMbF4
urvTkr1U4PmMC13tKZk9Q9xinYn3nV1CLgicntD2WgLQZlAsyLTyU9R4ErxpgeikUi/+saPum+LM
9qe6VMj4PDIoNnAqegqYjNIia3uKM2MENYrrPE3e6r2BaiUyIxfDpMrIDJtpM0Q5Bc1YE9/Mw71R
JUZb5Eb14cIrw0ANZdNfBkJbYQEDk/IGkLCQsXv7sJCsV4/iAQWeNqd5aDB5lmlu0hBLYcHMvEe4
nZn0XKN+CS+uD3mnDaaJbzWi7putnl2pFoeYzYWS+aegRbtNfbWr8zCc7Ht0UtcOxey2rewkYCJc
bqPlGHSqpmfzeCxgNrU0Q/KiSu5BIG04oNN2nM2KPcgas/f8+8e/snukFXe4Z5ohIFIrGcyXNeGc
epzetM/8CRBCTS6mt1ttZJ8WUnUcFfSpKYV/Wy5ihBui/Jjz+KEnvVweEPng6raF1eeO+V2K7j97
4B2IuazZYNVKKCBijCn72Z1YmuoJKAqNEffJDB9W1IwrEfX8ug+3ppaT8z/qUtit3XNGnj+5tnTS
s2yav+AotWo1IvkUqrbGcF+PQ2SduPIePyCoGJnsJEQBKJoaIm29rlHg1XcZrg3kH5CFq6uA0Mip
AMreYspvShnPiALfQLo8Spp67hm7WnKfyhsgvukH7fr1ygZ88Gq1DQLbM6LQNvrJtloaEfEYGjDe
JPFTkdFUREBW+UaRHHX/YpVBopm6SSWMschWkduXNG9tSiH9hR4eQxIE/Ofr0QqOPaKFvDZtBAsF
lprouhpRlK/RKDA/vz4Y18xdP2me9t0rhV0Pifu5Qtci3zyONtXbwLaINVTN78PL1dtDliYViNfA
lPIC9ut5ixbn+Du+okpQxiH+ChdThziXJvIuUXEsGvggJfkspVN1wk5ilAHEPEv7L1EzvRkPSIFc
Xk7WFodbqP/lhJOOk8PoAXHvo3wQgHua0bbvvE4b3KVhzlZ/9rLfracLq+Hl948IIysrLMiq8eej
0AFHAfIDEakIjSfC1m8bQGlS1ct++z0yA0cQHsaucQ5GAY6wQwKPW/YfNdkb0rOEj3fYlwurmD8/
ZFBLxpWlAFkVYI2bVmo14Jqz0idOQ4rt53zN3h+QQXefxtb4PKnXv6cWcd0u0OtETr4v5PIi7XdN
uxOL2g8wod1/q52CxRCZXk1fA9wVo4qA+pRFN+zlrjbekwDVXBfbSsK56+usgK0hPzlC0xAhBiPl
KSJRrkSPCq7KJwgi3zobUWeKI6FHmGGW0w0Dcpf6OcaXiaTIaHZroGWj8YmUKL/0SYgPwqJz3mH+
yWhE5nMIRr0b1sanPDWQX2j+UG4XEhWZvcM7TLyqWTxY0KSJVZL9mokucaRp1iKdbD7suEBDf9ug
xDxWICIw+Ce2HGsWKh5gwOZU8UYta6daz+EtmZgV22MJmM5ToGCpXThcqaX2iOqxIbQX7cwUeHbv
HSvAgTX7i6+mZQF/01vhgAwToU7gRvUGmCYtUpqc/YvEzKh6J1hraSs6gWSsNwKq3wlrEdrnhEA6
zuFyt2KF0AFWwrgzWxNqUheuvuanJiAcDLGcb10uQEsvnhTTBoeQA4WFmPSNXTjyEybOs0tEbqpB
5/9Qi+0uevAH2tlAg3eAdDMzEMZzpr/9VjFtVBkxytZJnYm4du2VY8tXVti9JmB7lRl5AqLlQHp8
TLrtRpAMWIe+Aw3SYvxsoeRODHlC6RW6svb6lzcqyY79c7BDBQj/SW0WOZGCHedv2vv/mKQUVOyO
gBojPdwAAxs4DkNK7KlBFngdGePQcZBUrs5FTKh9DhWArFDLI1mq27yuasFahex7rRrZ+8Ev+PwP
KTKbeu650y/ooBBSvFPs3T+UEYLOBCJCdLdUD9UOYsnDWXVQcyFSabqll0el7oXYlqvsaU8sNeLT
A3sa+VSlkiZ6lieHHRxo8XRGLoERm9IWZ9V/DiFXI6fDZoSIlhEe0EgD33r7vMzPBfziizJoOGBr
KhuHTPJeNOXm97YQI+m/ZalGGkeKKrMx9pJ07KdnaM8KnwvYeDqmRGh4uj0mpCNqDlTSLBykCMKM
dVtUk/ZNZwW2Xdv8ZVLytLCaElLEeDInLnmwZ10rKhJ4ysj54GsIdZaFthnrL+IpqWPZuqOY6z1Q
AMohOSjIr11gVa/NiszNBAGdCZjM9k15lVlTUx1I+ituf3G1tJgO6C+276lRDO1f18+y66bbFzzl
H1UNrgyw5YKSFMixcgZpORZKncZCUpjEMvt9ySGjmUbjB1+tlqicXy3+LG6tTLiqPD6nnuRDsGCq
GHzEyXEZGQoU2nubIGqv+TG+8abnjrSE/7o1Kr3ImXyMbYLgUYWz+pgcoMWs9beC2yWzPwsy9PLC
RM4if3OnNAhL0QKyLEZsz2Q79ZX7Yy1NjMN+VC4AhPqNowmh6sUlvRspSKVPYsC9YPvJtCqf0CC1
P5Gy7D5MCtYlniFGU8Jb6EdSDxK8PrTkqEimjCE4umRC3+KPAkJiG+5Ly0aKMVonu2nhFrSFbAqt
LJxV+aI1z9QzNSUlT8RHVLoNhone0MVR+kGJvPj4q5FvQkh+qtLTFe15DPCC5M0Zwwi8/S8Vsiel
7DSlitWlKq3l0DBGh/px7WCT7Pr0eMTl+1l/LOuoEFwpcst7S9se06cBPfv61nV5tAoi0Pgxj67X
hUeik7Eux2fKzqYyuHeanZrcjJVE0VWa+k2E2I7rS2kGEtsq+y0+zACjm00Gw8VoDKZGLuQXkaPG
nX8agimM/vNlwS8bIrikfatmFqjtnkzcQuQSEBs9R9bdhnPDLs/IwSS7yCe2indDI3LND73mh/qL
vlXOkoZ+MJX/BDWJKvkLJyTh6ef3BhJY9r9nCbrZdks6UCRMrycB/sORXrZH8oKIdgKmr09Ex7q/
4raHnMF3g73iKZwXXn3Zld1NN7HtqI8K648Jr1eKcUqPuKTBxy2YRUBvrJb1f6BXstIaVTzvAGYy
HMSDGuP22pcfCSnREt7c0M/N8VZuF+4eMwSzgx9r/CQEoHLRzCnWliqpcA7z2o/Sp7u6elohj4vH
4Xgk8oreGjBRxh+8kXpJzvOsdLhHTp/xL5jBHo/pEw1CLuf/uvBjzSXGBfRtS19veIb5lVu+iDSD
hn9w1nDXXrSYQqHaQqJledfhqbnGsXZ6qBtRTDkwgr/g7ARHBtBQ36xupaYEOBiiZxeUKptbZYRr
wmShKKBDnx3Oi+8sbjCNsERgRWJIDxu4afCew5DMvlkECp3JCjhBmzfYDso08al3mTX+G+bysiaU
fGkgb6nQaELFbZBO6PqhJiDNVDmbNJGCweS21mSMG59F9E/7za4eSImTEIFnvtqnN1iYVB/rfAZZ
UOjjVVvqtIZRvAzRA6M9FpYx3d9UwFySSQuQ4cKjfId+20KPZsXHAb5z4S4W2Lrtf4TKjGMPaVTX
Jcq9ABpyYkLhUPr/LQCJl5Cp3L7T/iKmmzZaNrnAq8jcpy1j8pXrpcCoo+pvoNcr22xn7+3ZO9BX
YwJRTtQsK90ghrO8CZ/sLH6NmSKpE5uxOMaLW7IoZtODyjRpdKF03pdWBPvRk+NSCUr1lRNWEh2r
5mqY7sYhOzyl3lGM9Cs4LQAnKQhHHYQd5s3GQPQ3GYPlpACYi5b8704CtJyIg9w8YFI0I2xIqATR
eFU5RVzTL1dA+oBYWcV5Tq1YylpxK0XTERMhNyzJBZu7cmQvLzCpDuD7Kv291EczIyEm2oFcWNrI
j84jw93kczs4feMTJvp0ARE/M66LJeWS5DGycOuIqcm3Lx8+h+CSeICWVJjayxiiXx44zJ5haolO
0AJcBK8fE7ORjtVkz5SYOda7OgcKb+NO4vFhVx8W1vYQhl+C4HVaPLbAxPe2FbF2Go2Ngjly/59l
nc1izqxWlPHKu4sZFAaMczKNwi+SyNfVeTGsROX6BIXDomWCZpemIXIpKM2JsNpubnTpC9PWqSQl
MVS6jtRa3J9IQUBHxcOlGp/qo+CynSIY9J4rx5K/E1WX6paFku4sdZVx/0VAGiNHdZ9zEYe+shVR
ih4vUFm3tLoPhC35UbXs8gEdtWQ9WMTQ5DKPlUC4cvtE+elUD2Gq9U8NFZlISaznXtrLifkfoOwH
CdlxJKz8fdfNY0YlERLGYArG+AzUGNyYR1RdGd5tPUBCrJxaepxv8cDY5Z4c9Szn+Y3mFGi/Vwgl
8qi4XL54DqPKwmP++SP6nOd21ChcWGYCk/M6UHRurRnsoMacWcRyUouISpujYnNEJ98D7XrIxp7b
6P4KcbWpMSYtKrt5ERMdzuvwPq4K/TAovTuxAiwuWV4Rw+lWKJX9S89OGRtQ/caljcOlEMXBMYeZ
z6XJPb1pQuDC/4uQVEsA3HBegu5gBnWGl7j2XFEAvewVvlPSTttKRRAEfKXMfMV0/Q33H2Fad//W
OfjfNCLiOTl/3lQF+ISVR7PUTFH8XZvn4M+lMjrJSgoIP+5yWnpHyDlu2Bhoxc4Ab6wAKpfTDmro
h+FGs07xrKsujasb5f0zujf/IRBd5LG4OOwxNUgJPFxEyhv7akk0BvtQMZIS3IZXC289eIKrbph7
R1dj3ot7nijdIZZ8ZlJFfbzhW2FbTX/8nGFl8SPtFG9oepS+mtSkVH+5kqnyBRrZV8IDkMlrlXNh
a1e93GamXqmUo/XyzMUMyr8qvKhxQKUrPPpFIL0KJhKzx7hS1JLLILk6CbUhV60mQIwu0H7de6ef
UzPKcyafUWAWdbP+i2FJPyQmxKn3UpErIZUTL0F1hmBFVVaH6Qsa3fXaXbpmWFsqHJfL0Y+0LHtL
DdPTk2cbrwwxfiUMqItC75tNm/0oom7h5r7GQFhRq1/2r7C9psnTBbn1U5YavIPaYqXH1ZngMRTt
Kzyw0J2nWd9z6ttzKsEb0ymrMefHzuzRPsGHaoZYlo1ivaprF75GJRFO4ANbjZnw8CKGfhlNM+d4
7iLM0qPPmJ85PqPjy+NL6aga23Tnsyyzo72Tko1qYDC3Z4UiAErq6SO2oTP/YC9B9LPmOHvJUOWv
mjcd87X//zMfO6PbDRPtsL9h8A7x0xbBp9PGZVfQ6Nw5qfpZt2z9BjUJCoXwU0dx8HWwnGT4YEXx
RCOxX+5wizmHlCdLN5NUIAZdrabSeZHgPceT1ut+SlCKx2j3YQfk8zkwG58wRCrRNz8Hvurh1get
P39AWRdCNg96Hpie1lO29A8kc7mbFC2LVE9U9hJab/sWM0Ef+U29/kPARiWT1rVKC9U1dQWAPnTC
9j+EscnFy4sw+vr/LfZsA5EkwQsYh2f5ikZln5m9skSv1sm5Rlhjj5Tr/Mmx12T43rlhSX14t/6m
Y99UjcXy8BsEJ5tf5B87Uw56YLQuIB09nMmXugu4xKILkpegTD12rzHbsdhpwOkR9TkclEIwPDow
3Yh2VioSad4rmg//JCVR9mxxrHm/6xoYDOiJEY22D4z9PLYOYbFCnudR0EsSKkQZwckE0EFZXfSv
fB3iDGPnh9WS4zaTj3YxAlbAeTe2OEezbMUfFdhSl9EJncI0xZaHIDzYhdB6USBy4OHzTFvXVm2e
dntH8XVLtJKOXrc5nT1uj2rmuXcaFWhsMO68FR+RiRkEfSsAYn3g/oqaqA66j2HkIUoDyehRWFSf
rCaxp7j/v2qor5tEiX+YbktGqP5EECwlLex2y7bmxW9Z4llSvnfK6ZdC4TT3vYcheY1EtzYViLjR
I0j/F0/sQzgOjoPfCEAGn3tY0dKFFcSx64Jtz6X0ZGyTXM7IUG/l8li0B/1lVgDbZBFE8hRvSvEY
9VujSm+b9drnqEyyp/Dy39BbIfvivsZAX8k3+NOTqBbSDQ52+ei9SmMprErhSqIDh5rwS8OqBeNd
PWJQ/22GBaCWBe7S+2G7TiD7NQrCO9LoEvYmefbwz++/b1SH0vhAFVOKND4ne85RGXUAjLnt2Gjv
nDhoE+OjV0RFaQjwJls+D6X0XspbXak5c60TD4MuJZj4SXa3hv8oA3E/OHEjGUGUC0G9yQfIQ+Yc
D9dybLIvjb8I6AdOcS2tMl8WEITvq/KCI38duSNSpI556F1r+tDqy926cjrZdbqX8pX2tiEp4kRn
dqysfqjxYft/DxSmtSmmn/V+OV60KCu90G3BhQC66z6OQAu+LFbIpGPnaeCfjOP64EW5IGas8eAc
R8NMPjDpP3Hre++P+jybYgKL+kEcLyUW9EH5/3vHtkrEokN57jcYzuXAhx+Dj+mAx8hQSpy/iM64
/D1R1CxZRR+eLE5UQKdSzRZLg92TAUuc8joBL2OySG1f4tYTldYR9VzkQ0Mv6MteODgIAHLHrZY7
odBvdhYU1te8J7DB73eleYjHr9MkXkohFdqM6ZeA6jXyUZIlQWcIjuEBiuGkPjERYBC84mrti3NP
YzJqV8pIxbwHr/3HmtbLSh5/iLAE8e8xu6fZHeIsfsJQmIJt8JrjOjXIQeNHFSPB7O+9YXo6jFZf
rclNfxa2sCAHN04Ocb3V4KDbL5mmcntcD26ZGubUs4amzPQzdjbQLzB87foCVwITTIog9F+/aOwO
vvM+K5fMzMJ7TFTkJeUhNMfOAIuEdaaHhB3+ag9z9c08CuYZ8gMNzZsFKTos76H9Uip6YbVnLc71
boiK6TunMksEikqAwNzvEP70udL7assLcnNVssPOaGpRfQyCSH0RJnNwPY0hjD7Rdx2J6Jy3E16V
jO1HE8Dhfw0+3I3n1eeNI7vKWh7+GwyiF9an5g8o6tXZHol73AlDmrk905QEaG1CHcS23F8rnYVM
bgxajhVq3wj7EqA/Jrs8pi0nfJwvuoLfYouLF5A55XcvDxTy2tOMUhy5RlRyAllwmfnh4+GOzKbe
C6VhH3ESlQf8f4W5PPkeY1pjGWkpKWhdKn5zGB3/X803pyK4WQXGgVHkuPf/5bUkn8/Y3IhluDfr
PI8Jc+C8eP4HwLw7/HPVt35yFhPgcggHBnCHwWi3eM8vYlN95hcxt05XkbxntJVsaf/+LYNhASaI
zSkSl8wkxPDhPcRdEFiKj6H72zDgVhIOBnAwxX+JIGueADCgeAg1UnnhB2BA14MVZ7I3IcjV9Heh
QsAqpNJAOEVentzy6bZ8Yva+UbIoJfN0SOO00jZubYUET9Egom9bNjOj8O0fDquG3ul3wwfaF3VY
9E7Mo0mmMdD3slI81FpWMW3osjRtn+i9UfHOi1Yn6YdLtMpCyB1qncxriE38h20drLMHiPXIJpVw
ZcHhI9uFJjASeI5uTlwIkDEsRQJcrcLATrZ079mSBwa/SfgYzU7n4nj21z4J8rChcuJUzeJEUQR9
2ZEDw00a2cMHXCtEY+LegMtlVhm9TMYe61eSZC/UU0PkkVSjEQ7Pk8B9+6PsULpGbtJa/mwW3dr/
qQ4xqqW/oow+Q4txXKrsxuXkZeW1B/xsejW9n/YGbZa+oOZektGkCmCVXL2VJ1y9kh5E/6vge3P/
+7ogF8mv+wfAQA1JPIhlA5TvQBVXoftAQcqobHe2lUy4JNv5mINW6THdd3Hg+qrX60qdNTNvAOdL
+e4HALuTx4tqD1tqjLtw5nxr1vLOOlKlsB1wpX4q3typeJlkH1+LfxqfYipo/pR5ZFdIxE/XWYPi
2xlC1UUBrrSDQ+718/utPR7bXRtQyWfYR9xYRNsxI4NM/NniBM8w3QVeWnKcfJgiBCPf53xzGUNA
FVmdDeXCeQ0YSgmhxCCMkr4bRpgJSqT64/eg8t3DSHdu2bIGEpBJIeXVeI8824uk0GIeGXBddXUa
cKI/Ni3M126A3QC9bOTn9A0ukbcisP/I73K2QAP9SnwY4WDyj7g7D4/37raHAjKt9+weDXv8AxGB
nNVNgYTKN9uC7UYx9K1V2gSRExbHr695UAjFsBn7MpNHGovIyswdEeARlyUUibSmpNXIaCAZz7DX
7YLN+hGO6GvzwiN1t3d1JUdXXvC7cDXvDJhapCiDASdMC6sFVdzy0NKga/uW8qyzriozBey/SSW7
wyJcdfoToDrGaP3w554y6UvTZgP85K8fJ7gcJ48cN3qUa4ioBVCzdyKt6D+towePlXJrDsXWcfQY
EOOtf5p38emcjVImyU2PaEoQEe7WzBVspUbd7t2O3lYBeCUfdvxbKznkKlea6NHu9neeMyvrcvcA
HmThV8WWe1KY6GpXvwGxaF88KbLizTWTUPjGMCS5SPD518FMP01KjjZW3pOa6myQeZJ6R8XakFpv
JajO9M0QjHmngiwvxu00vSOCo/tn6kvRNaKnJiPbXBF3McstAtsNrjgvEPrpAkqO0vI0nUScVfyh
GnNhwhnwrplT29skQp8CnRXVBgXWSLphabOPIgn8r1GwKH9fiWq7ue37RI9FAOkF3QvFwqfp6zhI
4cSBhwTKqsX6zafa+Ll3gR8dHqHPQYUt29M1KawNJoyllKGbzV935eEcPrdDjwatBFvqyTXT7ooO
0MkEIXm6HIEXONfPfL6w313YKUCHya/nzqU5QNdD8RFaMWouLgdrEIgTGq6GvV8UNmI956ST+TVI
eMR2MWxSu8nVPhk7ucf2B1bekkv9kE9bczXO0jygvaV5xMTd2Yl1ol36YK0X8ck4ftNGzKxcAmiu
ZznWjYAt2V2wM3GEM7SI+wGQv41oqZkH0MgssZ6Dj6DvGtmITg/3/oBa6e/T4/d654ucpdM4qeOk
Aw3ufS031tVia5kH3WZ/na6SfmmOJ2/H+ZwJvFGSc/h544fNfQq/yW2P5RHxpfg2Ym71gYndIe79
yGJhx8JcNcN+5GA4/OxGG9sbYhO3iKjVV8QDslRdWX8bdHdfGNtK0okiLs8CVuo41kNLLdm9eY79
75DhAeLcbiWLz2w+DEutWvmp1ZUwaHGQxi/7BEwrPHozzLSTfox9pXH0IpnvuV9NCQvui+FBTG5y
EKH0cLKXmNsqqYSIDiDq20sJi+aSoR6ajubHpBKLHLko7yC7nF70Yh/2tvfT1vGp1Q7fi4+e58Fa
4ho3udDyArSTDLvawDbGV30Bd7ZFDzwxAZGmvuaCZIUCkTigQGDY1DpHTCwgtEpwGezNsHVudXs/
bn7IyQKLos/JpBdNIQ8xgWIBppGwYA2lBOaPG5rOiiK1uuOyalNudNRR8Ope56xdz706HGCuPeFR
KNCed3O+6vKzRf8O8aP3tqMH9rZprVMTSprdrwRS3cjbbxiGJ/29pNGiWiy4+jT81DJcfdWAAycn
BFPBTeB5lSl37ipNyh+6RtdNmxAHK5Ctn9sI7PeCfUMfSfe7idmkrK1G08zCR4weT89sYCyCR30O
cUOo4K44+gzh/o3zdzjHO/MRb2JVYPOPO+kuu0J66xnpQrIwx5buQ/TsEkUmGg2n/bmJ1dF3nxcH
BcVv8zxrZ6vkORfnTGXEW9wHobDNRaypZqm3gg3aWsfOW3hBwJ8j7ckxhvoFvuTD+PnY480Czcc2
oEHCbnTh4GpQaZrhV5vlVnlLBk1NAlp3aBXuxNsucHwj1ErY5Pnnmp4OfKNR1rwk7fVrAY2C+nqR
rkaHK/H32AwA9tkI0dYtkjef3VExWPOq7RL8DaPyzQ3N2atvKzPl362wsj950rtlzPOTwabtizwm
L+haK5NI4pav9yUpKbZ+8UFCTVI3DxQ22tSVdLVbb40whNSQfclToZuUPXjqqHfE7MYENgRzUcyI
NfZ8MvVEvdDuim7OCCQ1ahBvBkjajxGLlDrrATEsfnlC1lqe+zhH4zd+LchJ0Dbd8xm8VOlqWAOg
a9NLAG3VJqGFYtZ/ZXC898pGdaYS9Sn0ff8TigBXwd4SSUpneiGB9HoDwuZGY0TZSRiGxGr7gKLU
l9OKO731J/jWKiKNSM/d1jIN9VbJnSCwS/FiB+kZaeXYNUGQgEcVCS8XrfdOGDXYoLWXMq2sv/Ol
d+ii8ZCTqhPkbdTGHv1AgevTxeI0gTpy9FblT9dMyQQp3BGq1M5thwG8SWAevYj6SQGPFvz706kn
0YLJmMLDHDwGFgOTeD/AcCU5rLwvGpsK0mOE1kSesMm9yAqz0G+nHu1/hMqxkWD+ZaUcv3LNRo2D
+L8YXErYt++KklQKyHtHxRVzq4ra8wkJWtTOFIwgUbjjkqtaMd6OBgq19VXlYJwintvpsebiklqC
lNqsp0rdlrniJmJRNAd5MpQ+yUilznYfqsYrwKohMKPuBaLqeRAG/+MgTVqn2b55VoxJqewqSTeK
s7NUnzIRHqTQnHq2iWUiISNO/9BOtCs55Gly6ui+tnAlVr4jXe5hCMmk4pfKfSlqH3EM+aDM5+ZK
pZr9YoWj3dNeMJBnKWLPaAfpYiLgwYAavaH5xkAgawYPlJH/e/tyNsll+JZkX+7m0PNqSennrs73
QIfQip6oMVcBtlHQ8ux1rE9Qew5jbIJTdyGPTM5oAZ3D+hbe7YzIxGtHktXZGHOlaq84OGH6otks
pBTuaQDnAEK8nH4eEmSJIoGS1x04ztwzKbGAfRkY6BkN2f+dt1ZYyawgybjQ4tc9S6eFXp1tNcAl
ijakRY9NLkaPhNpLJcbDCe2vCB9AwRehxKvjCRVevZgxDrDTV9saHsjvl/gL8MagCmt7eiyh0lWT
rncTcCBzKNPDcCghtXffxf4rY7/t8Z0wDNHRqxL4B5tWJl/93lqoEsH5EiEh0ecHKSC/7m0FTjpq
6cLmcOuAKfk+RblCxLqYzbpSppEfWw22BLRw8Ul6bXsCofMcGGTQclQds9C5E2lA2l1T7tNS94C6
KXqh4jjiYmlwleAspzJQDs8e/EtxAzvqlh03QelErOPRwTNWAWJhkKmFc7PbCpWO4kkqhxkwGrAH
UAbPKoL8Jja99JOULSzEJ7XI5iYsGG9ifUWssS+QFiCsZEhzissoKDQRPw8JMd9gSGCuuOyueMac
N22ThfDdNGIaSnEBUtzDRo3pSZzVu5OMziVyFUrA5OTxUE+OkdW4YuB5OqaRrNtGpI4t3lIxBew8
lpNEG07VhX4uXlyGUjp+c7QWxVvkF5GfEB86R+3mHdAiLwa1XHPa3CbqkmJpKFyECFUFf9aIXHjV
Us6RLeg3FOPF2RiaLS1bivVln5HHjlSpTzcdGXYkUdaeiIU3DDRK3w7D0gEpedyKUIG/+PXkRwMw
9uifKxcHXOf10hxY3n3BV3uhp6/yByxHgdBvI50ZVbpK7/nwooM/Eizk4kDapcJsXNR0thJ6QtBy
sBP5K+qRHSn5wqTvFv9CZGRhed2tnNdnU4Z5CPoycRek1mthemD4Nbm8NCG1eFgUwr5A+eWsl1et
Sr7hmNnq/MiWEHFKcJS3IbQgy5AZNdXUtMy2ts23YNvlRkRiuoOKAWcTKZlfdhtmHgY9V7oxsPKP
26zy1x0Asi9fEnx/w3nY4LeqaF/mruWLj9JRETjSES104bIf3fuQSr1kXZyrz/MlDgBWJ7yPnO4d
KqBNKrES+CgwrJsADwNoKFnBy1f0nNHbizOCNH80915llg1j3+5MxVRu9rjikbVviDSIa4uvZ94A
57S5EzSsVjtRX2/V/2PsUrcNfd/gNwq/VZtDjPF1FOrOtPnHybhP8axDzurEBxsBpzv8W4h5/yIP
4DlYBViaO7TJT1WMoihSInlfjFjIqNWUKfDvNIM3qqruxggszkOmURHm+7N54s17BDf6XqY7ZmFz
g+eUcZIA9QdVkInPeHHt9PuXFObkNa/nbpxzFj4jNLrIB4I8IEPqzOrLTVOhzAposvM3p5U+bgIM
aa/gVYUX4f2e3k4njoKreAZ+i1d9lP17KHvLehwSPs8nFFK/UOv56pyMFspkX6hZpQUOWcWoZdM4
nQXeJ+O6NiqMOpK286HgN1M+pomiyfaFhkPGKbaCoZKQdp1PyJ/O9MnBd+d+VDV3IGNhLguXaRXL
J6D4ip/0chsXgTqYSolUVpBYbEtoth2iVrdESqqmMbHIiM23nichkYVzKYocgyNStt2SbWhOkoAG
KAFtEOdn1wbuDhiXZl8FAbVUSN33UuING5rLaAILRqXvKCcIxgRHMIxUX9buZXTkCw1hryJ+Knj5
GEkugRHPt5K+N9wasFK3G07R+CyYs1wV8MsXELl1ruqMA9a0fXtQlN0Ta6IgWna3732RCYRcDrzA
cF8bTYlCnFKDIrzKNnotAtTazALHPmRedHDf/LFru8j1XHeWWYSbDy0eE3WhZHtCfGwnWrqj2vLr
Ngq6lIcbbh/VHzqTkXi+1K5GlK2bkj7Z/Zx3cuNbiD0OZB/H2vN3WXzrOjkGV82A6vbc2WBpOI4E
QaIwXVUIRppy9o/PPxvniTyMPfaAiUEYzGu0XdLDmZbPywtG+PcVFcafqwlxCDY8qsQVy79fo60H
Ri82Ifl0TK2EQM2n5nwaAUFAIMVedBldHkAQoEpr0I5Z3Y7DCzXzeDQZ7sojB/jZEoWfwiuyMKpj
PppQ6cF4L7MayjkWRA2f84Jw2JIPmpleB/0sU3rTdJYCRTNTByLGFRjjY5HaRc0Cl38O+lsJpgkr
WBx+Km2vvn1LV8f5q/o/+ePEaCcBvb/afLlAgzloex0YqrKVTOvlSXQaA6UUTUdyb1jsVRu3+Mze
prg6hqdpxTJRQ8N/WTtmggvBFhS+ECpqdTHB1kj1pQUNIxFpe6E2LEyKFYOEmCoD5k1caXyLXk4w
vaYijyRmuF5U+eqQiAR9wfW0VF7Hi/M3XRFa8D/B2V9+xLYaG4F23clsK1G0XEqW/LwmjQjRiCzR
iLf4W6ho8UmDDgGaj6RLh88uwAjgpPl9OnH/ok/LDuQaKjV5RS91gXhk+8rLNcuJ2LyoUw3bClWZ
dUplU99bq9OH+ok7n09w76iB9YEsg7/boWjJpXHHqnPB15x4D9Yu/BsBA4TZMQx6VMLYEoG7LRgD
N653YQVEVFyAa9wXx/GiCZFF8gbq5GR8SSftJ1ZxgTNgCrF9RVkk4lv4j8MvqHZlJvgEXN8TMxev
N1+dFlIAOporwNNVLkCvXe+tuExz6Bk3RAbzgrAANRWopJyto/LGMBS2K7eH8tZMzEtoPH66TIJO
XGKm+od8DunniDdiPdKLtvusmVH7+VukkCCJN8Lu/ZP0EYQaqyvVSoXD8swNKxNxUgNKecURt0Bd
WzuPr+cbmZnhmRDTglJtMjGuY/FZWNxvPNYVkO+AwhPfVGvsQZaZfjX8V8Y4QL8lLk5o81lFvmQU
y+icRJxCIc8Ql1pt2UJEENpJ1D+TvHM2rehZZNOCSXvsBDPD90PWjWbIMlRaomIzwk0v3/WBp7oP
/mOkDi5U/EPgGktmUsaFOb1zed8Fuip2WnA6vvNq28BtyEjGZElxk5hs2dbsazKg1IJjRizbs5B3
aIFMSHxamt9Sa35hQXEKgWEhdFAeSb/h6E8q9+3PyjuTS9+zygcTVZhJdGZqIu5+hXeXUypJ98fS
lOeEgNCaapVupWYzd6bo/WHZ4KTuFzr43pV58LRsWjdxJYCNgMfNxgtlcnTKa94gLmvjOY19aQ5F
q+LjQKfRVA/C93Q2fuNW92/a6Zp0oW2nkfZRf2oaNhaj/pCmecYQTuTUH2zcDHaTz51qdfn9iM1l
pzbuRb6urzhuWp9sP8Uuhsvg9UYIwki2cJd+XVEFcwK/Fmjp7mMAs56SrButdUBnyDPMVt4SqdUq
uaVowlb6uqRBE7p8qLStZ+bTUAacFwfHVtUqk3jVwohfvchpVYzWptNa5OcK3GdE3Z9LvqdkQpwR
tZhV6twF9MU3pDc0bVuO5Gwro01R2ComaZ4vK/jjCVLyN69CPn1w/FjSKlv6QPNO68sBICEmHWU+
4FyCClDxsrQryqHVy4OMORsjf/HXl5rqXNHg1rxc0RhZ/euvg2LYnQEKTc4b866bFexh8rhwoJVJ
R3CnIoKqbnpvGfkFco7emyifEND5wTB6eojvKnAoKoy1bRcHMCPVbf6tS/GnfG0aYqnlX1FHvf1z
OSFBOxXPJfR6BO4hZotC2+MCjZqgb6L2pSMpucMWLkWLj9UD0qt6iR9DCOm8DrQdopnvsjvsms/D
ILibuxnkw08Y5iDKWtE6fpxOBIeVHBLWdhOpvKJi8V7WbOvWZS7wZPEE9ZTKrrT6cTLKMeBVODYa
zD2PrI0TIcjhPsPYv4JVwm/BoiWy/go4iHbYmsQSLoIe5jSGqo7KBynpDMXgn6Hn2sbSCXasNO57
hAk2F0YQcqP+pFCZK77XOhpJ/BOfhUGRLQVZf6SjaAk1cGJIFG3tYMdXhoQZd2PB8YkDs+/CSTpd
Ou+wDyRULLWnjpRNjUdWRHRXr7E+EVqCArjRGhN6zhsRzzWp7NazFFBSyV33eF12l6/gsnDpppLp
/a8P01PyyE6A8jDLx7PHBSp7JXPsYZUfUnWVxhWwOeSos3lUAYEpTvvccbd8D4ZXAa8SPedAo06P
dshJd/lKa13UF/HqpyOTp/LCk4B6bDuNOvyGxfy9kCc235EtuzurnKfLqhmjDHbXKj1/Zl72flam
jftZHxzNu8qIUbdltlzkylA0xTEDEZKvitaLq+NkGn6+wt3M3MTXtaSQhvwx11/V7qe+sxQx8aFI
JkpvnfVSZIx+eM/N1q6XeGhfyxlC8fWYeDRo5fC+cs0l2ddLFNvACz7Lt3fGynh8eJZkaChaxbnT
03JVNHctKMAOfom722zVBRoKBTgYWV85PiPGYzoL16zItedC2kWYb4Ktw/tg5zH0BNsJzSDc/MTs
K5oGzqn342OfLrRaN1IPdGXcZEUczFRdrYjl+xc2L3eNtlfK5LSiNaRRbRclmiSRaT3qjtCufDGd
MAbqAqhtBoR0EZj4xu0vihjrBw71Te5OoaMHpgQVrUGTf0ONgCpMbEgHUInxhQBVVlA9o3QSzdQJ
Q8xqWnlce87OB3otRxuHWVNib8ubetV2KYiOx45YWHH/IoigUC0/cEAhXurLeoQV+pyaJfGuUQFO
aUqNrxvspP78PiP6ey3q6B7RoLbvVpGeYzYyYASb4QO3CkLvchwL6bifkv+/e9J/CBEPlNdaU9RG
5G+uY8o3usEkxzPdqFzgjYD0VJMWGZRXLuVSEeS1T0rUrvzf/+lnsGfUgCqNzAeYATjhlAAsbNtF
ey1ZqDCxhzmUdcJTp5NoqTJsYUvSliUgf9sAR8cw/FswfPzSa4fFO/vEkUjSQr1R0rTslYuZMwpF
lEpPELzIZrabDgfidjjfOL43Lv6y6zx5m0tWYIo7oR9SoOCsMZ+DNOKTWYk711e+ODT11NC+Nw2T
17HbnImgkSx2DOX4ssvguWDWQ0QTSHM1mwy3CFofkeQb4CQ3GgS64Z82d8s8pyWx2QJPHRpH4tXA
VyjuZd6DzXoRX6QTtQgXEWkdG4Hv5zXqZmXJbGAi4QzSkDIei3DenW1enSlJjfu8NsuB6FcdVeRw
pALQXjziJoReuDnYo2FpQ9tveocZlUUrXI2/fA+UXCZcNcjVU/9sZCoMcScHxbCwUwpFFICpAxiO
8DjdKbyG0LnQ5LkJVkdsP+WZ1Sw7ZWLWrRk32iPpMODjUzsko8UzwguhTwxrTgTt2+G9AszH6R26
7ClgXsf/UutFBCkmnmUT5PA74qvy39HzCC9qZSz0kTgch8YtA+u8iCkF5CnMCrWATiZjlW4sMZDn
AmNhxmbBDNfh/NfKEwWM84nceR9gtX1rG0cYyqJdPshNA0NkOUuZbsCwmHyRjGs0pzKib0dvXQR5
mfeMcGl0Y3XNjQ41pJojJuC4WIVDum91Wgaq65oLAHI39v4n0YXsQMdldHo2i4FfZNPWd8560wXm
jGBGUgAFB1u10wsCdfkmvdVnoicDgbBeNvTKmKnICXvvdazW0W9OFvfAIMFQnQ44J52M2T/jnu02
u9Cu65orsSSv6hNCniZsItLUXmNcN1q22UBrOq1dU1SC8qc9KjOzSb7b5uUHLzFXX6VYN9dhpPT+
OUh1zW8rG9aP0CR3LuKjYzRIqhFbeVk7LKTcMcZjiZPommprNCiANAIR5UJo4groduznJ9MJoFlg
xAL4SWO5Bik9zCuAy9qZAE7Ei9lOCI6fTqwB9XyUoyeysbdQNw4UJeSHACWEn7LEeNhu0x5Zz443
ZDndDGG2Wtwz3uTZG4wjxq9j291b7PEiDGRRaST+bum7r8DvWV6L93CrizAq1AchFa/pU76rzETi
yhInZirTitps14Du3T+GTy3L9xmilzJ3sVO4//EJsBxfCfxwSGs6yn1wwvhL3IFCL/X6ToAkohbk
Ej0TJSeJLhu5V61FDWuQBXRHOZ1Jd1fNbfl7TECnWDjUKAU7QXJ9m+OR7zTzX+KqljENCZ4QNaJ8
sDlKFjCxFGglsPloHGcGaIQkCnI5Ku3illJGRWx+Ew4n4n+S7//beyKk/9N3pWx6mnVCHdjRD0b1
+K0xs1pNl0y2Y/0LmwFkp1LE76delpV0UzkdeginIYt+XXltYuofEGA7ond6XIS+TfhZYEl6KJcm
qLCniETp42nCpJWnIgy62jQ+rDVZ1yfjK2jtkagfx15RHuSF9zBknV/CZnqmI/RPeqH2D5c/ymAY
HC6WvcyZwWM7qEBdqPhL3ocyX1f6R3o31bs58Z9EF22/7bZjLn/70nHk3GMBhYlqAizAjSmzVTUk
oOSQ0VSeI9buz1pD3pCOdM0SJ/URBWcKmUM4pd8iYATJzDK9YHhEr6vcG8R5a/tJYMeccrC3wyFN
FoAe8VjUmqpuQyopnIkUFZNvMa0mbjWv4zZD4hHf+Y7aTo8EpjOsPwP/SlXD6OZ5oXuEz4bwPcbJ
d6oqZ+khCm5vwPemuDfU/x3RUZQLQHzJfzKHi7KSHXfox4aKLA5EOwdNKYptu3v0s2oYs5OGQBvP
ZEx/7dEQlNsFt4mrq9vMsKipo+x1++yGoW9+ykR7RmLB1KYyG/+DECaiekmAZoj4wj8k8GzAS+HY
W0N0MLeFDcheK/chzJi0hT7/od4PJMcw0rCvm/LQdFwwKnybZO/s3Yj2S9QwSC6nQCYmIty8v2LO
LszV0FhrWjcndOatXNdFl5J+FPdBiYpRLkjp0QdLU0ltHm9NehDpz74WoKlP+JPNvgaNT+fzjiQW
xu7rEP4ZHWs7QATOS0h6ZRa5W4dEUo9Q0H4JdtZxot+cXYROkuHqAwb1abB6fEEo7dT2m2eoVqdH
LxTEFT+o4Dwt9q49x4RCk4YGysRN8owe6qJujfqGK5BK1/DQ5jsFLkTFfTCR38zTHwVuD/hSAct1
/HVcTg3k0IAM7kAnLV5achOAEHZz7QBHj0j84NMNCfPwZZfUp0GIOfPpkRvMtyTs22mCKOc15dgK
YzOJx+DVR1cWsFSOJEY0XvwwNxiNMVEAs/3tb1wdnTVpRXe9W1zD5tNkq0e8Sm9GoOdlxSuLMIYo
KPTlBZBA+QcNDunbhcPE/9DzdO2VlaQ4OtmjAaUJGCF89QTv8j/yHpGurni2XMN2xBVs4eJlJrOw
+h9mault+QegbmK3u7DIgbIR0JuauXD4x+UDEqHNK7XpWdRJhL+mYmci/PqHQupMqFO6+jtFXDVh
z95U27t3oig/jNwiDU7CMgpKSK3tfaB3veLWejChzzPLVzXvqMD1onbdCX12vtTkQrl7zpb00+d7
WvbjtUusOzUbkgervrYknjCh3Yk8kv2bDQUKk6Kd8mulSEVxR/SLw9BHqjItvjS7BCFZYE+ixCyk
nbRhtVqxxaX2jUvY1eRNln1SrHzVDmIsmbW41x+HzudWiRWPRYOL4cF1ANTdO4dmCn0ncaCwmPcA
D32z+qqWY1ym4WR5KAesoQNvRQInR4sLxdz7sW0R6UN+NlDTq2qOrPCcP0Hu0dsEZeKClmnoUaDP
xsX9NW858gDrZTYxKkWYYrZ85m6DscSQjv1qGtL9rztnXyh2SROwxQSp3Inbh6ubx+npGHrCLS6L
sGuilXSRgUmWzdX4ICCHCRcX1xWkXBAh4yTCVGIykkbxpmQ2FeOyrEuCZY6Cyx7i3ihbzWbFoA50
lkYKzNFuiv0OKSxWLrzqwyozsRy2XEu35sUBY+Di/STsk1qM/O0wjX6x3RNLfFaBA5LLFhfebknc
Y8xkDp8E8lUWn2kUnogzLOt4Jo5eGg0J5eB3XxgC0z28NXTCOH+uaZQvfVsUS4t3HKe2p00NS+gI
PxWbUpRj5BYmnNcDh4EBlxCIE7i6n0lKR6XhWOV+0yoog5HxLBdFpn5hH4Op6QWPt1jdz0VcOxoF
JYUAeNDyqhpvgmaD2fEby5cX78+MoE8p5aNPQChkXpYQ/yMZMQdwviOCY447LiYZ6WCOWDNTCw7X
s8hn+ww+r1/retHPySDpS17gEv7VZ+U9RDwlUf3YfWdw1qidd027HdOGvj6z7j9b9v0aTk8vFOQy
K4i9L8i11z9jrTqaigD6LkuWFbeKBiNrr03vUJxxk024l1lM7NY0T8qmOoCsxq3c8b58oqPy1UP0
h6L/VPvY/f2jzva0YU+PYUf5l8BDPtwBRoz5qe1dUCJ9uwSJyRM6rL1O19bon3lsUfCDXUw2HFLj
lzYLdm18Hk52p0XizDjeIY/Dg5B/V1jIpxD9KFWkZ6y2uSGn9JQflKipNzezTU/6Do+Qldv7c2Sg
mi4CMs/10SsvxYn8cAc1EiBAvw6uemhUyWhUYkXSSUUZwFc/rtcyNHtTvdI+LRIzxFBaL348VmBU
M4ng90xx9lCuIy3f/X87Jj7LkfLFersqMYd5xxcT244lXJ6n6cZ8FXJKDdU/jOekhzq81VVMHMn2
2TvPyj775mwRTMqQQ+3Be+ZMWDbBG33FB6FWdZOiIHmmAJ1DBzkBGtTCkAPr+cvgiuNXarV+Cb37
p1J7RQMiC6rh9xyRm6rul+ngtaDuY1TR2CZ6gFvQ/4MO6IOaSBj0RGiCqt7Kx+EFF+EhBTYR8CGJ
rAnh+rLTzymwc11PEaMzp6kmqbMz4TaQ/i59MHOH/UTYbuzr81pSgNva2twF6nyG5403I2wVwlWk
TnEB3sPSdSN1RhTU0hauOB7NOoe1OLs8lQS481kSAiFhcesxcwo4RUFrdp4kpYJeLXeoZm77aOM8
1RgihhUu744FVugd15L+S48REdhOgr0n6iikenLHrNzBfdAR2wN+CAbjcjA5IY7m01H+5/G/zXAO
x1SZ8w05uQVlsbaO1m4M/hisna1NzKL5HRwfMPD7cRBoe9DMishh3VZm5FBlvW6YBm6WHY5QtVsJ
JGegsbAuSucv7BAHsZztS6WdUS1WC8B/i6sA0W9ARTxxuSbHhL4EvVUkLUry9Ze0uUQetlzHBwNS
h4KGo7tcL81r1/r8HcJQIhQFXp1O9BX4x5CybHzrXGNt0IOWGbWl18zqkzJi/rc8nOO0g9zrgRu6
8AUadMPcZMFXVwGBecNoptJbTqqltnqQiMuFwyZgiCDCEm+WkZTCfRji3SFq7RSZKEDssroDV6tR
MaGECLMD1N29AskUolvjPnvH2wucAT+IIEeJWIuJameXEXJk6rQyLFmyVL9YwhuR4VugkMvQnCjN
TV2ij9KZU4mp6fJUMJ82G+BCx5HckYVo2oJ3hp9gj+8ILd/IhzNWO7UUH0CzA7KQsl3G6u1Gv8iF
fbMniM9edEgsW8ci3NK0jfT3+dLb9YKsgBhECocXxQMu0FLRvhe9ODBPxzY3r3YS6CxkawH/uyxv
ILB1MDCX3UtXLzL7sqT+wBjiruSfb+pB+eWDztpS59MtgY5PsQdea1D3qaapbzkURKK9T/Gi3N9d
cdskEmBeT+kJ8iiWoICbbmghSg7O/3RWsRQsvs9ViKmS+8GzuJR7fHr6tBecVNuF9LePy8NcDA7O
m4CeFmiRviZQrPn5l7H75y+LjDBLn+32GSDEP2WjY9OiZ/1F9RFAUBtEeKbwFhJ8BZRMXKTmGdSv
ZjvjXKfzpfVwzFzNvtIj8Ot0SfzsE2I4p7F/oa2X4A5tp+6jwIrBOV2xRSXh8h8EM8+Swo18I67q
YS1ZlOvgSE4+YM/HJK8KTL7zhyVoSjmU/u8ZE7kLwYaH79DBhEcy0zmhtHCf3jLIHJTpxgo8hybw
5Th5LEsRYO6LfdGQ50Vbmfpxl9fUV7prIEgoAgFqJB0GRbXHHWvNqkc4Bil9XDwxAIWOBgLiuRfu
YC2YJRpzrgzKrl9s22kV1UwkKXF1vJemVINEZjnFKCZhrby/wEEBrPicBAm2YFHJwXdZFLTavIwE
zSmy/fBLfeSZW6lU1br7KKeaEHb81CgUvk4RMWIr2s/sqR4IArybTObG5jM/hw7jmEhpE8XUC7hs
uYS6kre2URRSEQioEDW8TF9tTjFBIhfgsJC+Xafx/IBd77VaTXf26wsvpdrlxyhvEhGO1X+llJFH
YBHSLZfqVz1przbjYfke4ZIVVENbUaZCkJ2tJj4vaV/zBWnqoMyobyTE2SGziODPAFrAFYMJB+DE
PtEMXPW5B/3uAlno/I4P8cFZXFlznACA0KNYc2tHqINaRr45gXo2rjvNZObq+yPuIFZUqoQ7tPyi
wvEFEDc4MGhqd4k25sdUiF7MVZbln/yYeRYEGGEjQV0kZUBwP7G4EcMHjVCgYdol0U4C+CkHFBU6
M7fUPG8yJlIZjC/e5cVEtAvhvSzmfLHqp5Z1jIHm6M9NlL+yA7u3+yppyop6JQiN/fm8MopufM4+
vg0WObp7+0W0T0Lu5ugknJ0nSpBuAUM71QwPXNCVHCkyg0XD9lclVCIvZGfOL7Al0Ueb51mVtsW3
gOUPOhshPtdcvk9hvmqU+thQDAtOd8rRPCXsgR4iA2/207RZMfWta4R+jRu6Ei/Xzrqn2xBQBD40
u0rYrMEKcRr7LbZa3qc/MR7qGg/27628dFAiuzXSG5eFJjilDUSokokiclWqNq0gX1M14Oz9mIhh
sGu7gqO2V/Neag6wyUro9iI9x+DnNDP3HDoPgoP5bPheEmA+sP6xi04IbRo51Uyd7VXYEavLppKW
B/IA+V6I+oj8dgaHgFRjGGjUAJtQdfIx/Ihw5nyLp/BrIS/eTMdmVn6EUQ9gzftBfFUi6NnKrnaG
6jUDnJ3AGAB3znp2DZOR14amidoSulRP6TI+I6q//pJWbBd2UJv7xcb+0ZDQS+MOgLfFsdQFfHj7
9m76Ty/UZ4RbgHfov250f/eVzCSX6qzLukP6eG+1uX4xyQ+qYDv8rE8uCB5anPSIycnyLooTKtkl
6MvCaipVBi/j6OBQyKMfBh2pDe0cCvvbFmjGKz+4FsDgHXSuGmb8amonPtTnWDTrRr3YZVUmo2N/
C6rDD/3gpZwWrNl39I3TppyCbmy/VusjK6ra+G1VKXUmGyMGC3lkZOESkbKnq/4rhUyKbwgTR3Kp
5a+qnnR1/9CE6ifoUxhxLqx2n1IWwWhtIfBNTof8BhEDLf/U6WQxmWzKQXIgs0OBUtGrYkNANFF/
r39zrYZO//MYhdibNFgAbmaR7d2kvc5oaRt2AeyvWiw2uuZHFkxNH6MNfkVE4K7tkbC/2zwMDVOv
n+Lza5nmYnxlurOnlwNOHVPRFS5qv3NSwErFHpxXUBU+KvBg0Mx3A4G9Y/y1oHi4mh5EVPquT+Wy
1AN8fZIis4GjazDqYJkx+XqxZIppO6sbpsTdIcuuEHKBEGF+MF0BL6zcPscMXCtQVIQPcjZPPab+
Ys3x/uTRirUD881XUJ329mgP50aGsZJYvSxoSZFiwewX/QVyC22G5zm6J449xph4S3ZAQ0t9eG9Q
iXo3v/X0YQso9CeCiGXEztjjRehka+4ZgMCRlp6dGu5rzaKT0kP9iO88QmhDD7/1ifyyVmqhQo7j
fEipo6AaJfkVnxQ5vR76OdWRRhiMly7vHzRWlcsAor32jNCNKc4KVKShZR+Ybt3DHpeyjmA4KXZL
Xv2KHD712ccPAFNQHkHcjZEhCxFYqP1hAGlKIl5NXXK1OsTYNiw8zBVoH615RwEEtspZ6uFaDcIC
+0X6AaFWV8bRkjFkb57ZNS8dHGy+7ldcOaMx6RPmt5Fz3++RqH/V3+LbxjS6Z7dFdGsCvrcWjb7L
pEH2QawLk8O2LkcEWG1T/Jt0nAdjI1mMnyZQAFxDoVO+id5e3epne6jUyDzHZzOfb5meo5PvEH+a
d6YuN13vfKDQsFwNiKxauxT7YGz8nP4i9bh+ZS+SGqbA8wzvSC4UtP+wDPzYaQiY0BluFr5GMaqS
+H8IlQIoArxFNl6+EEfb2E+Z13EOpnrMSM4YD164oaifoAiRbBNjX0WeXmIft4On6Kj1KNOtEbsr
AX9SPJRFR4MAzIFptIZ8hQ0mlgsxvjELvXGgIV7zZdklxyv1zkls2D/ZScpX66lVh9uPeYRZ8j3D
OnPLHmgkauav7feBNyL8hCzJg6ByYBTd/7dywLDdFgLpKzRHuqwu18YQQWNMGoQeD3zPjtRP0BzF
Tt12X/xW+Z3Z5wLRdqRCDZQC8aMTFSV1GYz7R4p5AAnxg4Xd0YaIiNyfNXFPq60pdFqOOOph6OBf
zZiG6nmNKkSFMW64tBD9QbIZbYHWTZtLDJKhBlVqDNiOjakK69MXGsC93febKjds4dkl3vQE4orj
MgThqtdwpzyGv6urZc71QG94dKUULBWdDDbHSR+IVi1WDiuBBFwoLifeU7JpNBChDy/kWu/V1vZN
xL3m1altoxIfUqpe6+Ify5+judqBCnCp3pG7EhlHsh4kRmGrOjqiD8np8LdvoOUlpITIzh1AfHrY
I/OTZRkcHKkitZaQigDRYXUw9T4OzZw/ovlDJM+y5BubHXehDJ8gyi8qEKJZ82Ulzd6pMiZOFiUk
zuVnhXUvGzyIJaAq+DEVsrkpU6JASDM0fj640jXn59JLELV83cJspMpyMrykmaqovfEoERNt80op
EVhnxTs+uGe9ptOgBSALVrQR5UTjTd6kZTDCvqGUxRfPyRHXHB6BtRIIoDNjIc2TfsSTYIIdoOAR
qGQ3sW1LrCGyd1nItlIaMJRn75M8S/KucUFgvaYx7GUhT4Q4HBe03YXzGkB8VAF4FeWktMXc7Lcu
dY2MVLf/J4FX9H/mLkCJtL0qR5doUsVT+x3iDRfjU4RqxaS94uVzeeq+6VWJ3y9DRM7wmQEcHkCa
MCGEpSkWbLcsJ64JlWKYgHDNBVmufQ0xQZ/Qz93C1+90SgMcSc2p+QqSvSdJdLSCxiLUqjv/nQSz
8k/o4Nt2ffxfaWMaZLz9MRsK3MsyBzz98uaOgg+G2LJf6uvulLTaL2VsDVhUykFe3RxptrWL6kOu
r6uECP6vuRWnFv/76gRMIJIa8B3ZwpgU7p+6J0uSKgE13E1VBhExAEOx29jHBjUjHeNSI9Hiy9WD
OadTj9TS8nt09u91/YpWGQtozHnaZC787dleTe5fjDs61LJsA2Qoo4/C9p/pno3yoRaIkojHGk5r
NoVUuwXuaU+f9otX6x2P3QCpaXbxybfS+QUGf4esr+mODMFf1j4UnsRj+d04a9g2IIz6fRmbkzjO
MT6jhLeDLNYZZ95QDJX7zGgeISvrgBFadOnKonKR1QuP8ketI0z8UVCLuKwn9CpPmzZw9qFQlOSt
bgzkyyPoagBPOxOE0CnHUQvzRTgeChaAs227aQNm27LiwPq6qiAuYyFsBMF8iph5Tc6m1JEoCplg
/mGj4uHldGSsPUbhMTtoeus0gqGTow2s5TdPRXgwXZwOdxBcLSpE41idctTgpMyY9FvB7AAJm0Fa
1LMkidpZPM0Cs37qa6JXKgjk/nWLLGCji5Q52kOtQBOj1oaTpUQUunOob1d0IjNNuyNR6xpjimdd
fWjQ50HLru0eFhlB5k4U0pCN3j35bW0KFPOTrX/ie3SXMEFhKV6xg7cPxcLzhZC1SeS/DxtUFldL
fnT9gZSsDyVkNbuOKklAj2fGna/FNeB1oS8mVmAL8BPAXYfPzNpXqn8QIOd2N2CZ46o2VFxeOwno
Ip9SEl9nLzyCa+01gcDAc1kxOCH/vF+3k37sEJuVhGzvPGYtijEryjg4pBDEY4Zhemg6SbIYKV1I
G0T9hKF0EQWiOqSRGdws24HPl5LVuSr9QTxCCc4xuJbmf4lfdwSH47TrrZSMd/+UR+aHe8woinng
LTBP62zOT2au5FiLiok6iIu3YLNopsxznxuC89vQ8uVF8G+rB4GgGHyNsc+q9NJP7EbMfRysO8nX
A3qM5j5Z2sP0emuyLepVVKaoIf5J4QbKDfjv86HS8Jc5zeHIZbXMoyJJAjIFcpVrr+FZuPRGAgVv
A90oxDFcDK/4yImQSmb/nQTn/2eUz8mDCDzOLx+TKednb6UsY/qokH3cHn92Bfc7aGg3eRqrKamj
gra6IhHGYIN75BHY9id+v5qOPW3iYWcuDdX7LsNtKuQzW3veQdayiB4dhJ9l6f4XK91FClmZ/BZ6
A8OLyAdUdcaIZXKTjUYG6sI6h16G1OdyxxdRFMVjPnNvPNi+AmFNkftmmdHx5S1zfxBY9T1H/SBY
R8mbSzAeefd9eRZZomK5AFLj+UYQP39hvNpi6IE7SrRlRowcMwBJape1ORN7sy3Ugo789UmUKdws
tz3RfH5tz7YDhNto1SJaCdvE4IduDv93uHzNiS1a64zWfJS/4bQVcE63n4FuupP0ZvP4IVPzGVcH
IEIYlDgws/x3xDYM2btroIIS5fNTqks7lKxsOAqmVw7nd0mbUpFZUL2EhvXDBRjrPyK8/6TwziFI
f3jLcrnjVKDD2C6Q5mzoYEffcunnPGlksdzJat9C8r6HmEivprGUimDt5gwn3HESCwhlvdnhjeA+
tr1tcRkULH1sj4sSDjQa5ANTbFWi8L6miM6SyDTzBTNl4n134+iD6M5IO91o1BkSrjA5hNLN2PTq
5kaRfP5zBtmJQO9pOxwrHtx7a789E80YrXRCWYHvGrfuoFEvzL9fD+kOs2VnmZ9FdDMfiTCTLUZE
0CVrXR9mYTPR0kAYogS8H5K7WOnrStPx1neEwqd5OMeeazsrhjPY0HbQa11Ivdzx7aH7vH3WiGwN
pzmPW2EkM+AmchwyOHIoXo51SjvyXeyBZbtkbtTc/S8bqFUDgKuJU0g309SrblcNEjrxeYqtvPN7
ZsPWIFovcDKmA1eHQBrr/fOO3PX6FzE1c8RMEhzdmPMgi8Dq8Hwci7hny2dnFCz6suEnQFC52ITv
VYRfJns1Xz2mUHeGzcAPKINWYnd2zqqpT5JJDJ1V8afYKz0wrIdF2j8WG9puIJw2ijlgZwfQnH8A
IfDQemb56IkWCNsw9uU1zZCxt8SV/tongAv4fbGzFYRpHpQFvU0oRmLDjpMJ9W0lqRwjmoob7oDi
u0dOB96u1w7hG7QajSqCjIgvTGYCXpEGR+1SL6+T8yn/iWt/E7kBaep6KTwtrp+zpnEjNM44NS1l
UZzA0YGNNtSviXqjr8iCnpry6OUhW3bpwqpUct4SO+rYFN1GmaxAQJLa/aMVRcaHUn+IdTx8rq2H
DXpnq8lqEYt3AbgS8lwyIDIhJm86zYNQOvc8EK4Ldj4EuxsoPyJkrGTB+EQwlLMIj83tOZP4kKnt
9ci3+c/V/wUD0a4HaRXYY+WE4h0jm3/khPQPSDehvHIEqPkJEFZS7zzPup3yugsGr7k8yLvpRAlL
5/Y1W4Q9yeNBUdzB4oxaMmayEUUcEY0RwmoVGKM6JOV7wft7YS6+MskFjcf5QiORltXBSZLQmfzP
j7599prS+UQ/FQO80fFrvmEqPkyOcAf4N9c9gSphd4CrL2wTTpyLU2uCceScc4dpv3pbn/9IRCTz
H+KKf0yLXO71IkJJilMl+Kk0rKdTBmeKhbKDZ2HKohoesI0/rOR1KTZmg0z/C6y+QhHQ8jej15w6
fyUKKQsO4iV4/SquumJrT4Mc5x13FCwMnxphxqjI5ahlcWsK4K/+Hf7cJjplDSVXiWZRoJeCW+Kf
r8jFmHpLu2JHa5cx2truYMS9MZ5UbHavDsAe7kFvOiSk0HiAMu8iAPHCFpSaX24MbB8bNufHeaEI
xQ0VANaIUmmUJNMX/Y0DfMx7NRe9vmSj3VPTIj9qfcApNq4IIbkCcEvw6BqVhkw1KNljamOYKyAF
O7RE38wFuKD7xDRQ74MzQiOPYCGm18eZhA+G+wPnVwXfdeH2kIbXXwK2e0XuccdP16Rns79l5oLo
DBk5WyD1TMXx+JaAGMDaC3blkjd8ZKYdceX9D4xMRqIgANyT6K1WEdp0JINZfnjr2zbUJ2a13mBY
DWkE28cYRiqAx3Ow6K9Jq8SGjCsoLiHZyqUm4bH1MWZD+twav48g/vEDJnMbRzlDoX6xkHkr2ABd
4d/xODaxWVrt4NgbexW/zJmbhsq9JfdcDJEHfegJeTGwkg0REFDQHu+wyiL/Y6gN5Aeh0RyAy+lG
yr0XBAPIUpgE8ZgQx3PPeGhjXp4JajKa2ohw7opU6ZVftiyNKHvFV1+qu5gE24Z6XX5CVmUQ9I2h
0zkoh/MBjIf9zIT6BUpXDd6etc8AbN3d8coM/OUchDCrTUppSUzABY9R0bXS+V3T0s3jF4VWF1Om
bRdFRBbSlQeX7pyZWcw5FgH2vvGr/ih16zjv8naMazmjeMhLUUuzbbJDsWkbeHl+giGqqsuLMU2P
wmGhfva9jHjLnCHjHqOrla9fFG8MK2u/D9QlFiZxXj0drjh0u/KZg7A2l5gU7WvOb/57geBWrEOI
XUW+quZRiFsO+qJxN2EUZMohNVBpyIw0H7n65ZN/De+VOTlrfqNYefvl2sPfliOr2p8Zu8ArS7/F
6NB7TX4wgohVrFRlnCwHf64iANlfbEPzF4nS2OgI4kGK8pULF1lIYFB6E1tdyWxW5AWKis1InPre
ZPF7IHBZwI0pxiHRMNmIdpOQ5fbLAOyN4f6HWSL4sxt4WFWo6Wb7Ya68fQuGeMvH0blce0sLEc9A
v1wimH+iZOf7RVHb6wgY1rkCeblR0nzmpkj+Uo8+fxPYqZ/MxcOotybn6bYKe+DyZ9VnLSWzLQih
mlNDdx/62agYFuYqmTHODLknh9gA1tWQVF3zg1iPC6IJaOjJDKySkNV83/Rx7ow6B+2H6HExYHv1
79CXcVXfL76TE+r6UmRLQcq6pZTr8rVuo1oxYGA5JqtWEfBvAeNg1U0qqtisGh4VVzfmkQSz/ktz
syLxZ6Za/cEW+ntVRvl2LQQGA14wKzBN7NHBm7gCQMhRQgOqnt3XXbpY197Bsz522qQ9d43Sz6YW
nvXZ3jgyECds2ORJW0sv/pp778RcnstNb/cdtxCR6IfARfl4a+iJA1IxmPJhnifhVA/9jenweh4i
fvDPhebcf4tqCmlHjnNQAm50tWkk1c4FwASk/6g3BCSjQzl83OmgXmChX824XzdSok0EFufIkgr2
oUJs1EkOFgASch4xGF0iuDD5HoYOFcN9x9dI6FKusFub6DIGkyKumQw/S+8Eep5sEIbuD3Oq7RsG
AYkf0MASlSKuIox5//nP1EVUcpDtSCHyi756/QHLGtLXTWA6LA1CJRGq75WwR/RcjdkdbBYVBDe5
OOvCHN3fU5zpQ0FMtMhzNzHQMa1RWqelHvF1skwQTlGD5hd0xK3Vqegk5/+id0ZCNQtMX3e26Ct0
lXeULHJM8Si6GUf/RcaMf3XwBSjGI9WZsXsuh9hyt5pGo/rMm8l3efvR+r30ILaUjls0FUq2wboS
7mUzw4R5dMLIDQF3S6OIOcivEvEFLINIbMgWr4s+0WNY9IrUbJp8SAJlOb1T18T37dIr9ZIqzBzs
C24YT/fuO2dtWXNMQBfUQ4enZPcR23GR9VUlqgVBWMnCBMGhwUcUKdfdCG5NqxQtKFRgrZ0qo18c
a2Dw9OZ160WbZWc6dOOb7C6kHs0pNPXJc7sbpCiO6v8AJaW+exJ2OyB37l0NCOAvvJm4nJ998sNn
CagOraVV0LkFz3B2Wk4VC1kcgAaTGAuSIrzbC+wSkj2yJvidOKT3midevFrFlVaiz4ejB47BlEig
tojPyuD06wFur23M763v8+xi9k0RZrnXYhmrfoY9kGQ0eUgsI9RkOb8V0j0fKbaUsEe3dI2BNglr
vHC9gUwRMgHeTiKNcyDa2aYFuOnCC+kaYMGbgn8+nonABCHU+Saq0z/83bwmq71IRJcHqo8iErfk
IF5gd/453ritEnLrNEBlyMY0mP8JmjOfMqcml8zwBJXNHXKZCN/AkH+Di3VBOSUxsyliDCCx50cQ
UvMUHnLMlPYtZU5xM7ugBO8Ba8exdGBaH06P5G/By5vcoTcW8nOPFTZdVRMddwRnKKGJ3QYBksRL
43w31xQkxERlkvt3lD1ClL3sxOC3Puiq7mGxInqoKL/1ITtujq4VygJ8c8Az5ix2FY/hhwGQQgwz
y/i585KwGJcekJBmT0+qbOuYslzo7IhxlKg8N6tCzwfbFmOZyxyQKRc3I492XrS9OL8ZpRJS+6em
yi9J6v9JWpszaj1M8s9LuY5TFbvDiVSmR5pA2CTK41AXTpiMOuzWDKrspY+ZNXW0PAK+h+BJZqD/
owGylLvE/yMEs/tqXBRz+PuH1oXDbkWbYQsH9sgsvPFqZwGa/N7tPKs/RDZm/JDB7xJinLg0uYmm
3inV6v1RTdu9jYOvcA4HGFyWTa3rdnR+DCSzeInqRPzjEc4rh9S443Jouim1KweNLUDqEmtcI5Ov
QXwJmclFf5L8bNCIzjljcaeJ/rt8jJHfnyRpMKZLslQ6GvNhOa/YbI6VDaCnvmQnQy7GcaJT8uzd
989MUMCny1IKCV6bkVFbMvR29gFoKWil3sLir+sDh0AfZ+HaWoAoh9TD+xDNtnTP6U8vlBJnddZt
+9F2wiLMgJRlFvhw42CKbp3kABGh9l03BQeUeye8OSIAh3RzD12BETdyCQZxiTMOwbNoaa3xXfq1
T+gBZya4DWCuaeVaTAyq3MSDK/b/HR1fPCbpmou+jVqGPENmHZxOAeiPkJ3WAPahBiYmwlms6TyY
kf7BMG/n305vblX3qiUE26EEZCqoL9Q6sF0Db7xdlaGNXbCV56vqEPhPO5CdVbnHuh11ft1cXhSD
dANfwNd56tPhrywleUzxFzgNH1JA9TBniiOTgXXYsAIxFxcfa1xTiDmxescnrF3fxw4yzc05MJzN
CriWzUadgH5c5Od0FDI/nPQ6DF6SnyNmO+2VAsDe0hxpt/rLN/eqM0o1lFkWV3Vv/Eg+txYEzFI0
I2/rbn4m/1hHRofpLzbmyd+r+eSAlo5rwdrP+WfpR3ceXOkm8awtlUafpMXLwNUbr/PeDABgXcSC
5dwMsBqqjMdebi3qp2mkYCLq2Aav71YLH8FsCZH+Cvzt8lv1RAa2nosX674enUUF4kMMwsWag3vB
mk3s61rDThcFWMjqkINXaNSyg0RJtsLSMWoRmBHFiexd5UCPB3/6v5RQvCY96IqgkjY4bht4LiTH
CVjd6xr23ZiVo4rJdnpouow0sOf3B493jOBVR0yPOVNbJfPgz5DVEqx+jZCLc4DP88yHwlRP/9td
ms+QPBwe/XZO8B2feBG13ahKEx+FR0lqS51gPbJsudI5JJp796Z4oFnAYzpvZ6qoLZMUZn9ZenPv
T0In0c/fDJooxshRSUVPSWFet5W4j12QaSppEFsifpr30WOEsddFwab2Eg72AI3MZv0v7vnNkEuw
pf+dsL2tITuPmp/VDYxhwnx53u5ymIcDOKgYKTmoG/J8BwfYW790VzzCybRd90XveRGndoijXRwd
jMi/g1vXI/7Mh+H6WLnHfFP8SWCn2wsUrmzV3wsnlVLEqkJ7wtrOb2wicZ7SJKxpizaxtuQ0y+Gs
ru0R6ARWXasIB3hWM+dYwG1X29cP+Jc50xDOehVWv6e7K9iWvQka57rwoL4DJttV0GAAUFbL+zb9
1kj94hejPsoj1afawgIgBkSkz4chMsafMhWK3vAymJ8gIUUg4mK+NBU1OvkdRjB7byc3W48Y7Jyf
vIsEUukwMiButgoV4OI+3fD4GRGYfB8oTb0jXfggQ/eaMCZUCVF7pUAfGPPcCWzLLDDjTkEI1fhn
E+WrN6mSllzQhmtFi9N5fNKov+Tp6cTkqOKpTHfaRZPQyCs8v1Wpu02nQt2Ebdww5BjoLZNn2xn3
TxGSyGQdb7A8fW+suQnt5tEkUFOIxs3sb87+mDAYs/gVB08tlXzfmdrs++gZGo10Hs9MdFL1Jccj
UuuE4F0/adHlbcF/GxkL1IU2x4wHpy+M7wJoefxn6IdgogdbcEvKfw2mCWB0+xjoZ39x7LnaX9wi
tqDPvfV0zKmtqLQDqY+R0SadNI0YbQ6t57IMrSbFU/js9nIqw+uZNHi6Kjwxvm7GPfIBLfbAxrAG
NzpItA1GktmxlBjbQe+mfco3o7o/Anz07mUl+fcuwQSLltb+mH5Vfwh6YUGa5OrW3s066aN9t/Hn
SNNUD9Q+bYDm189Fp3AvuvN50iHeWjRsWh72rbaG/jnzC4g6xZLyunySDcq64irCaESjRuIE4rG4
TqU3U5uBbXgLM28faRo394oReh9F4lKo6fe9fiiRa3u0r+kWp7Mt7xr8wkyztcYYm0WmzrA3iwnW
xjRhFZ8eqIjs4D6nRUsnOj6z83ACn9cD4AoZiZBX+dQ2UnXygYJhzfM1HNqU2gyrA1owihbP//+P
EFHTtyYbEPEK+6wzGYWfa9lgGXqausN0FY9TVOlOGYNW9ogHfb6Hj7FMviqlcglaSHZRGgAkK8XD
6t0MKrSzV0UzyySRYQY3ttyOLrxXdsOqfGNzpspHrSAiiZtBbOwN7v4hTs6rE3GMgI7Tdriitq4H
21vvRUZaPsPN6qB8BhWJcrbAv2ro2LjEsTne46060ED0iwPVTn7Y/BikFg2KLL2hN1sCZywL4tQT
YVNAn7ANj7WM9sdlAvTrX/qM3G7lhtSLBk8LZi0m1r4ZIsdiYkr6vaLKgumRYpofhtGuw1qFwpwI
0jIAbOOV7gbvCxMINM8vf4fumtCLboon8nqs2zrbvcuTfDJMYJXDFcjkv6wf8Qz036rbXOpIOYY9
KAFYBcqd46rOVtsvsSwb/zTVrmciN1lbhBh4le2LtjvWftzxhLotqEEGMR2+f5OxOcaDE+5Jiahx
BYzCRSAcsLFlndoNXUquMFSnglufstmfbfkSFbbczLueEWjZhmsQaadL6MRuSIHGqm6WMzV7DApn
/4mVAmvhJvncrHRrz45fY73d2swe4pCuHqkXeRZuCxJ3Wfgjyi7hZUF4oinY9rSAsYSFM8Zan+To
6SlPq1XQGhzhHDLC6jzhIxxyG7Uvx/KQYyeiBv/HH20muqZZewqGuOOgqOLnazEKdJjniJt+/WTT
z1J8SSrB8PVdTABJzM5+0KYaYWm0Rm74/6lBwQIlomxLUsh8VHYubd+qsH/4h+s9+9r+FBaL3jT4
7F8rBshrn4wllPE7e48izBjcTSmqwu8LDS9MXDBkVoIKvtRV0j6VakNzSK1AF/i+CimKGb6uMzAY
fEyZgE3gIFbqIsmFgxICOKcElgk0jrq469AydaVB2q5R6d71lSfFd1tbhvlkvz6qW7JJkQ0U2Njf
krRe4C97axUkjvpCpCnN2pJyGoiyXTQga0lYvjF2AD0aCEy9SGAia/O0ytJbz3SxpQbrjuD/sLkM
4WELi+fJcwE/fN09ofQ7Wgwp+Y0V+Bhx8GR99PWdvPqTolUVe0t3/s5P2ni+ECAXs/4gZF6Fvk31
kZ2RTnE/k8rYwFB4PEvVAU8NWixXLxD4fxuSkvM15JfReQrpQLBngwr3VmvpsRmIMcnUREiSsHbC
x/PLr45F/xz4NsehEcpyR3RNf5/ANf00geOUre4CUASWwX5Zpxeg4Suf0lAGOb5m7wCgXM1fuKub
BbAuGLGr5qQOktREUfuRjwx4sNBxbvwiEXUValvL1LyouvEzyK9DmOaIStYdlwNhwgv6ritLLyqv
31BfhbkAmPFJy/PZnnM5FgOzuxWOUPPTZQA78G7e7ReiQhEFemYXp/61IhEjf0MbqAQjdRj8qIWy
NwYd6oLhMlWo/T9u0mpDLHQh1kN4FqKXvpe+eI+6nqilMcgZ67LZfOrMi3Fg4JuzE3KDBt6kC+iv
s7McfoboHowPV9alJmxVJ0BZwGdaNc9eJG0/9sjNifBlKe8yaKiil2Je1NXDVTUswcL18ifGbO2I
TtzyVBq+WOxCe2asY4LuDiQkGr01Of1Iv+noz7jLuEojevank20QxSFa+qNsDhP2CdmuUH+6mJN4
L8RWNaWQKDWhnGhD8bAcXH4ooImuK17DzigPj2FVBLXKgGIMNdg2j0S3gf01o9BqaxFBqjh9dX4u
a6SVxYKbB7XllJPncHAzPNt8r6yf+5clQL0c/yyV/wIU8tWnosuvs7ilmBNqlLcvTOkv2VvBCimg
DTh2ncyGWIwxGXKtWfO4hyqeGtsPYTGZQgFoX2MEpAI8FpNUzcHubTu+9ctfwHxEc97SC1wjh8zT
ISskQgC+SsHM2aWD/rUX5CutHNzPOLNaLyIp3B9ANbypLNZCwAg487rgZ+dkulCamJJHdlTehuMU
LTrGdVkMETSWwdeqdDM94McpNgvqZruqXStv9slA6P6AepnjTZwbPCsQMXDVVKZXgUsJz0IVZtJZ
LAIPQicQsDTj/QQ2eKE4+kdyfxJ73P4pBs94XmngiCp7TJ1YDpYnRi2nzMPw4QpfO1thtW1vrFcU
J0rbn4ElOmEyKVPbhZ1sE5ipWgnG1YEwr4Fu5pRK3PWQhUljKW9VVnRVwtmja2gROxR2XfBJDz9C
gz/CBB4BGxrPQIM1rz8kIofnc0djer6tRsFafd7HJIeKWMF5JpT9Yh07GHds6Ata6cvjchi5ON9x
dv0Go2BZG8Qjsl4Ih442GKQYwXEHqiWmm5ULda7g1HvSID5QNtnqc6eFMMVqCLDVeFt5z7GrmCqI
FO83Loga71j+72TRZIr3j04YhMmIpRxmF2v/tfOjQRv71yCZv1Xb/pPejldjnJtyv7do4WKFQ9sO
ayTLBCL6dh40wU8eJF1hcSOltFv5eIWBhgBPwQNTBiEn6dTeFTXsjqcicuzt720WimCTuviJvoiT
zzPitE2m/UNxiwaogu3lsoKd6jfH6FJqFzmhW8BcEmH/bqKAWnK/U4pGq6iyjD8aLIm/2Qvrr7rZ
CwwnO64KlOmbTkC2oO7mY8xJneeFFY7GsUEH4hDI2SS4xMNSj4ODNCP1bZhbjhVUeMysvH8e44Rp
WvTTkUrEpC9UAt2mS912t8k2OTw1APqbIdf9gCNa2VYSsxWUTOkkbggd+g74adZiEKHZKcXAwErL
I4lVnscQuzdEZa+9VBkKvqBRHTxu4nCEbIVyZZInNBs/xl8G7fg2LPp0E3j/SlxBH8XVPO4BmszF
Tw6FwS4daSnUeFgmZtwVaYfvvo9lAWV2z1TPMkoZ0qkobNaKp0l+RoVZlUodLgDn3qs2/y8Ns0aC
6TmmqKSRpZZGVOf8aK8pAkl7WrhVKD+dJZ8UZIS2blp82pYxQvxZW7OR+nPfKfi02yY9Cx3dtP6n
QvATtvIu19ILZPuoVphAwTlPI1FaTcX1fVS8OAlWmBoTDDC69bfCJ08tB1BGlNdKpPcOsDZ8+Buk
DETbiw1A9/dR30bByYcfasYM7FO4ixkKr8PPic/CT4arCeQlcQTde9Pw9LT1/ZGADjxYu6L/XWaB
Aw5gS5pXzmgaBSEf/uNC3ajQHkmuJKJysrqAEH14KB7zQcn4h8jwR2EG5snzxQbsKmBtcKYvNGHO
G9CyZ0jBN5G2z3mm5+nTkwQZy7YMdMiXNLJo6Sfc8lx0ZZ/NS4P6bjK/C1oMLIc68Mnp1kUthXTx
P+h6FxJcrdSh45LUaRJIIXrrULGOrZUnoYV/Chq9FIlL62yGbPX8m/HTrhq8eVLV8XCzYIOyvOyM
dsA1yM9wKn41vhc+S0d5RB7oDcYoOxhzz/Xl3duRjxLOaxvTpuFtO15e9IkbV3dHLUdPfi0UBorL
I3mBlk1979827zpig7JqGu6Ai11yPkJYQQ5jOU1AOnhjihK81imMc45hrbuG9AStTOgA735K90e2
QI9wjvt0rqRquSJSEZt4fDV4NRrPOPki+XLWk3GSB0WmhXpp50tUz6jCVGZPJqMshaPHcS0ztZF3
D4nUR3/SE3RXksv9zahQBuvFpjU64g/BGXien7yNtVXxaeQ4VvLRFqY0BoKO5+rPTY69X3TIn8s2
w7m4iJU66qiDGwVI2roQsnTzZs8j6PsLYLFAEEJc6KN+gkBQk+vdlE1grtFRMtE35GOfTop9uon1
69u6qGMQuupySjPlbeGw7FDm2RiuH+qYS0R3ugah2miEPnCjlcZJqyhMzSCgx8zHs46CPFYfcseP
8GASKGmWZO/UTWhRidHyo9MzSLqDhzCLK68atfXX0jBRq0w1Il4XPkm0PbxysPU1cHj2u/Esb8EZ
HoWDQD2IIYyqG1qVjLW+v6nid7R0DzgXRSVBaQWxlKxfRJH1jODHPEJ2WTPasRie3kdL8jKt9ij0
/DzdkzxX+fKcDVZjIqcUUzm+6USbKX/CJwTs/av5V7DrCZSRxW1oqHId/22Vy23tj4lhapZyWlcH
aJFW2Cv2q4DZWydYtDi68n4bwVpgB7Y6zrcQj6qXwXPOfiNbUa68sB6XkMp/XCqPfoqK0mur3fAi
/OefFVTTyRSghMTHH/2Wztz2gBkj+HrOMAD28dZxApVpJpYWNyU8MPUNtmjhCJJGBvv/CHUYZts/
5df+FaV79W9bPOzYnChIGIAOjBbovGG210ss6Tcylf4xoqGt8zOfY5NPQk3U9//8dkrNd55AE1+J
+5e2WaSiar2Z5pTg05Yl4E/bW1Yw81g/bFhyPkb20/b2ys6DbXyzXiRZPyrQY+EIBW25H49uuxCW
i5trADgAz40wAYD9wLTxvvjKkF3nKESnJBFCsU8SmEn84JjtVPBgE4ex0k2OGANVbYe3HByhzfDu
++DXB6Ac6+yQRGT4eGyJmrr5bS9rTr0w774VGhaMHm0nyIi7aklpw4DZMGjiI1s/EhHB+2tW6fkt
GGiKQ+lgMlmGg6bYnwsxeXmuGS8kOZtVpPmYwyywqW3G7cWOrJp4s3o4Rnc+KsXhRBC269sNyP/b
rsCuiiPyVGZpUYRvW4fVI/ZSBrZ+g7rscADpSQUOYUPVQd4gbaruTghoODXGdoLyjRAWWpguzRwy
dz2P3/XDcyC8itw7h7S7cUkWDXNvJmwQCri3iXjZ0hUBDnUj12KDdqsdOnErM8aufbvMb4uEXati
bH7SL26VvxY8ztjarjCwjfyDl15xeyUybw9EeF669z2iflrpk8qkUxDhFi8NNVbvFhDx3Fdnd9/P
gy78ekdIFaDGHnzm6UWks/w68pxrI3YuyAp4oo0yAvMldkcKS4EBoxlyLgsPjNm8plMZloNO+Rja
1R1JzUwGCbOJ/WpKSMp0iWR67hkdhbPPIlx5uoZ1aqbbYoGCRkX/9g1L4TReiSwRt4EDVg7CERKi
LuT0QcH9lpPoMu2/U20VGlo84BFND9SL6NproDgPbB4NuUQNH6R8wF4jbv9zUo7XKdCWJ1i4y7fT
xIhD+3k4vyRTd3aYIWRhfv2Pj241vu+ZfVdvtA+1nM7j6RCVZ5VJ3y+ir9+r0P+6uHPM1JY+3UGs
1Qs7xbCfOzieuoSqnPoei0ImcCtxjZpz2uR1rmTiGTC1lwCZs2wvvlbQokVYMJLVLwrOwD+ShTb4
kFrz41SOKZdHozRD2aM7UmDYqjfcWPIJcyzBllg7tEhlR7DLOkUAYlmZgshOg6DoG4hCkglOnNSx
O3xWWCyQbCPqdZYgiTwEQrn6M3l3D7q9kGGtz2lspqLdw1ZJIY3BI2YHmjjq6xB/RlPf1J7mmEyk
ZK1ZqX+2EdjBCVKh5IDJG7Q2lq0TzvkAlzoO2MpEoXlZ3GZpuJeTFYrkCIXPi1iZoibhEd4C3HDm
4KXJyuwx0gNyi9lp+vL0kGyVPGxTSQKMg093CIjhphEJ3/IYpHH7oAsB42twi4qN07VHwEtWCTnW
aEInF2poLubARVg53C0h7VCvwubjSHJc2VER/2N9e1yF2y4v977ILqCw+leGMvLQZ34q0XVJHHJu
ShsbLyUS5jh3tjdMerp0SYYCffyyMehuYlwCJKLQKiedMLnxXwXK9yuqtKJPyXvnErOTjtPNFlBF
BNTGShz35CKtFbzhuafXXTBkiFSaPqviy4aKPAvZ5Jp26MbolemjmnyYuhm78elj2QgzqJ2uZe21
fg9lOL7uMWwFou2J7iNUrdQMBzzU/kSeQS9mdwEWNtYM9uYcr+HFHDs13VovQZ7Hp2S117ksA9+v
F5LmCDfETy6qF/nk4GfGMn3RwKC2h4Nfxp1XJ7pvlpmd7HHEaKppaVh3PdyqNI9jlU5y580DpADK
O/AV5ORSYW4fpzUqdbmSUwKi9ne/avkSnl4o0ajgDxK3+NDIiaIUFikViCHBA9UJUo8oE1si9FZT
ozDdvoQG+yy2AgRkQC90exnf6ZQmp5u5Epfvpsj0m7L8B0m1bPKP1VFD2/ILuCUYezn/ho3A60vx
H9W8jPdiodyWl4mWOfLXgWLVdcGamo3isKLYLEjO5F4IHvEDya+bNeemuouxitV0DadjHLHnoWj6
tZLOzcuoUjA5PMW12NkuX2ExWrAhz3dUDOCj3OdyNahGCQJlx6eD6C/lsIprW4hHFOLcn50tklGR
YRS3YeIvK13Ng/Vwm0KISYdfLSwr4ndU0GB5V8VCpunfH3o4CRcg8hkubUGfY3Sa78E9nUgNyoik
FjIV/R58nzrEa6qbP9/0dfmx2Lmm/vS0KtxjzcrXJmbUvCKSGurt/wWoXHyXYNVVeF7875pzI7fj
bSVv8GuqjylunA3a14hN4qfjgHpTyEifvGxl4jgbhecl07gF/7C4oiHKBEzAj2AOwWKmN/+OLeSr
hNGAl4uso3aFMZhZ0GRTf9fJWRNUvKE0g3j6okeVmhgwTM7/4e+rbkFmA+gyln1e5+4hbP5isd+K
NzV0TV88fXApgTqHIs0zXdm3hRVTs9Vf5kDdbr0FIWsEKaMI93YmrEGxTyvkgIKZacdPHGV37OGv
9tFV7tPplaBTjPdJ6Il42oq0VhvoJhDPiJZXPMPdVw6N5wV257k9Dbd+gaxKftsPgyGnImvZiLNh
W8I+2CJBNdPfNg7x+ec4LGh/N2V8tZ+CKpaDqBqKm2yo4ckVOepDpTouBb5u1v/LHeFuRaKKnU2y
HiUOUYHKYWvNPiM8aMPMSO5rHz/wrL7/IqJmvcAAEdWBWiwkLiCAkb8zFfSYEZYuxOj2pFnENaf7
Yx9KUM9S1bZq5fkzsnBbG+/7NFXfl31JORREoWybu81mec5FJYtZXlHJsHU/elOKCsr3ud/q8idO
3mQT3a0Nakgb6b7ULZNh4DVknmEydxEp8CH0Zl/Vz2xwA7Rmrr7V09kRGa/6yF5oW0A2akLbVUCY
LUDYnCKgvbdrbPceJfaAL2eKjadNURaR96KBrHPxrwzgGHZCewNFXG3NNvIH7m+4A3JmGsrJ/3WO
jiPlol06YoppLHxjbZofmGBEZNhu5JTvL3uzvxo8hVGLKOsfPrHdqySOFKMIKUILVMRCyN1mWGCr
HLj7PyphKHNVTxmY6+l3JZHdWsnEqkSQNivOZzc1iXpHtveTAIJiD+aZOBBZXnxJIFpkpQuB6Rfa
IH8928VJ26PXho5LbF4Z1D8jpRq43tThJ7MYmyF3FHuFxNEfzObTF7dWdlJ9w3wg0X0oAa4UmOy5
MQtVV2yMFf+U+YXEoB8RTxvAsgZndcWwbJaPqAqpN5HYEir/MEnpsL12eK71jA7lz7zhtvFjnfJ1
I92cUIiStVFJSLcCjxjnU+MPa1BbkW9QFkgq4ADyQ6HXmurfp3oxngyhcZV+GKQ2wqLtAR1U8z6b
JYas+AQj5tynJRByJYKT0BBzsoXtfejcoyctAa3j6mSVTK8L1I3nEEJy4p9Ohdgdofrx8kuusa+1
qIhiBhRLnjf+mx08mto+GDOsKfJrYjMY0hTu6rxXwvuCMkAtCn5iJCK/hahSEquo+i6z21sOhfRy
I01aMmH9Dxa5PvVRSU1R7ICmHWHEoQD/TYZ2C7/p7x7gXsV6wHIJi+vFEYASSqRQmZKrSEeAcJzj
16fTPt/elza790oMBAjsiKncfSUZBG3RK1m8ZJmoOy7Ts7K/l8bdQtKgkD5OPp2X74lJOu3Sd/jT
UJKf0sNIYJphHHABTajsc3QghvLkPSR8Pz7rEqMC3kDLnxzn2GvabUQadoDyMJaa4iWbWZCuH0XH
IvMbwMGgGI7c6FKWKQtRhLUgkGCnWut5/CnpMU8fKsuDY1R8rXUS3FoCL+TIE2RlXF+/3pHm8941
2JC4XfQsWbYCHEOcnB0+LPffGVDczVg9O8GALVfuldCCHGljIsrkaxUK6u4uqHIE19tftwIvxTHe
ycSJJ4h234Whh+b+qYztdmGDjuoF0XHBSfU/OIMpgeMmTNzQ9bQVxb9W1QxQls71qApATFIaKzCH
U3yUx7nV8ltej/0PY0iZWnfTKaPu2uMZtYEMYIJRXjyOXFD6wHtCy6bxWNgAoW0LNj7moZlcf8nX
GAczokq+vAzPk9Xy4nUPxfWLIejVbgy+BMBynE1KUS0MlIpmYtO7EWFrtSk0JJnVVlhKpA/FZ0fh
D1zWiw0MYE2GLyqHoXoYTNZtqknPAElqo45wr/3tJiCJsVAR8ZhZac36nDkqHHLZG502JncOwUUn
a7mAyW033NWN5K2XsqH1DzYeSHIJ8Mp5o0n0mRyfX6G5Fab/qNBxwCq6jB6KfQSyftwOYot0uHSP
E/9/jm4aCRtzNRKwJRCl3oyUhUulQXKq4x1Y5bmJ/IXwkOsxWJp0xK6PSTh+gly80FUYtUpVBZcH
22aKAp10x0Yj1NZWBZAD9kD4DeWXM6LAM6E6Px6xqavnlhlooE/7dAY0luUTXUagpYyWphfow6h3
oUKh2A1nX+6dhtwdh6VZxWVvM/Nfdrc9lCsDffjIHekqlywM1endfOrGka4W8EjKw7kq3GIAO/Qx
5VFAHOwwK4BEt+VSY3G3mmPYpM165zpzO3/up+3/tVmB3IChWGELIFacHPNgIP+cE1/xqRD5nsaB
67QlMONESNJACA0Pbk5otvJquoE3j1kdWao1x/k43BUnmwKWoFQNCvuokEX6TZpNgnbUOZZLX8D6
3RZ0uC3jpOvhi16baG2uYHwnjfzMn2zZUlJPxLYmvsk653AJE5w//PpwlYxhNAj2RauiuYtoML2t
WjPPILLRikoDGnsKVthKUPwJUQ8t0x1DZixQ/TUAhjxZaqMLOg09R/oTVODCjHgPJxUVz+llPBFm
oF6F/1qAu/0s5tPKDWQdO7EUc/MlzmVoMvLmh18NiEROXPQk2e6TQf/G/z/VjFMUfG7tDdKRDh8M
PBVwmNggF4SYVC1xC4EOnfj2bxFiZJgf7Fj0WFk0d5xnWWD2HqveCcnVA2b0MgTPbtTT1fnFl4uR
0x96FCBEch/i7IrSAFotnOp3v+o500PFM+7Yot4Z2z5r+79QlEVITA8wOgOFwr2MyIxrBarD+gpM
yFaYmcra685IuLMIktqLd3wY9Uuvqj8KfH0YPR+Zt1KooihxfmFSipD19Uh6ID1tFsrWMPX9q6jI
eTJtMu1Lv4SkW2gKBIWsgl5jABOOiwFbmst3lfZHWhS2qw6lYPkZx7hEXzLY/LoTLQp2xomtY57r
WmWUhCMP0oTOlA2z6pEm68U8HlOOlGUK5rrZ49zi73qy/g3mLrQM9425+Lepxzow00sm8zyURefG
OYrvpa8tZwVWZsispx0cRkNFQXaqxQVG3+5ZHVv8XtMao3DhseRYrpT+yu8M8d934z/mXktlZAV6
FAp+PATzxjVfy5R6KVXTWMEl8jdG3k1WxRbEptH5AkZllW9LD1EG4aQHdV1j//CR67eUb4BLJgiK
k7pUVNA5QQbj8WSaSF4y5lcdQnO2XAQ4UnADRWo7bK7gyV5uEj0st+GL/YgsPJ6DjioY+9ILJlg6
kXqF7NqH7ndpsYLExav/sCJpbUW7zGzijPWgQK0UB35El+icbeCqE2aqNJ7Tt6RMamFnXULKi3kr
EyJ2yOdW8T8Ow32gwhg7JTOeoZPfgj4w9dqdeCskQsBBmfvPIM4x/ezBPN1hev3wsAVUCaYBYIeA
5/yQwNO+4jWR++2mtSu1uuOqITpX13Bv4nEhFJ2XRdDxwnL/gWnuoURWMQ0SqtAXL/mbp+oEJJcv
ie6IYN0Imkt8qYQDZYPV5PrHQymkYlsq/N58SbzmHBY17Xz5ayJPnJ2G5jqVe6FZiZ3EHtS+LPbL
vuqnNEWw7n6jGeRqHRpiEoDwZNpbw2MR36+bhXUOj2MdB2to5FulKk/e7FVgjyj6rnWZNW9rC8od
T2CzmkOX+4YjPoH2bNVASKGPIsTKQJ8n6BgwtJcv7gC/8L84GayNQFoVNlclhpnlECDYz+bUdVT3
1h2UwZnAACeX7LOu27drAf4lIJGdbxhj8omrjDVBiXfVnP50+uqC64pQTfzkH9SE1aycxKl+1IHI
bpICMZGal0tleMXfGA+wN8Rbe2vQlY1/VEn817r7z8XyPrvToEbt1K2iHiMgBxxptCRvtfXp9Ykr
7mPAYk15AY4MhGWNXWWehnPKTka3sGhHCm5VBwCa5EV5Gg+qhmg1ozd4YBMyO76dbRhmJmNjjnAP
fIWd/6nIBmmrU3rRPTnrBAKbp0VWhCzQH+Yb9YImX03HOX3YIrn2oiOf47S65l11tV+IWG250nBV
RdUyL/7r8G3psqM0BVwHBpQOsuOTvRqCqdd4e+FQ9ExbCRwOw2sXsw0CoLKP3O0wFhLzMcz5txgx
Deds9zJdCrL2k3iYOLmFmJ3SdkCC66ja01wpjFGuw7R18kvFCLxk6FuqtRa5Aldws8PETR3LWiKn
4L/c2A1zTX7znO5UIJUMkgE5DiJPMqeUc3mu9xy4ZZI1gLpoAqvJiOLb2w6oCOU+q+Yz2rOVotej
xfWiy+zpnvCl5Mqy32msWNfcxvyNCJnvcUwfITHBoZZkcmbtBG7vvMC1jAuh9IvAp3wNvoJ17kmw
KoxH/8uFYVcP/TEVHo2E3J954Tu006NI8ZgJ/TlaCYwx/GpEBqoS9u9nIASDkdc2z8jcq47mqFVi
W0Ok1PZtERipD/qHzYpFCFuePQOqlRIVYOUeXdJcir7r741U9DjCUrVPyF5vkvgv5ux41gIkH1E4
pZ4/gikMWVnLFmzgTEpYBwStl10iImiqk2rZN3sfnKbZFvvCyHbPJJ0kAyjRh0OdbzDh/14GuotB
Az9XcMq2prsLdTxyjlqREnd+IF9xjywCfyvlbqP7OIeC0BATJZNHWzjwz8cNekgndGzSOaw2GppB
5sPWfU3ZdzulTDK9gzcT3ZL0Nxmagkmk8jjd8Z3qkIrpLRslYyRuP7+fe7WvWNRzKUSl+eiPdJ0W
PiWu0aHIddBInLY6SXHi9RHE+1KWoXTdWsiO2NhSUMO0mE6vHrUpNCzPTKbogv4dNJEbcDJMTbY7
Ot9oAJkWbxLCIifEMMbmjjtyDIQ/FbWinVdNSjXHZ7B+Zm4/BK2Uje/jePpDQ6mBb3bMC2Q+DgZ1
YJTFwCaBskrewQ1A59hMWoab3xAymMtaRazawd894OuoZeV9oqQi+hRFuOBRTq0Hvj/6svkX+RcS
ovLanOAtm6MAOW8nXXa78s8ZRSoUSV+5hklQWsEx7BzFTVG1chQy0czJI4hoKGuawveQ0FJnVn/J
IsPqD9p2mxq/vhh/0VyOhonG99Eu/0RNmXN3pZp2DYGoRIBo6cwKkRGaeg+U7w60KfvMDhGjJLhR
/Mfhb1+vQo3Dbu7bdaUcJCT9tn8ul6COHYMWnUWWa3tYARwLfhB/ys1LFK3+ivO0coWqFxBQj7/7
7QabrcKzKRFXhNcl7ILt4xh6DG87xRRPYAXnvNCOqeXXf9bPm7smBC+anUrHBvRn1lKRNU0R9GgQ
kfI2wh2huXk3Ga/HTbQm23GZjQ9BtEIxC0J5/RHugkTkDDbeaUBhzv8jGR5lnaLDuijIvowbIUhQ
qIfLHKEvBDaL87X3d5WsDAYU7WAyAncQCDGUpVV2iR2vQ4q7h3k9ro9FyaVatZokZ9E5WKauLt0P
CznihCDroI/DiQDst7r1cid3bb9JblGKVZnF+UgFYRc8w1kF9gCqRyrVbkzlblriRNKbcHj+zxY0
62UxjbalxF9IuZZA71eGB+v6J/u0xoL9dJ6uPpCggxiYRN55wJpao2GCqTtvsT5efJJvD+00bIkq
7DmKN8mn8mrQpP54gqW0gzQtsGBLTtANzKIk00/IWKeMpHxr7PAQ0uDyvJih7G1NitnkTY9JAWIJ
6raIXPuhbylwr678JFYANJI4CK2b+2ucVeMqL12CcuxyvE6fs6x5AQ5wgP67AGT3iBaJVPneSEwl
s/ph/Lup3NVAC1r32Vtlu63xxyvIHXIqC0BO+fih0tjlMJNLhS1TXLUCli7BR8ooTZsvWWpEOzKK
9U+8tWH27zidvjeKKm5BAGTaD0JbKlKhFLOtqPHkoTYhBmt7V8uAJ+BSRP+MKBnAQQCCAhMNupEw
Ad3R8HNBANu41h0tC3dFwdRjW+l154Hfb/W4tXpDrvD7GRncyJxy6IUGkrJQ7deqHtU7IQZL2I4I
EX1f+zvscZ6tEcVKx6QlhjLgSNyDWeB424aR6pj22upATblOMvY7DvUm5O2V1W/EqXu/3PeF2is0
GeocOpJE3E4jtJjaGBqrMwBU3ijmnVXfusqLWdBPDhnlCzHDElpSrRIEPVHSTczYzbZiaACyBegT
jRtbPW7v0QqW0U5OMHCtqQqaMG3mVt7JhaCvrMhdf1bXiC9PjfRMbfY4pR9Hgrzs2c66rkOEioBj
w+IMxTxeLAR/mwsKZ5HHRHx2LeppZau+jaMrq/s1coMfOTBq8FWylFhzTZlPFXTmNgFF1Zv4ydcS
p4uOpoNDkmd9g6AeH7te02m/KAAQGJ4HcBKLqUQs+GexZ1uvKL0wpbUxqbJ+nJg+QxGoiO0I9iVk
qQyGG/fCsvA/7nKKWLi58nWfGgdNt2mxQepJDmjozzNIxHXpBlJGjES23uEZWDwp5J+GTTHGlgma
IqKhSfcP07SgdAW6utXXA9v4PLNH6z8U35MvY6kjaQY/sNBwWP17+ysOkzQX656E9/Bflf4LvyLj
b3BK1ugRrvABpsKD6GGjnmk+ha6jQIJBk+WuaitbJzSc5A/MmvOp/yXY1T5KLIHvCDMYXMyRZW7w
7TftsFEI8DwAs1GEYQSSKonMhYJSN9vl7C+CWgVtZfYyulcpAVB+yeQ/VfdJWG27q7vVAqnpTx67
HydHGGcA3usJC8Qf3efZsRpYa6oUDYFlmLrOp3OPNLSAsG/MLpCRBlGwEYR9ExGULxHlqnSlA9k4
aTtEcbk79RmMfEf1Lb1j/93SMCDURU3LmpZOtpxqDKFgKN4jp4i1HA1xUuc06POQvSwmXvWShmmp
cJJshIiJ0fHDWeRZ6V4hSMkztGDiUv2zpIMscieC2aTZ0l1CHVjOoW1aMQZZch8cgAuzgNwZ6mgD
unmk6vR0UmoGiWWgN0n32reN8Rw5T0mMBzBGWTQdE3IF5hLzU5ZNuHTO2uWWGsbykpVdgAQ67Xf/
rxQeqpY0GGstYrz7iM1kdwn7Bw7xA9rQVHNUysIQFYG92p0T2uVG+l2gayNT2ShLtsGzcCka7/bR
yyIAH/rHbn+I1DMyt2+VtkT9DgQIP48TUVGDJ3bGCjwHz4WgivxfDmNTWqQ+mAHyFt7+8rbOYixW
pdWFUXRISrvchxiqmYOl6bwneGGPwHisPcHtcOUPdC6sZ3MUidaQNWd1V8pdhbRQFR5h5pNxb+pY
7f/iu4q+RYAK0OZofi9+pV6OAzbDFciBFxgVSEtq0PSJvbvvM+SIhXK+bZqh8OMwFiC7aHcmVtRb
9GNFBIvG23JwRFyLZfBatRAq+ze5zLouQhnY0dlyUSaWJuh0PpSo2M/w6ZbL2u3KQqkYUBoOkLUc
2fccy+FFYgOqVv2TpXL7IRYKvDkvTbuI4UBrT4aS/h/+RB/K5gaUU5YgxvY54+HHQtcJ6AYMBdNE
ihxJeRZhD52WVdvNr48iqc7QcNm6OpS8aTkMyqMRwocFKjWVehDX8HXnJlDTQ57z7fxTM4y0ZMXv
/Bel+ToHn9BOE3N/zao+0dAirc3dMUysal7fpz7LXi1sDIixOiFLUw33Yy3tAACqLBh19g/BIpOB
e2mCXvq7YioGKHEMiAWlyyuqVK+dgYcYtDYdhbj40WU+jIMeU/N9lt7rkAhLOvJgXlbEQnngHtUm
3LSt2wTOyJHcm5pj5Z1EpaWza0vABTsgJBuuovn+rTmOn4wXqLxKRSRJiPZAZe95ESdPgKGRvkig
5W8CLMu2LGy4RBo9A74YN2M4jb/LIthethKtuSmHTX69irEkZEcmb6K9Xc/7BRJQrvb2Y3+nzANE
cV0hNcP/Qhu1U1GYK5bn7djHex2A7LLI7xxNov9/JM4gbo5qcGasx9/69uQigwWDSbUYHUmNxdGN
UBq7Wn9qcOkgx3fw8b4T57iBffxm08TyegXWBOxRr3nrJCQ/2f8lOW4bow0nBGyq9t9VodZRIKtH
mU0zZCkF9AkKg6QSAti6/6SXmeXc46SNqPeIVEYIFohSsBae/5PUvZzHu0vUD0evo1/Zn1rEVFsW
JlMPzuWeFZcDStFB3wxnusHxZbPBV3EXBhMRSuhYvBNoMIlIX/oGN/e9963mONKR+crbRMmtBdse
88y2JHAEvCOYZ1fKo6D9uRCl8eFsXYx1mMTefKd5XLtFhSZ7dz4g9+4QzsU31Scd2szk03C9wl3g
sJxr4DxyimLliITrtPfNsNbk5+RgX4Wd3qmJy/Sw7r5Glf+UY1w83TXBfonaiRuUVrZgBOmBpSNZ
OKcoSoBbJ+tqgDg7PFd/K11GSr48QqIutX+c90Xpe7O9xZ8lZ0KeVs+oK4M05+NzmZmgVuAxiwi+
U4mSTBzWvkuB9hMsrV+Oy/kaG2FQyxuW6Z1SDetpMEc+7Q+zJJZULhEN7w/bhd5LdETsk/9EQtzw
XWDnLxW/364OPTFUJwz7iPhC7uxs3C1ouSUQ9PVJxEi1H/4Dm+A6KtHYdKmzkvGC3dB9Ik0uds6+
hlYYAtzz/iCeinJTLnaaD04cqyz5dMt1BX42mxVlptRbIq/Z6+KmwiH6w/Bx5btfJji2rwCXJLow
Y6jVvJTGaovuIV2p7N35tVvEBbZ/ORg+UVaWUqiNUhgXIyEa8X31G3XVY5D53t2RqwrbiNQKpbBx
zQfkA59a5Ck7QLckwoBFDYOT6ARQ20VCCaLnlCRHrbvCM2gYIlITHyH7IHBFPkbe/ZIeJ4YltsYE
xl3YBz23L6p2uQZs8Q0s6sheiFxca9eCH8MiLkhYurBTtNZucd9jSJ9bjwWGLw1pccU+w3cg+wS6
iCbDvCKl1p1mnXJ3c5s0isfgn5IlF0CfbC1t0u0XK+Vquna5rsokztqhbFGkADPHZ4w30NgI84qn
tJDfMrEPK+mb7hSfTEKmxjUqXwHBLev/pLvSfxXzCcH1sxs3j1b+/MxIsmI+PJvWvd36MyxKiltQ
IltoonEPVP95Gn6pWKniDB0pFueJw4DtkuRU16wWxDL/uGqSCxvGTQlJgU/pe0Ty4SlL05ZYya7H
73Y0cGkTY9iZlJh8KhtNOxIbS18iDeVuZa6Mm88H7VY+LJaN7h+WdVDrcVJPhZN814xqJUIOHQpj
bwm3Jcv0vW2z8N3aXLx2hZjUpzqHwQDwpFR5HGDwqhbwFGj1ildP3yinS0KIHGdeqmjvIPG8fhWA
rwfkrfUp619kFuiDJQdBQ6HVTCyRVHSdlql9aRlC3ZkTDiafVVYmqJEXYIg7GTXl1ZAOsbcjmADa
qblRNktAe6+B0zFKfxmdAivfKFcGsyoUh/sKOgI/5z9mGe3th7hSTJXXsHEEES5t2YzZMTlKEGje
n3wCxsCxE4uE+01d5x94hPn2RUiceq3lzwhz+KCpuIeDH3a0FharQJau7rZXPMCVfYTX3ZYwosKm
+uFRwVIzAkrfQTqj0sX5f8w9uinkwpqNOPCHAvrLMJAuGYEM0YSsP8/jHmTPXwHtdZ275P+W57fT
/T4uivhmhdRLxpK4NlyiTUtGDUQmc0blF9hrq195TTv/Jtwfi1wzUL+dxfxICBslCOlMR1bmbhAy
Ga0T5mb5yA2GrpLqWLzKLBWfb7aBa+eKHSt0YoCVRy+whd4dPtcRQ0TwS81IJc9siE6wc5gTgYYT
Qb+xJk6k/yeRB0IsioXOIoIqHtRgINpcCqhn8yC4rihN37ftwE503G48SHUlRT8XLkRH1TvHCNAd
moLTnvLfdUJmiq1ZFFpFlXNmDyNblMToAqvOsKtLCpoP1uLsvVcSnmuZGHF2gWsFdOq4ta4yGyle
gKfcZnOCZF54ttSvawKCoRYuCzCRx/EzAJNSCFPwLddkj10PVPHqW0wYt04VGEFWC0GVFuGFgU5C
GRWyy3pCAoYLpzthCx8ZRnOgZ8a38Gh7VFKk14KYs6bxrx94kdkozlXrYeOPD4SKWYafvKDB+Hf0
XrSf0TqS1sVX1tDkV042YvSKyKcr0yOIpNbMUb2HNuFIsGE8RX0a0i+eXhTfPXXPTDNjafRe4AJA
ZCIE0MWLt0OAv2lMCRv5IydaS02ELptvb17psYlhECDnNi43G+0HTkRShiVHnju7scO4drHSsfCd
5TmDpvFSS19EWCidde/yTsc3sIzy3t/vLLtJM4mRuctjPAePMAI2WL5Qhkk+zH87065iJN0oQD/k
A/BrNIeoBjZlBCi9KmsQZtyDQfjPHieXGcMiiK1VxGm9MB+x606b8Qia9gIBsVZdxwFIU4ytW4HZ
Imr2K7vB1RweXEwaL07b36VtBHP011kX2u0J8Qvw8NtnJT7JNqDgQTO4oDbaUNJdXcvq35Od+D1c
aciDXJSEnsluy/VpFD9cc7R3ucNBLm0jtNPJRaLD3Kip5Rx0DE+T4q9nb4OhNA9NuLnyB4O/XWs6
7h4RqMFL/1UObWvAWDAsmUtHdCIs+q6OlgcRTPAqhRfNQ646BCq8ywBLwhnP4jThx4IOTkFppGzz
Xa7eP7cXJ4S1SI/h7SntBXirKhicjD5CMlU/O74TRS7obWhfzecbWTBOIJwM56ip6XpQ8pBntCc3
VQT3Krt7VoUNZEXiO5SC9Xk/4KZ5uk3oxxzf7O0dWlyBLeSaF2dbzs/XzqaSdUFBcTMpfpzaFAZ3
qDKcX9ID4lM9Oc0rd+DqKwoi4o2PaWSKYc7355H94sPkLbjDAdmSbFGOYb1WQRCxud3lVl/XjDlO
KaY1du27+D4nIcW9bs19oYeKt7j7wwQ05/ea+txOus8PuyCrubqJGYWxDY+rRe3oYpkPeQMewUHu
5ntCDL3UpIIzNFGnvZrDjdwaTxqBLUWqMJKeI/UlmTrLg9bK1O/NBe3k8AoB02IKPAWFhlKe/HlB
D8oc80XffBOcPH8hSDskvthV8mm90R0k8T53AGGwHofqDEGZtjX44FAZBPjLXvPfmbqvWi7LxF4g
dKXXjDESAeSuGCXQZqT4b/J1caEteD88pd3Vtiqd1+1JIEk/aTbrqgwExfGFd8MM2qVWhzwnRXbB
vERG7TKgHRna8xxqbSdgJPB33jfZIxdBWSd8FqSm8nrZs02BEQZRo92MjNFc735g/3akbw8kDMm2
BinrZSySynj2F5G2EeR+bJXg0jH2enjICitysMUs71jtNGbOCGQqnluZVAODrcX3z9I6Q3STI331
dLgBLPbdqdTmLNt4eC+pwoLfSIRB1roxU+Q1os0IFHyAs+KM0NiMDScGhMvd5pxl+vaQp6v/OR2m
y9ZN3GCtRD4XcRU34Tjk/ohzT0GVCm/JT8wknD95gmezmilhVwf/JE8jb4MjCTjguYPSfTCWIfMe
dipydw0SWgE9nbS/545EnDVGvy1eoPtGtoFJcj988QOHHo+s6IvEH0VpqxpoTuREsq4vznZHhMdh
Lcf0YdFDvirvziy0kFIMKpfmGN0aF9O7DMBfL8oXdf7ORWOsdrHRn7LEYPrfbdroICgBm1HpxJYl
nt1CgZIHAE1ArQzcbA65/CiPrs/yKp2GvkKXzjl/VjH6NDIPCQrCDT+pvqXdMpP9fFOLKcmyZ/o0
38ooX8M0v5S0PqmY7FQ6DAoKHgTB9VG2WQVpQikuawjcDorVWT5Bi7I4F7a4hltg/BB6zlonhH15
tNup0ZLiUevqqyAzXMYp4uyMoGHLna30k+ExJofUEDfkoGb3hQ5UVWW+kDHiUGm6o9zwAXKsh9y2
82NN/6+UqNKyJ2jSZvGqVGHA7xEA73ioqJ3rd59PruJ7qHOHip/g4k6Ak2XpZNLQYPYfxAKmsyeL
Zw3CbCaBfAAkL5bM7ewV5CASmAjTnDVSCd4YQr1vR9f1vJvNStMCVwOTh/CffybLgfPBU51BaGE1
bOySxqtAliH8TYaQuQaIPERBTNRrGLyca+XJDxYPpHZSK5GYgG+M0+X0gIajIIwmXMegOc/t/NC4
tUwAOvPVLyztF1YxxVWDK2WZUYtyaUIbs33c/EAAgSlFG7ryf8UciCInO0DCd9Xk696BxEtJKLpi
yzWObQwEOBLbDGDCma9yJvHWB4jtwsI3hAPlkxjedCIKDshnOvCftUYbHhnqYrs59JkRjl+MPKbe
YZ4P8VeX7bu4+ya6XnWmfzY0B2FE65Y2Oj7/7f95Vg26RsPZX4x7kcYGqYFrbGXdJxLkKjefX8C+
ThLy/Bf61UiybtHt/p0xNiqSFZqQt3J11R2VRM72vkgfZPl7gg1SOAb9kgCnmSCxBawkou15nOjY
+xKMrIckMXHSpNzkbe8JFWxbM5DYe1NnntUWwzxfrbVNvYH5NWlctJ6z1EEdsW+xO1WopzQArT2/
xHSh2lX/FFh4IuvvOEctt0WheWoJrIBZWZl9VNnDZIKccgNvOrpLPzIcr8kgbd+ObToz6//z2SPU
qwQXQHYGyXZQmK6WJWtN35fccbe1f54VDhHcVmvIXbZJxYhx4uHQ4Aq+yNmWoTD5qSf2d6VzsWom
ue62Gk5cHCy17GG1C46MZftsAobxxIW7qGZ49OSG6PFds+TJQJ1tMBqT/R6NtKitC7L894Bwnx+C
yFLglV/BtjAedwcFgtANczyjXemTwLFKGjo9aA7FO9fo4ggGUmzdr55qEKZGhC5fvWjWa7uZv/MP
asDxhg353dhQSvgpBXIZGnXMLXcIoVStL7AFsidILn9GuXLJSOotaDwkhg7fM38kdkX+8GHDah9v
1aqM/Z0kwkRlnHwKkVqlw+9Xl09kHTO3hRRPs6ihN1QCLmYS8R363Dj5ow5a78NPkRuNAOF8JP01
dRusFbnut22Xa9KFXdMLtJI/m6AWiqwSFThseff1HVE2w5AlToDWV5/Yrq9DSX2+j+NRqTtdW7ee
dXG0GE/V3WApJnQnOtjfdSlt7hKTkLKdWwk4zM3EyCmrZ2Mt76bqG6AvozmEbW38tPlKl+uZyP4r
9D8EP9/A0y1GRS5qgeUbRNIGK4072MmSwyxeL+Bd7tXIeReoOnna3pp11p0bdbJlawJLkzOyUgCX
HzrXVt4GRDv/ik+cSYZKG/SzHQ7I3BvsoM858mNrmAlb3sQOzguPew64CbidyMZ85Mw6UsNRXMqP
hjY/USQGz71Jb86m3RxLNwXtX0W/X5w7MAVBOu1N8yJ6GHo/2hJUh+Ewa3yZ2CFdjQ+leW0OxNJa
AfbkkQZIushA9tTsAvCgEKTkpxl0w8DJ4RCd2i0aOzSs7HYVeJUjOMoPgoWzA70egX28Q5Jv2cEN
M3xMDS9N0qDE7oSn0HLoCNafHmc3HLxbdlIBHegKFnz/15HZzbi+LAX3iIy8DcTPvxpmtfiu2Ho1
2R/3pIIeM0ajbsl53lWFR+hHoyzTOHYQWCq1akTMXL+5wt5rIuOU7CuuFzYEkbhrqXZLT7cRzhVS
m3VuTfhfMDtOBOaXT463QUMxhAhc0ZrMIHYeEzi2ZlBiILalNWNfYbWx59kWzxYtzAFNsnSBR3hI
CSnpit6miHn8a9RA1jxYn/33FDYlGVRLcem6ELnAhAR72NMcFci/pVImtUD79x7XxryfiR0XtuKL
rryMUDlRfsjWio2T7HQ5DtXn9metoC4WkCLk9pAzteMJCs4eN82HyfDyp2fCqcaNnW0cdG0pRXCW
UhMVGE1Je5LnbN7Z+5rLaPtZoP6codGJxfVylxbIC5SnPXnQWOAM1cseopI9WKTxpBu+O2YLAMdK
AN+r+0cr8Q5wGLFYyZ2/7Oo+NqhD9zf2jkxzI3j0NKNTo4wVWCzXjWfyre5JZ4jUfXJCuGztbWBY
b1XffsmjB1pdBAlyvxTZHIFLm+d23YkfVs87H4AWegiJc0QFGBvpqc9d3nyFdnphFS9hgYnhwSGd
fGvFikN02HIXWflRcDm1+uJZZ3cpzDzqXZnbSAoQaUfEtJQrW/CWC8fzKwFSNAWs48aQbwObdyqb
hH+KxIwYLxblHF/vWRGwzobkizCcU75oPa48cyzl2VEu6NybpvV+wWfUzNE3FuCkRx5QCYs0W99v
9ygUVFzDzSJLbAuKr4g+5F3M9+l1ZICmHdfDUTxE9zaNojK14L6SEJyvi+0plIS/bCOhVEonBAY1
hMBOzc3Xpg3S8dcEcoftQ1FBWgTmC9N1B2SDU50XQWPQxck21JlwgvlV5i8SjhHjtcuoUeUcwgpj
orcZ+lr9CdlBsNbFdL1w6KLrCMdiVFhpbxyWR8NCn5J1+Ka+ml7meqhWlv5BvZqBVz2oYLACDcCH
TsvOeQnlRTkwLhFdZ6cievLwm6rh8UO95U8TJTIx9rp8kDzRSKqpxAMPcQnwB0VQ6pB8PbDdNCUA
7HgWEBmVU9Ei+dCa5/SNGpoD+TVfVmhs6nCfdR+Oyz0DuoiRcBVS2pny2JM/LuqE5SQKZbmUw/GI
jt2/404HM5RKiG709ZWU86hgcPtVobmiiC76TwXUOUrtY7F6hN9YEvHTUc9Sfs+hsQy1rtk3ubq6
+GYOQMwFQfURcIFBNn77uguvWjwgmnUK5Cu02Ti6ijVZsaURkY9JQoJhbCiCrNoW/P7FbpmPf71f
KE3Ej3QfA5wJ8XXzV92V0Vq2sb/Y2COF/Ik/abxj6O5iYL9OtEWCHVgiQkzUk1cxqnLVDc0OmKUC
/qeVYYlkCw1RB9dwsZ0I2o3riaBLPBzDU8lg4hQ+M52NgWFnnmxKL/ZMpNOWWtrbXklF5uORDB6l
zLIrZq/05giIrtHF5CB3gXO9UIPx5GaYpPC7Fr0T94i9Yk71IFJVJf622NWXVwpC/awb2izoqwtS
ywUQ2dKSLWFgoKdt9AJYB0HVEsCsXi25aEOUNfUKGkxZ0RIzZw2sL27thkcXhdfkOiDM6XSY61yj
Zdno/3EV/TB3moW3IZxbzdpWRzuI0yp50WmNJwbgNywlogvJMkj9TlJJq256vSkjuEKjHaSjxWHs
enVkzNy7Taatrm+nWzc7jYzp3I5vNlpvlyJ7edSMgNAFB/7pyV8VYKQ+UkSYzwYJftWb6cuiheof
O9Z2wfX1hI6ABE0SH41mjx162Dm3SaGV5kx4orttq41wAg5pArhFbzNXjXwKpO1fX8DY873HUrWM
ql6s7+oUxmPTfH7NWQptqBuQMAoDy8XAGon/1Vdv1ltPMSJ6fC2s86LMkfJINndMhX7algGWhwWA
37DjnDPBXLDKCiDWtGy7vQk36MPcqII3s1A3s3y5XwMCwPyio9TbBo2CK27z2edEZwIUXVCIzDFV
giWUkqm6kfwjzyQ2JczNqSW7bVIHWT7snaU6Ty+2AwWKRsgRradYcILlqXKCAOpZIXCNHmhq0Ub7
WlzAB6Yym2bUuVMMV1mJzEIPUrTWIIhfFSWXKkvVBjLqY89Ki4M0dHGwTesMiDPmNOItCIODAz5o
NWCXS7ikG9SQZMoU/rBRtL/bUV7YIj9+l5RQNQ8SXa9CRBWq9/rfcec9VQkvpwCVIO/Zb1bDh7Ki
SYg9RFxHhNSXI1vJLqmUDalutRXVme+twiHDBQvejGuOdIU5D9l9eUJ7SaVX36UuC9wMRXoQsBG5
p3vM2opmbs70IKEM2ZUahGFgGDpXw6HM783dlRSCGZgfmjf93Sk4u47bRlIKgfxuk5r+zDMY7+rr
GgkOQdETFvfWZONmSUUCtwU3NNHghyiW6XGUvGekOKZvEF2LsgU8ZyxB9whzz9cXb/1YzA2rpGgY
/QtgZ7cb0loe9G0/qa1D4SruFTZ9aczQgyG575+7JcPBcJPOBEa8GBQBSq2C6LOGOwlNd2blBuNb
sTPdk0n8TCbcTzJyeXyAaTm4icyOsSBUr8zVdXcStm2wpkenHyhYgiFAr5ljUtACrVcHj1TQXhfe
UjXQ6shye1WPFqCCfiKqDHStGArV0akLoNKtvDjPSeriHasXjE8XlsAsXcb+3ANg5FKhA3g58mVu
nndzN1CGfmOJXqa9Ad5uNzAIWMjVwP5xD/ICAl7kly0Li4eGQFwOEVkRwUmfVLdhOcOrQliijhKN
G6PqHOAeXMDhWSFJMWuBvRFRMpEflYcTxW8Fet8VsqqatMQyaf5zYQEI/t21IM1FMZcec1pONKqP
2cBLh4lS1fybkY24PuOHUyDE3IS1dEQgEUvksatGNhMGOGSRiW6q7os+BBD80pBXjDFkHDOmhAQL
d7RWYkYnAlrAHaQeewsXMfOeNGlZLUKa9dfOtjCDCx3LYvxXGDgKfJmtnpfiv1x31WzV7xkxRiXT
V0HnKImpP2nOcFfaP09f4sdigJqo2xWP8+yXztYD2lYSa7LiWYoIA3f1fRkMI4wuseHzAc4DsuQ1
OHiEdw/SUa4UhlAJ59Bz7qxd/LOmZ1tEGwdss92seF2Mooi8YelSr60QQkWdqlRRod3rsk56UYfd
95R5nIbMd0bmP63gpcfZGmGRUKLTe8igY0U2UW9I7IEx3ZsHvzEmCCZJ1HKT5o9RzpPisARA3Bg7
wcp6jEXFehL9EcolbQeWIjCgDz68zAfjwaTJ1bkIHjWX0kd6lHqQ8d89A9JJzsJPlHIQidRPIJOo
Qrwe9+BINofcKq80O0tYVdG0FA4ZCpAykzk0R+xLvXOWGdQajZQgbqxnya3UxlOXHBtnp7xVHk0h
qCZ2q35Ru1SY9Ukx/Fdihtv2JvmRNQYiyZ6w7dfdryd6aWGH3aHBuCavP3TYSp4lgXbC2cSFcGGP
Zf0SMwyIkPGRWFfg+qCF5NlKRiY5INu/gGCaTBKbFWeNRhdNcKptxhB6GzJRuu3t9Iyr1g+DKjNX
63V+f66gssQvWB7oUn/OBp2LNeXSoYMWrtfmeWLYjBOGDO6I+1ION1foP287y2i0vw2oXVBDsAg8
j1DFn018SpSeqmAdjs6LY4iG8aMs0Il/Smc+ORJQDlG+EcXHimSTB5cOKSPi4itgaEbqwYcORDoj
ZJJnS46wDM3QuvIKtJzcrGke+TWLArI3DcbmAl1SMgjdtOPCHxXpZM9HRGzWp2IGb3Iw516EttWr
f/pEO2H9kvG1pticvYKH8mLXrwELrL5zYC+DGp4+SK7VBajMu70kWb+xtjLX++fYhKJ9PqOFhQ8F
1ultXIVKxkCUSGJdC6Iu90xT3r2y6bD9VDTtx25MDSFhRVYJbA52gTh7dWl+3Mu2MB2nWozbtxXI
4gnZhlA6OhamG++3i69ukvJwkO8trEMH+bolFLjWLRWVrMa97wEYaU894H9kg1hggZqmo0g2et13
5Ai+UuX9yfq4zKFl1Vd0SvRBflkhNdhm/TuHoDWWOr/P5S+QKBE7dnZ/EMkllEMVdhCeuN4Y1z9a
/Mk4GKYsjI129ps6ejxkGf0fkhrdCXS8cpNQ2O2ShZDRe+2VoxzPenkroXjbAD4LVlJL9LZTxdkO
yMxTRalP6ExH39YbIrH8zG/xylA6xvZ8KPRkTllphGwlL8YniYNQkzjszcyNgNSmV5y3TfyK0Vbf
P6LFGk6x21AyZjy3pMwYy0zs9BLJz97yahLhWHmqCSg/J1SFvCyXCqdxxF35gA9t9e93OaGlkjrS
QDRYfwvci0BGh+w17yuWXfv+56SunCJW50gU4lX7NUl0JR5fdEtXrz8nYx9DBilhX8lYnqCUNb2u
aGyPTyCSB6wogBYMYt69RTSGZeTH42dnIQt8isu8TzGzITpupRZqxQcaNSzjjTgP7XFIdimCRgym
IKTNJzbB7qQQk+kts099/LEbn1EuZ4tk2NivXELOskVg8Tw+BSwxE2xQzyZD4mR7onX3m4VNZdm4
xG7PrNNT3vceA01Eu+wNg0IOQ6GNjbGUFa8jz/xZ90NCZH59p7IarDx0EfJuuWhPsiVtkiSgfHtu
dpMJG62I0tIvJhFj6AU4jGtIMAvB+5IfBYT52RzyK/7GyMhY/Pgz9Jd0YsD3mHEXod9q6s+HV5k4
nU/bU6IqvFU4n4ivACdpJheEe1NB1aUq/EX3KAy/2Qw34NKta+BN/s/tuFkKhDIGSQihePRcjdgr
aO2SV5QIbYe594enP8kkCp6rNmcp648ARMyaXH5BAoK856lbHstN9nP8Qvovdru4KIh70opgfX97
nLLERNdg5vljz6blymZZCb/1wKKYzskckOTUx+MlAOZkqeMe2qoK81KSnd3EaM5q4wqf1evPZfmP
dIfMTQoNxlOgPWx45gXLqUq0ZbHV/Ry9w8E+7mZonQhyhjIvJFR6b0ZTmRnEzf3MITYn3YwU0gJG
HMnL78A/KYPyDjYOmq0dE5sMOhXPIWZeBOvw9xyIUF7yqTwpdoYymrsUH4YSxYUFumqmmJdMYLGk
Q5sUZ0cIibt+q/Qg66lthnDbhdhX4gnPeTphP8qjIuyVGe2tlv82dsDqzgrLCrIyE7vSdcjlBiZS
zs9F8oGWFrtMjoSNcOp5arcUlVHStpbZwHuJb09I/Rxz35Ra8lIIZxWas1efgW8RdMMt/aEc4Gii
XvNI3OsaUxvfvyDEgV1uRmduD+yIbVW0kdd3vBxccP94TVBkv77RCHsrdIIJddskBS/BI00YHKcv
UFs0qpKqNwofDBaicAXoG/efPVSL0k87I5aU5uOpxe43CwnXM8Yvh4oNzCQ0DgXchTlzKOpMWyyl
6lpRWNgtiSJBjIa3OTuhqlKaaf5jtqFn8rqcFh6vAFLHpe1zmuaeqdZxI6ROXcHRF+wbzkyMIWf+
rDswd+ypm8k7Q5RAHHoyETC/JvZWCCTgVmg2+wtEBKv68QRqFAXt8Fg8uE6Y6wUVyldRMHizyW3Q
cNIVlIfKyivX7Qu2hrU1A5XRVD+O3NIsRQkgrP0F8jz30qc3RE7P/j6mps2j+RBQ4col1TfQLTFr
qPNccEOvJZECwmEI+CxIuJo54u9CF8oM1gB//8prMTrpA/d8fTGhszqYSp97WWlGNpodrd8sjIeb
Zzd6LTzOhwTCf+VRjYmgj+0frh9txZI094hU9on46Fwh0yb+keQ0WpgNWsQJ+QkzakSQsfviTJFi
6cgSkRBJ6y/4pXkRuF9YWDeE/tiS4ELYnpHt4LiikSygu4/Wq26abiailx3ygSV0ctwkeg1NYchu
UeVG+3KSjkQRQtu1/D0gIUq7yKrlth+65/ehpozkp57+5Yq6x9iSZD8Mqnqq8udlvAqqkrCYJQD6
YKkcVrZScDsLzpitzkB4/eIEvfpZS54xxraLpsyKe4hPmOy3CdFBDOMrKOsBGLL4sNZ9z6ifaQkT
yD47eudNKWZJzI7EwT4kJE4UQiLvoL2drNji1wRhmzLlSx7eXqV/FZudYnKk+6SBdx9B81JggQxF
UCmJm46/JDmCplzjMaMUWzR/HFUGbuNFzoO3snl2aGSE5zQ5gc9xQrL5kJfgjioQsDw/C4QQg5sM
58jDF3ErIMvbjaccZPUur2h8UTFWCt+jBuxKTcmFrLTllN1pdC+nQh9NJUJQazXm3QawVgOqW61l
UQOb1VNpkzORWUuBVi1k2TzLChMYGt6ZbjDhXM2jlzE9bJKLbb7lw/Q3gRpeQ5B8B23nO1tkaZ+p
QGO8ISWxWO9pcwZY6o7WW4bM/bp3yj/HHaBsTCirRGYse9694pQUI8mVl/0GI8AbhT/0kK8lvyMq
Tc5F5QK1Li1pkkNk6+Au2sh1z1ianJdgC86DuNPLGkZY14cFIOjgS6oygHm16FwKgRIRzd8uUz+V
c9wXM5llBsliXfWii6iahDa5ng0g582Oi26UFGksWnx+WrsTdS6am9mP7CfF3jYhaDoR7aTXgzOx
qEYC+w3jp0nEeTjODElwJ5G8QvMKk1YbVp1omHieFAV+1m2Ic16MsrfA0NtutJOPdo90QBgFJxw3
qaEo2oAL3/OCGs8CT/LQaAL+1YMqHCgm2T+3clEHcHRK9ONJHREfkiNnCdJsnTCIDvyH97ccgkMn
zUsEERHJizzLJdBDEBK2wjVsKcouJ/urLV34w7GES82Aj9bake38z+kXssNaxnQJkgiaiwuYcm8s
91S7iLMEWQO2frdCTAYV+LXKlQHjDldHbaTTE+Or1cyKeUYlCnI3PwMRrRldDolUVGGlffVaLlR1
KM5asWQ/7B045fq/k751W3PYaWC4KEwaqvdNf+oJ4UR8YWLvncOjYKgogrlb+GpQ6tZ0FTlT7X5r
tG24nR5oh0LQKQYwWXPFPgPwBTg8/g2kfo81w+Kt09hpmWf/hjgqvkPr7/f2RWuKlloCLPXzAMtZ
dfITU0Q/ODvmS7O5mXIpHxhI606BWLnlYmhFgN0gUL+PJ0OUg+4c/aH7GQcht5MXt+q509MRrobA
9i5CfrhBOHrkrRvpsVWM/ujU9llt2ccyKpXq3KAwKGu2nsJ/U9LWEr0BOykE3tDNwCRjMPexsi9r
C0nM2jI0bYPRsvNNXlWp5Y92vRexWIlEyIlnWKtZu++X/ov9tAXUXoW71Og1q+knlwnZaHU5abvu
G08gCdffURBfW8apsf0uOyNhaZKyKPxOoFH0VgrHHLklWEegRslyDLEELP6uB2QX8+KcbufgyrQB
/tVVo0n00069qkA87hecxjEpHqrW4OslELprgMJoUBHJ5lS4oGqEI5Wbu7Pm5q3WOG6t72ubXYYf
D7DgwQ56jdNNSVzwJgCyRygDG/I05yLlJzjNF9kwh6ivacEjseB9mdlZf6ny6YW9x0f056KC7TIc
wOZ4TP6eNWXdMlSJyDQgNmwqYuY7Kc8g3vC59GA9hGNp+x19QpUIggH9cMccD6a7wY7oqWH+xKqC
9YZjuiRrLOPReH/GfGr20tcC7o6tTdBOO2Uyph/soy90WXpiEP3cbQfGpUQwqMe2bph1ttM60b0h
dlO7c1UZdy+wGtxtUP6IYCBspIUG1KK0w4dYEWQ0GQEIIGf1i1DyrA4toI8HUNGdhxwjFP+sh/p6
8rVblion1lPCQuBJyJm5r/1V0KG6oF1hGg2lNPy/lrRdbXhyRUCIJcJnmPkLkEQHNgHl484jEvi+
UTBaHskbAlc/x6DoAVDVvgy5vxXt+BGN5r48h5vnGfcd9DIL918VSJc5aeEjIY3K/1Xriy6extXt
hkEpVVS9Du2xj14hZpzo5Y4seJN8x9vCx56UMHoqd+PjlCP6om5Lnv4A8BGwOBxgtXrfzK3fB0/p
80bUEqt2OwxenBwehLtJnYEpV8Hqw2UV9Z+R6nGDZCtWZ5QWKujd+r9TP+WI1QfqihDwFW5VwJEB
0iaRLl7TcF14XWjeDh1Z5dNLjgzltLG/195mAvaC68P2VsjjtUC3z4ateWHGhms2hj1N6s4Um+g+
U7XLbDxhzUz2pxbxnOko9BC4B/NvWH+6VLAvP+dpVrCUiQIOtCitYPeKkCtR+jZT1xmQyApj9vre
HCS83kti+3qdhpAB4P2ovyBXjr/1p7SpKCMl2G/2rz5U56A2OCnpG/WFTcGdEIxOwJGXJkkUuOmm
inGSFbFSKDDcXaR5+EjkVYJgHh0sUArTjVFMt4KsvcMQMcGMgL8cp4ulxojRcnsBM+JcylUoarpz
PhbaABg8R+L2RVAXmay08PKc4xJ30B136K00jy46oI8C5ZUWXwaeQaV0YHSIBTlPznnUZ/MOAs6W
s/4CjLsY8F+mx1wfhEWyUz08rnaCOnCW2YN8ZYL3hSPEu1JYEwQ31gy0dAmDT5G33vZR48jhqMeV
U83hOY5k+0DYcEjuc5a6DXp7+bRtfca4fXIjWaAYpeUJyaQvG5K7WWOddGIH88o0HjbOgC3AZaHH
VSRbm73ub45NJuZIRmhdi+xWD8ExrWDDGToFBlAPdVoA5FTfoGIdqW+18NlELRMTORZ5j4ll+yNa
fWuhlm8KkNnZDMB/Qe+Cz5u0EshSTUb0AmYV5/30R/CV6CQ1gwe8B/ib4iZQzQcEbMnn8bQm7SD5
jF+dmYq+FMj87BfLp43/aaCAP2v75RKgQKbpSam9XsNGhdOW3uj7N8WfxM1KUc0xszSi/Syyz0ZR
qExEEJGMfhj6cpZZlOoa9X86g9SU2CWj8lK0cRa6XJCGjnRe+X4GaJK29Q/hKV1LCpPkQvpUEoDR
18fW583XEHIWEzDNNNluyv4J/sy+TIY56p66WfNPUDZDl6NSRLXXRF5r5OrZ4RnueftavTfnbaza
X6mxcx3ko78bU3VavNdOLORu+NASg9DuwMRt8zekM+ir2Z1E8Ng8/d28GeRCucEljI98Oaz4rzVS
LvGIATO5ZlmqXw5meGe+iZrQO3XqxeTWzlzPYSFR9tyRcMxoquEK6GZQs9Z4usUlFa+K8FQuYopN
25tMoRp4LEyTCq/eYC+tXRPuWd9Q2C9ERGRp+mJimaqH6B8QXJpwNBma6IRBmoMkg4Dw65PURIcU
k66aXJpAN4wQ5PEt1/+YCx1sXORY9WSwBuvG92JYwn1Pqs88E0k70MGYUQC7WZWmXv/8DH6WvhGt
ZpZ6Fi1k6vk4BCW5OM9m9KqJ697JUnj1MIX/k8DEKTELfvYVT7tY8AwPN4lz0IDC4L21kYxPyLrb
GDa2pDl1W1ObWHi9bWF2tipOHfSMvijDQoYh8amJRwW7vSLJtIV9AtwQ2UJUZF1s7iUe9wbqG3BK
VMaLXg8CCTXWtb8mTA3yJ7kOi/2f24nTsDcV17mYZgepYHsnx27+K5LCqsuQynkx/J74eH0xUwJm
cKzXT5arcz/3ob2CI7bW4iqLddfBJuY6R3H6ufJw8Zq7bx4ryAvyhGFecDAfcXlmlF/bdYYzBf02
L9yH/4ckIQ06KtX3OpkcvisxXCCQ0O88E+mk0++lZgzFehtNV4o6SHBqXuc96Au4wf1p2C/iqpw8
jLtyr0KFV5a7oDc9TITgeUGZEi8ZD5S023vVsHzK1Q72sQNWWjehvtMJxnjTTMuo/xplCMMSXMUh
NfMK0se6wnwDmmHG7qC0pJVI1/8i68hDz4Is0IXajtk3X+N8KoQHwr5RA3Oe6UDLH5o+am7Ob+jo
FkmZ/0U3D1W4kXm3a3CAZ+ALy92n3AVYxjdIOsYUXb9kYQIgfuDGvE03rp09bvPby0KLkQgEliRB
uDAAjQiMbsD6/xzqTS0ADpYp3AXRmjm9ord/UccRsxjAwON0R4+wiXCrGpyTMGN4pwf+4PQ15dJP
tIc2LA7I+mCua1eVn1Ml0ywprFqpKjWA9bjnvvQhOG+avX4pdKfh04SYv4r92RiWxtoJnhdGVzWR
Mvy3iJMn/7kf+TVdOsVx5Bra1dVimKxZRssHHb0OY3IAj0NA5b14dtlikcq8OOoP1omHf2C/7LYL
/QuHqesCXPwGgPDeuvHNIBYZFJYiihgOSMfET22qxtZb0+ic8TFi6cVLqCHAJzhCwbs/4WjPGsFz
/8RMlW12eKZiWdIVhfGLCTMqHxNZycAxofI+HA1Za6xpulYSw59oWRFFAAjiK6qgzKjRtOJk319d
pSqRG2i+5J8Pzvow96I0lD7YcTG/xco44DgDQNSyk9acQSiGpxCgvkN3Lf5K30yKGTT+jYkSZnNf
S6BGEEUVBKz7nZsWy6C2EeIYzOIBd3TSyT2kI3TToYIPlrMgf+d6hoUp0675j9s585MR90Je9J9h
xXLGWpzjjbsd+Cw/47BbkanQ9oIaZ2KK7aeHM+HGmRwQN5FLJH6PSz22MQ/4nbFD8FLR5hxAvDnM
u9SD187hankmhm90RJZABzUNnLqQDQR7b+ZlGlq1d5o8CmHTzYO5M9A9JM9bR2nHRQf8dWX7oWAa
8fQsvkXzEmvxJI9Cl6OyfoCqDPfM0t74oNFSbt1gzLxcfEdfSASbBJwHAOtRfSzATfRDlRXpQfQ8
ukRNKLL35gAQEe5ZBBT6npM+fsiTlWjOt+awE4TV4ELQVLXEDz70usmnY6Dja5M/bpmlFX4A47m6
pjU53EOD6KHehvSsq5O0q0CaAWl2ZoOFFhJxZjaPajBLbN6BteH5/RTxK5ArE/tgGydQXQfVViqz
Q8wsYJ0NJAlPuKYyA0BMLwaoG3TZOKy5Fs6Yffx2gfsd7hgeuPtQiLdkwpxmmCCfp0ABgtgVoBUh
gIILeBcrIEwgWlAMK31YfOnlNO75IlJZWL+r9syE/YrPrhc0GByAjlv3UeX80hnDNOlSzvuAlBt0
INvOqHWQX4Tw9SpZbOBHk3BQyVwOgFOFixFDGwLtt6WI/Qa75QPwue3qdPXsG7Baq65O+aZX3bwv
IxRGWSf8/gSxNaoK+7l5vyYMBVGX67aR0OqjFNYO+d5o9cBxbJuSm0kpJ2F11+leKL4a9Toxr7F7
wqsx3ncXKgWqjfKG1x/OBcfV91AQsaeaTGzpMCjLq4Ca0itAieKBnsfLEGhuqElBnwODSTRe+g4N
2rVnquZk6Vmvtq/Q8BtIjL/WF3ULIX1WwBh1xuHzQZhC7++hbyLhaxl2dg80YLVmecs1BXvPUtiB
tnEoXbVxi7XgUOdGV7mdQ6KKK+OM2iRLNeK3hewp3HIdeMKByfpyn5abzKLae0yuW04toC8BwEcF
JgX9qmQp6JE5WXE96/FkwG6pQtr336rowGg8V0GMj5tctvGuSrHs/TBIm37ltIQqnmSqgEihja8k
eKu5V5Pz0QSUzLHKh3/SU+74GKpb1vLm13TzD0ACUlbopZlU6307NIFDMfLDmRKLPFrgiBku1NsL
x0sNTXEFgcTB+i8T8hIiMneBWvyWexegF/GSYhZ3aqwB55KQvVIVZKALTPKq4EvJ7R686HaOSDAC
9oSmaQa5/iY0TWyZfiyOhMBN7GzSw/xZ/eEPB0NRaGjjNSUxSY4XQEcBw/mSD3IW5sSme/lrUXya
5Kn75dp7tGk96ChvCnY/zFD878cEBT2DYRMvDgBScF8NEq95rXqNPjsjZ6iiicxnkeVQT1+KB0fM
HGjz+sBPZkGxNiOv6jKzmxAQ2C6lmQDyOuAAWcJlC598nqveDu+vQ5WWh5hDzKgZv/e0KI1JsAjw
eb6HXOUASWQrr0Wz9BVhejL0voD9feq1whXaXIxapE15xOMy0fym8w3813Ni0Q5KbMaPh5sNOLzZ
Is3XrE5MH9aMq5ZGL6BVQUTo1tpmVAHxuVmBTZlXQc7kDHGz4RpOGzgwnL8RahudLTnw86AxF7L5
6MlqTKe/KEs16QnZIobADKBwZ9UohH/t0Qya6BMaftWZsI8wd1c3f9Th+/NZoVb1g2Yld0ir7dek
lo8DC1wOBUf2nCSUoBuXwTgThN26Y9WF8Ad7QXx8c9eFYHY7xfYntT68o9SxyZiawm+xwPjXwRs2
UceKxd+clrnIoAvKr6th++DzqFCQ7FC7Gok9m59fPdKwGFgHsqK4WuUwafofb9re0P6FIY2FNd+a
0k6KgIjEVHqsa5P/IVHUOWiVmjwI2zxEVvGbTF/CotvoyZkLYdsO5iR6tWUvMbrc+hClAaRKtH6u
ybl2oQNzrNIEm7ypkwlPp/A51DxIr6yk4p8e+0T1TWR9U6wSBXQNfQ6IN8UDa0Joqk5bTC+g/cla
mWQZwjGzNagoV4fLJvsUMscGpjbwqn3H8tBhjiWqkY3kUhOc0mGeUH0TbZlbK3SYA7eyz8DgnCj7
X7qMuiWpOGKr62/U6sZheiLiLdlNWybONPe2qgbfEwzgHyrfPOfF3KUe/xFNNwX0y1EmXl7h3Bjl
5dAcP34VELmc5K7CUxU3Z5G41x0uM4M/y+w44NtYU5hbTj5XUQfZFyAJHldd7lJ6H6W4gnLZOp/9
AIFbNGnOC7m2UsRai3ILWHfbSnQcplgKgV8y5uFZNZA8tDuf70WYHbGMkcOQg+SpuVygOm4QhTyT
rEEF3YdLU2HVvGQQGKS5UbW7Xnq9lZInOUMOokyzsMbHUT3ZSRHicVan8+tH9BJ/rHELfHqq/VXS
Wo6l/3V56uHOzVfGJSkQCbdw7g5g4U7TP/4Yle8eIUHxMa/rSdaSNnO6MgiEWWVah/TT74oFLZIW
DhJgtEX5BxPBSnftKVfVJetJ99SxIqERzt1jnMbGBvb+QDSkLG+alnvx6Kelm9rHZ3NiikS0gooy
eEbI8yrYtaw/aydw8JQZbFw3gC/KI3Cu+BFuAb8f4lrKESkTRHh1dXKBCrV2i/1PJwcdyKD2NFbE
dJb92riXThmhwRT6MnsEshtuZpJ87zAU32HYK3NeFzeADz3izVk4RstVmEysWFRx4NIVi0/8FFYf
5NJMiTSkEvGWjXMs8dnpGG2bIwu4aU9RmYHruN5NRAcnt2L8TnDkFzp25M1yhhOBEKDY1Z9hBhHS
Q87OtviRLVJMcJjIgA3fC0m4W8W2vOF1lwXqGn9Gvnvg/jhMmde5OdbRSVbSbazd1mmFMjSjzkEq
f3k/lzieYZZYkIPBNJDkkaC/wEVowEQ8jkcnmMxeTaxWEaIgZ8tSJ6lX1uV8kf4ceJpk47qrUxlw
y7DyCILx7AyJhdfzdz4DJN9g3+OHVwbIFYk+VDEQwIOjaHBeNKLTZKEDqtKV85FbfCsNIjK4YgUn
cLKq8nFT4H4ysKvI5gTKCjiJchjY2NAkUYt+trLuNCP/fre9eoC6Xec+1b4jj8Ik8vB6fTWO9Zvh
ORmsHgGoHQyzZOXb+KWvHUB9nvQ4i+xMKNh0coTPJF/0hpHx8ehMAWh1wAzTvrGmRDAMUFcdeeI0
gR7N/0B3ciDgfqGTfR5mm+2/04JL5YaJgWWhJIoQwsNCCVvgBzAHTcmadGT/9VjgX9COxouVqUp8
hppV47IEjGx2kTUktJPJWa6biSKjxsLHVDm8DTkfP6DRfU9yOEzdeo+C52VcylOb6aqZT+9oM6Kl
pKcx/fS9f+GKq7rRrhLc3uS6IKV2dyVmmW1kgSisOyoqvCeEdbvQwteGy3/UUvfds3GNIOlgvmM/
qgxCykIWVnjcCKgcn5o9WpGHHZ6f2OZ2a2+cNGdUrFqzpouBU1M3ZdjBVnAFQj4Nvi1dHmKl0A9i
QYyOQ/4VQGhtsGrZyI42SO0YOs7NUQV5TLVXbbOXQv6qw5uhis8A2lDA/mbyehVwq27Ti7q81p8Z
hzYa7w6rhkhIuXTkdqXn9Xy58XORF/J/slKS7MLWNceW00bpd1iZnuXKSKciMeRVIGEW9HpClv3O
gSkToJb6z6kQBS0Lv+wWKTGtlPgslpggfGzDdHHm2tpPzSZ6I2FBin7HYox0MDLYnJddEaduFYUb
uUWpdHq0ZZt34xgo/Sg2LjnV/T1ISVgozmHKjje/zXC3QSLDKnXv5JcCour6xV1A/56LKHASbeti
LqGh8Do1fn9zKl0nAHir/oGYb03CXJeJPPkywdJpcRvnIuQQZPYJ47mm8/APlwz+F1AF3BRwQCOs
yID6HKQS4xoC0nCcnxrWP0wLLSZlq4WFk3b6Ld19yrvua71xOKPuhI7SjoI9gWDW+GZ6tNwEPpdL
xwxNC3TbQxqWDD5RE5b5Bjt5JO+og/vYzfKPDdJughdhu0slf2uoTJynL4Kdcylc+MG3j8hNMLzk
bTf+2ZXNBgXyuxlTU311e/Im2pgEKcSJGuSqZLjLdjKhSqHefiaDWU9iXlJQYaT466faC2b8dHRH
VRnc62h4jhmV6/rMQe99twDmAv3/57pNnwr5S2boRAMl80JpVZ99wvVk8QYP7sKzmYmaTVADudI8
Dm6jH0xmvBYIP5s5/P2zEz6I2FIb4oVq+w3SwqNFj7qpNW0iX/1t77DCUczQgcdmJnVTwlRa0as6
07IFtpLEBadfLO+15+GTb0frhqiHst4ChawHs0hGWUTuNPy7H0C/VE6I09PKR9AEmbGqaomVgN/I
xBhKwCWMuu/XrscUoqI8FoJwdDJhVHTa0ZMYu6SE7RXtpfQb/npKx4DVjN0lBW1Qmhs5vyc5ci+M
nsBbBAg1dOG4yB2Idoj4oqJy7WLaXg5JcEe7SwMa5uyB3JSGRTbUnZzvj51t9Y1AdSflfYKh5RBZ
0a0hPpiz032ndr92vkWztaFE8nDrn+R4H2Sygsx7ynmAdw0mQ5sL6JWkEubgBp0Sc6wkXCKQC1L/
H8z2Jskyp9HyNCSuFrWY0rbvSVYOc/sPP17LY9M5hnRLd9HWLK8p0AkP/pdnhiqArrSlzuGZspR3
z0rJbFA72eQyzc8GgDeQ9fPkctQ8v7cqYAeddTtpzPAjab9fhOZMbp9vhSMpJFfwXhbG/k8iMqKW
UV8W7ziYBAOBkIS3beA3KpdpsMvlzBP6SeuMgZFOcmmU6mWob1eYqzAX5hgyfie+lOYV2FboGQo8
zXZG7rmPliulg1y1/NscI3HD9J+p8OBo0Km/looyEiPTwe8HdiUmVC/CYjIbdhwE0m4NURzKtMwd
pDH1uQHa7+lgod+1I5bSVostjz9DnFSFhcA8JeI4Ly2knaBFYQPFRyq4Ho5GUTz/iZpfOfDGJXu8
Lz9SKpIQZ2m9jav08PKNWHM+PwBhXF2IGBIeSdWMKSx44FJeCTwxMQwTSbto4NBgPK3tTQY3cK8N
W6mcT9hVwVhwargkkOCtCaXg3AxTiSz+OVCpIsIvymsU/LnFkevUQU+siHJIZs7dxMy57NIca4Nr
qmxwK0L/Jobnq1GnWewZZy4kqTrufDQMIrQn+81rHttCj+D5Qh9VImYC7RbMZTDRjBmef5q/erbG
wX1wFpDt5TGXuK3isijmQr0E7+jMKZr3yS0o2df3J9kPF8ANcOoYgplljpLH4zy8BF8XztHo5tWH
qmiU1on9M8UH891yKJY8Nxwz2XguKigZJuoOchBc9mR1b4O745BxU/uX+MxarFxQi8bIPMP9CBO2
kbjttzdNDwe1TsBwZVn0ZhEJQ3wYFjL60A5SrG8R2mQg8hKrKEtxpJtZZDEEuE3ICk/j/ejGBNW/
83IKuZ6yZtGXAzGAbgGPp6zuiQXgY8K3G87MLLgqcZhSDMN2EeZEyL5L+0X1DnQp9HKqZroM0SPI
C97ZpreVlKT+21ZhDdstJSXBM5YrkNzO0s+l59UHLJpLbwmQ+EKQhZhcKPfa4q6HtHAKTDCcMFgj
Pc2lFIpOujiPJEDmwDR6MNATyPEr+NcUbdxqpLIeDnqBh0F01dqiqoZfRDmt6hmFBkGlE7fvi60K
SNJKpaO2CksNtK+ydICjAhYOPNl9f3NhlepAfGydxLR4lUmtRSLVHwaMMCQDLK8s/Xfta7izYYMo
05lj87dhbrSM+Qk+MQX+PlKeWx9CqI2g8xPIJldi2S1RnYuj1P8DQetMrcW1baHQg9CaOiWXA7aZ
lHOUT2FLnNkC3PdRYP0ioFAEn9YvlIoFphfgYPauIOPj0HF7O2h0Xaw00u6MbGs3Se4/EkEJiZD8
bXEsffDiNvEi/cTqCVZfo9Jzo1mqRFQO7P3LwYSqxmK6S6q/R6yjTVeNtlXBYDreL8h4fMnD/ra5
Ss0Uorl0Bi1J87RI/ZZ3C6aNT1YHVrPXeB2VWqC0JiCXQOvZzGIHcUToucc7tdP2rCBw5faXUaTW
CzeKSjZA8k4nqB5rmeuHlorHQUEq+DsGF9fztuuVEM+RTkM9WBGGIv+9I/OQEEVpWw3R+wqq7lLN
dOMv88yGVaEZKmi4jqnvXAhZR4YqoFzyKuZLzzEPzq0VGfAz7zDhzPcCUqSYhQQ5ViZg7txWYdb5
8V3+Wlk8D+ZHkpghJsJBGwAd4MLATO9TzgtDq9qWFozNTflmstP96MzarPOIU/z8oqXnIPI0iqqs
5cJ2dTDesGxi7K2KsfYLoYlPHg0m+w49gAan9kw12AGfi7M2Z0H6tR2KZgUDRG8jIt5utqpqeq1B
Bndjf+aitP8QyIlAo85EkTE+CPzyBWK1m2Uum5ujV6VjNPrXnDJrqPCesyioM8bje1UImkd6vF22
IMXWJUVGlX+pmJF3xqCT1g+JYVangsuhqFm2zxqu5riiFPHnVIUdr1spoTc2cma8wOognkjphn4y
S31/F1j2TQ8bZ2JVpwiahuM052LOCefV0JlTPTvtvFwOh4xxdiBqOAIRUzPg3NUuoQih9NT4HDRH
oN2mdjWu/IYVyk+PKhHkEuEgoG2z0YxVPHYJ4+H5qvG1lo4MchN+Sda/IJZzyT3uSlzx4rBmco/O
nii4w2QvmS9qVWYQZ3kOZ6iYZUG4VajY0HysL3K/NkvVAHy6NNlFs/9kW2tZAu2kZioF+Hcj+Gsc
JRXn1RdcPMYm3Jb6DziyOl12KT5QJ/4rhR5vlfNgXo5/i/4QOo1qypa6TVma5f6IQ9ztXbNTd73Y
XAwy3esbVfzjD9CK2yv30jnLid350wr2diONQ5KS7rv3LtzrGFyTLvvS2RtHNz5HtvjSRZnunBPB
Ti84tgnCZxOCS4KVAs71hlX2iQ99A+aevuuCWMnvlvHUn7ykMnDgybvT152HoBgO0jpUp/H3fdGu
Tmx+gs4sjfWiEjD/cFUFlMSc1Mz6k3P2ojXe+vSTNoWqBLbyrIMI/wXBONusm6JohxKNCJFah4cz
MbNmGS9cmUb9daTq4+2hW0WwYxMCdN7DprlNTJVetfb/eOWrHC85OmyEfyA7dkLUU00Wa5kRRuSQ
BlLI2R/YBrjpSvkJnrecVOCqIFCvVSgQoeIOeQItDc4s7S/S9w+8pgUwMCSLDpPAjgjvP7ZPxIkJ
FMS04rU7dWM2fgQAGl38G5yW3BL7GvKjbABJwIUgV1sxyM5lc0NrIZWKo2HcbeV1Ys5WpTF9Mm6X
+OhEht0Z5rcitYi2vyGTKKWrRZr8OP0Y/Dcxb52AkaQdKc8N5pii6bNu6SnkuDokbzMNWw7D9tua
qgumRUpb2QWttZxJkhko/+d0QrPxkvuSLgLFShBuv8aRT7Zb7sE2XavFYIwe7my0a7/dunYrAjti
2mx1jKK4tXBrMJnHZDTfvtqy3RelF/9JKC5Nr4EWpK+y4qyda4P1+GWHveeZzdJVLgWjFLhjI3mA
GOv9L/wLtsYPxcD0RgNi5nWSN10/vgc3NznSMyb1boVtBIm+6YL7vNO6EIRpfPYeTS1tMrgki9XE
/KicqzIQIY6HUNifLlGOnglSUuY3mxJR+kNUmPtwwCsdCyt/7Mjjj9g8X9xVwCoIkCL1WqaYo28g
bOQZG5eQDWUOjE2Mc5umyCKRtyPzOB7Pf5xG4T+QDVHtRUmfiCLm+ZlTVeI7JP5yCsEM7eWO03cg
BI885t8xZqMQUl66LQZ+Gg0O467ncbeDv4/5NS6sc/7LY6hUmch51/+jb6JWbpRVWtKUWhqbqzfj
SR0KgkKXz5RCsG7RKc9iiaVKhUHG3r1Px1278yT33hS0mWNoj3JgC6asYRI0P863GhNBdzPORomG
oezdrTKwJ6jl1cDprxzW3MS7fSRB3YYNneHQa8SvCRhGIaX5Q8Mpo1jQ1imYustWR4a65uy76MLZ
/gr6O4vwWQb8FvAUlwGMrWy1PgHmWar4B3L7X/pnuKARYMl4cuexaImbVubLUg+vFNm8pqRq7WwB
sK+SeqAZeeVed5MenWUzdMDZVQt+gaXfa3sPpt2ig/pQ9Gmg4QYKhhHZ25+vi7H0zCD+6F1aUsmS
j8J5uzefmfTzNcFb2bIOyuEvGrV6kZzmT0izY3T3h2z+9umMzMEaJWZ3/+UKCKja//TP/69UWRK5
OceD11ynGJ9II/iip8MxJBYvGhrtRy819yUKq+A0P9HxVbe6iJsxBtw16ULlf2KxfVsOE0lsoFRW
vs5SFC7tyr2dJ0SVjP13P01lSkhaoNtDZnvf3Wqb+fBMLFcNtw7XXlGKIUbeQz07dSOYoSGxy531
FYCzJa2DDLbHvx0yVNHcG3Jo3Oe+JqCfccs4pa2xId/5b4ossBWlguFdQR7KqwXK9REXVfXxlHhj
KVxEO1DH1h6kzJTJrWvTiHbpumKAzyoDsWPJIHlwKzGzhg6dPLakwZOQpWPv/EHlwrCLNMlW+uBW
P22OWZAlAmGsZ3zWjY4cfixTgvDImZhdOfkQel//RxvsxntWTQ6n/CAzakFwR+4az+Wn/su1x0tc
fmP8yex7XI26AOOm6pagZbzb8PdOgnogu2y9JmzSMtHRf+FYywR0vZ828k3A97msNAbJ8m5WJusx
tUOBHQnNco2ebo1AHRHVGmvsc+DRME7yuS8fu/dphkvRUwgHf1nDUyhVHdnAJVr8c1fwCuAxLauW
FXrhTJZJydecCvjS0p2S4Yw0uZmDqnKdEO0Le6ZJfOKNb0Z0ZMLNR9BXTJ3OBkMa/WHxMOcyNv+5
tt8tMFN+8WJdsX60m8NwMzszZCcJR45w04i07Y290PiAYirk5uMXALCTVQRkUWiQh7IuyTwKUozw
pYUriSaUXwiCyHGOJFhxUyOhBi/uJQHLa7M47BqzmbiiZGXsEIgoYUxDzgM6nCQiW2I56jR+GwHQ
S2/d/h2D7RjpQWoa7mBn5CuXf/hGfGjN8yoh6w7g5hNsV/UeDNFPtsqOClg3GKob2rLE3puCz4Fm
fF8NMUzQITd1y9oeIalOQm9AwnjiDbAivYDJD7kjyt/k4vVTlIEGP4l30vD/ouN1cl07ApLAR+pw
Ok+l+YELIbBg1LXX6KE6R496NFwYi6gFpVxZLAPHCu+8sAu3kDEjJzAqxNt1/k7lJM7GysDVJifu
1+mP9/L7jGm2upLEV1ME5Zv2vFbTvGjJn/8DsPFA5yLcKxiioT32txcFeo4f9+CDwuqVA2m6tgSH
e6mObXT3P2zOk/zV8OageddMv1sVZGWRg2ZfKv3x+Idln4eBKog5zPxxLZwDalqDuyOaWZfv1BU+
Amwhku5aD8/EVXgRjs1cQMytRwW+R4QoIyCGCO/s00l6dCM9bjehA9/KeGdYbeINTRicIX1EDbXP
6EpZYWhFC3M6SJK4393p/vT19vOaTQmodh3pFxUg+O0HIsaleeMjc5HWIAsQhC+6scrvoMFvH87/
hqZ4um/l1TQ9Ks2djJa7U65lVZY+3I9sUWAqrJguwuA68iIBew4foXUvpnhmIW1n97yLIU1mXYrh
KFU6FfgSLiSoAcEDJmkTwR+XNoaoTAtett0V8eMOKXEvZAV1QDl7H3wSz0mmUKgKq44/rS0har26
A+JILTLKC/BRIsr1To58+fqdUrusrIBlQQaiwOs+yjHaKHmyjl20Xnz2GMloh42XaAnsAjvgUyQA
fFtYYxn/p/9p+HGgnGdUGz2pFOHrGyiqg+5ygdDo23rswZhpeRGYcUFLo75qSGfe5tXvDdjVSPA/
8Vip90B/fUkfTS7gdaBMVXxrJW3aH31UvOR+1fF3sdEhTriCOzNN/XJLXSV8mUEP7oPFYIEGHf5Q
7/eDVh3dT08SzR+2ML11axSHLpzTNlkP3AKNsxPk5v5pa/UJb7q4ZtFNSyR8xGVB4hYokvZHA+OE
Ww+RhJj+URn0a2CtQv/auUoeOAEgavoE7C0UgBDyUZAMHndEKi0OuaMb918YGzziCzIRo8rLmMkK
/Gn+O+43PfbsuzANzVGQUJ9QldZWs3gomgwYekWRYp9Dl4GubtrtOd2TjD6EOB2/qGiu8Hq5xa5b
Oa3xbhOlBg0xr3PVSsWOnzAdK6muHZo/0Wy2G6BnNR+WccwtwbxwFmpQUhKH2tqP7zuldgJ+fckP
wGf74mJH5RYWNbE+bv8CMgzNvRHZiIUZzMlGwKieE8aN5RcAhuWh/w1RjQGJkvbSO/2NvfmjNsSH
3kwgYM6Aw0zV74HJeHu2yg5gwEQnRul/BRKzPgjH3shnFZaXJv1QhA4n84wYK/MxxUIg6ttIP5w8
+hldSOr5AjjkQ/+UDmHcFxEe6koHkkLEVFuXWJSEcn7dNVM02a9xkRdzRIvK7EurUWHZmkiy/TYQ
2ERsIK+51p1xCoekKztUrgzcFGycnoZr3d0kCH/wGptaskZ6dQmFrl0iluzwOD4KZpDrYRL3Fq++
IHRyxmE2MgR3C3Yu7Rqi7P1U/ecB3A3jme6NrK+o66uOmHssgzK3VUro730i0JZxcs2jC768pi9O
whp2IK34CeeyB9V7T61JvWyuEVhBCfIspcqFDnh4lHRCTKcGn24rYEYJVSQbNu3smObUqam9Ik7L
zh2Mjf7iDJp9bzqh5Lnife5whPmHxJUnk0U1enPvuP4jVMb958LXR2eRTtolPceW5WEwz0uFKZSE
YAWY7RYP+uEHltbabfGLiYcaRIzvymwAYurLRMTwSRbAz6jXdJFHOlEcIyh4FeAUQCLMSuLgpnYn
M/OlgARFFAouFSzz9gfInasuSTTRD/LTA8hZYCrw9TKgBBwt7bSeWnpN37JNQP7uZWDSll57qXwr
5UT4EI4OP4lZyZWmZq7wcCN+AvuBfi2F+X/NozbJWUfe5JKarnPBfMezoeZfRl1KW9UyCYq4N5uX
DhMKt8wxZtcK8aiIyTKJopimGWQhz8yx4ih1GA+SnjpK4LBQ4j6NpoxcSF9YMpnJXhULPKyA+q09
lD10O60Ll1syxFn9VkSArBwU3TVlUJfbgHH08L5lDVhUsuXL74rDwXEnXVZuKwLvaCyL/BmtC3xj
Al5hkEmHKa2EtJ0N3m3YiYFBvGUEWGZEncFfZnNP88pwd1J/Vp2UEFzx/kNFTGIqOAa71i7egslO
cURukKYZLz0rX2pX3C0YrghYqEQK5UjmRrnZRq8VbClXPQmAGoUIEiYHTa6+niOCSuZl7cu1CgsS
EKCdgBE1W5q57+ShdSVOJA1M87t3XdaG+hK2omjTfHxWmJ9pYkc87/O9a0TZOnudQ/DwUlUtNXV8
KMlquENiILdDvGau62h8SXQmTAaJYWg+jSPHmuYr6d9HgJ013wc48vZrcnHDMHw/lDUm0pts7p7w
hEDWQZcBrMOhV12bUnBzVyPbABeCetZ713UqZ5l4JXriFqJCBEt0FGlNt99WqMr5fu/O280jm+Z8
2trxFDSZWEE9/ru8/NgoCo607LgpLHpUf3yIuLOI/upAe2I72oGXP83Xgnkm/JUcWmYneFhx4Kw8
rqzPK3ShaeOl9470OkuaAm5oU27KzGhR20b4o7fzIyWGLIIxJhlpwLLdCmI2AmyF5qvE5NzcoKq2
7t5CMwzBmjwglsG4Dfjb0LDK7/yw1Upo/0EFUi/oQJ9MoBlQGgdxQYScZhAtRBz3ebZNAD2jOmqu
XvQaxxHCF7pzwmY/nx9MH7L97QqS/FoTkkhsWROYFjqT5UIVvfWNXaZtBuZIarOZFv9BgVPuT/zq
sS2fATE6a+SeJOA9mTDZ3N+81DlR4256gMdR13hm5j2JL6dkhtbTQIKc/psxCqu3OxqRVxMAy+yM
7zTlHhVxPvIkE156Qa937U0VEmsvyreEadggyTLxnpwolHk69c3zjX3ApVUVtLSsp6ldv6M8lF7o
uNzKlg14f0Y3scqcs1modmqZyRsDiBwTM6RMHAkV5MNvmGTg9uxRy8iGSNh5jDK2LrHM1T6TuMA/
D7w0d1v/f8OKw6De//IGoZtLIIVeTArwbKSB65vY3JfA9fDPNDWgXexiNq8ayevpUB3Tfr/8Zhrd
sAKPW1IL1J2TrUrkTaOrjt81nAPOzZS4liryao/HvQkji3hV2Z1GphigD6h+S+x57OA59/FNHPlK
sKjGh/dU+42XUY8/3Viz4V6ajWe+0YmpDlcpDsF3erMQf5fUDoUwKihL0l36k6v35oME0geQ7ULM
+ZOmCSU8LKqDwkVaqveVDFAFRs5mnyPZzVNuK3vNjBwI7Va+YMWrLDFZaZFvB7l/KZrnD/gIS8Vo
tdlmVqurNH+9JrgCFKEmPQg5HHkQ5DZx8dktbaD3WUEjiJJJsbqmCFRRFX+uFrhkamoiMHmzpwRN
RxpHL1Ye8atehfjl6gdyvrkokUvOskHOKGpFvCjfCjok/eUw+D4afbJ0dfE0q6aPWNL2oDz/RmHc
jNYr/K1JLNUAZOATTnVNMwkG3zRjmOGUvDkMxQ1dgqkp3Aq7IdRD2Tnw44LqKepCBMPxuBvIKAQ1
7FwxcvEQgdw+Dkitx8eHbDzvR8NxKVC0Z0cMLioivNZJyUk9pf6RNI4Ycm7TG0FwBXkgYnxeCco2
4wYBQmsqAbFRFafd0nMMMM0relbRhgRPMdUMWnV0KMYc55cjVH6yWG5NW/wt3JB83xq3/FA68C5O
LCJo2QyXnI9y1jw9Njl1JFz91KMIDXCwj4K8GNSXPlZh/mECrcjIHwKVXSxYtLc0iLB+1P8Are0j
6Ds1bpyFLXtjPlhbkkThsmFNX2jx6xgDCoS5mtdncs+LiVCsmx1EVFczSiRxyd6QlQli61KKoC9R
IdmLncYJ9qRFAXWd3RIhQJiZixQKNGyKjUcu1aZTJjY6XQBCanhcKPSWVCi4rcFnS2n3u1rYFaHF
gBxz4gUwYqjAM1RrrxiV3KN4KNSNu6vuWVejujBsrwdb797oBT6jmMPcVuInJ6VeGokFdD+YfPAY
lbycT4dS0P+fCzw6AsErs7BzE2WIFLyFcjIUDTZPkUl8ZFJ407wYgCKgTDqP+FhMytWQtN38+VuU
1Zp7n+QGIDfOiEkQmKULPxC11yBXOiy/IH4T8waBIdIDvPyKid31GwNFGRGOyA55JtrM57+95y2w
47l/6DZ9rLJqE2XA7gcs45xpcm7OUN5Vth7rXMX3gj2IcDC6KfWcBVYGcz5Ol4L5g6Ck0KgetwVH
yVHpi39ZjkBK+l5/QhXObk12hZTZDRu1H199aWbNZneCbFN5eiSr6IqYxjQ79Y7KWvSlweV8UT4+
NaupMYA4mmi4alpNoyUGxs2npetX+ZUBgFYfdXp9LBZ11BpgM+7C314d/nmda3yAnJaY6MBO5uyn
s4uzvK+uMACU/teW+WB81iJKZYs8xJKNmpzXPMBKFYuctqCAUPm61TxBtjWzfrPvVJJUCYww6SoG
9gLTBBLomYQFo3oliHdhzT9GPhQCUK9OLfdEKHJ/nYMXw9mTfoiG7OB12bGqhpSenvm3PlEbmFYm
Y3TTx4Sm/F/fGrzIJ8wE9LflBJihwJDkBk+Z0TqUIztlwgIxbWGVxkXYI/c6kG4j3Bus101VyuKd
tzvvtuahAvUwg2CMj1xZYa5wH54/JGu1n4XCpLBn2s08oj7nFbTuf893kwB1+fdyK9VclM6Au8x4
n/Y49UWzJc5/RQb6OiADvoq3pxNG9rUDOOb0RQ6nkl1Abb8ii++uuxkerA8w4Z2aytm3Ex2HsXwq
Kz+OXdvBtjnrQR3SevHxFLznVOfUEPMZjTaDsHhKEXQwkCk+80PHap93BLI/b0VtBqoof4waE+qW
GaK4dXxD6P4JVHULkHD5dm7k/wzv1pA7cgfjy8GwG+zlhM1AT/O+cGtrtsnj+SCasL/S77rU7Iwx
ZAVkFWhBCbKzUismgmiyB4A2qJ+vSg5f4wIIKlWsGq7fDZJDbdxoyULYioXj5vuAwcQzayDa+Vnf
tsoLEOsJwFCVSzmPqaYKbEMTQW+uw3Gh19JTAycQ2mvpJ0o21kI/61pWqiwztkiVI3J55gVsYGRU
hFhaLWi0lVcR++FLXxi9GCBhdhNeQoU0ao9HZRC23eV+t9zQ1RQooyUA1ZjNrZtUgkkOAhH5VKgb
t1f3CD/geINxjA5WZhV/UZdU9HF18B7JApPOKgIm2a6Fsd1SajEI14oGilP3Cdtha9wav+QyQ+n9
GWnJyqoA7z6B/s1kIZDXpA2k6hVcFhSz6xrEWSFYePftqOC+Aoq7szrDiiP7migRutx7hz2oYaom
S+zQY+jN89EysthCqt4RCixcBLTIwfsmL/sPi+QYMRJxz2LRilGzwJaCuV2SKCph++G67Qcwpmvt
zSDA2H0faV+Q/fR90fPpL/5G1qmAn6+sM7ypqlg65nyyfV4Yj8LCd+hC2SXQ/kE4M2gJIUPxjhIu
6AX9LBmELsg/eZe+JvV75FK7JffE4ZBmfQE2fEXfYn5QwGNgpG+955dXeD6/b2qq2a1cHdbVgHGP
U2QkwNBRtdtZwLq/QywkVIuVE9U1kswWezISBFRJwxn1QBGT+/BZyLkrDB+O2e40t1VPNIyfm0sV
eQ8dwuRhapN9cA+IaLF40nurWF0evFS7MjfzYp+yVKCIeYnCstTCbPomnRWWg91h3ZmC3Q4vYodo
Cw2aXAXDGaJK7fYAK63hPO+vO/fTMS2nQtez8S14iti6gUHumeh/nGjhZWyCsIhL8xz8vJOyhaKE
9hpPHgZCkL7FKNc/p5COoIgQNMbS7PwaWPGLbwMTz2aL/FwJp9MvmxMz4m8G1s7ktgYp1WxQ1oO1
6Nd4Jg4F9QOBfRxbiKZfU+ctU31AZHc4QjJQKlxJis5yR8EJn+Xc9kAwt92Nwfqlh+d0qF31Skzz
B9UrbrZ+CddbY6VGM9mNPWbE9Nwx8T90SuUQlb2XZG6c6mMDGghtIbwEVuhqlqL/CihJvWiBACKw
mYuOYbyehvFPIFjE1q0LuLx+U5CUuyhumXGzM23zeHh5+BEu9fQgAJ6h8+M/BrFE/XV4z5jONzuR
bVP3LNpX1/Fl1y7s3btLoJgPTBVqmiwQg5phehcO+nAqw9BhQ7x9VmaoEj0AyoYLUpDDCvZAHxo0
8bYHHwk7WHxI5/wmslWE7NtAzMc0zPxnNoLrFe+q+GAF6MYs/8jUGM7cCwgDhwk3WyBn2K6M73is
hneADL/idadQwcolA+TCYx3Eje+st0oxGxMD45R3R5iAQJCeQ34dl3sMrIkg3nrffT4h6BPNr1DU
2hMdapbp68DJT0Gg3E3uc/Uypj3i1op8vSQYANKQbxmoUvfhkRUqtGB4HM7n0TViJ4T5Zm+LWhxm
bR1FVYbxlCIhBievKFVMTof+lIQImgqBYsAg2SadZ49jJVXs/AK79GEgNgBWHKTK8jLTvH1CyVD5
81X9OcKdCc4GhxTwZsOleygTT7eh4aOudtbmqN1JwHt8y/WgjPOmPlZveGqroK6x6A4c1I9PS7fn
6x8XmL71vH54FSgX6Gc1bYaJe6TjRjeO8iiY03cbd1EuWsSrpSxHV3W1aXxPRvcY7jUDjF9oMEpc
hw2Pc4z6X1crPe/d3MLZTBUPA/IkivFwvsKKOOd8HpHFkZAQdj1lLQCgXk6S1pX9YrpzJMjzEBH3
ACriC3+lS4wW57MXvSzq7jV+4jYy6oKrA+5S9pgp/XgG+uDwZljCRVJVcHzjIwkRN6EnQFfwpqkL
vVzIikBcgOpUkyx3WBne+L/4904alMK67Ft11kUGOvsp4e5y1sAXDijVcQvoD/Z0O7VmKRsjaQfg
RG+/0a7Lo3U7dGnsC/Z90c7/L6ZB1gD95w5a0LfvKQD3xhXyLS6bAo4I0tyWqUdbzETG6QwLpMTa
0SPe+Vn3IahyFZbP4Sk8SGLKo3SRx8HuvjDXY5VxCc/9p1HIfZeVY/Mt4/NOz2dXVXu1ytqAeLMs
aqCBB10pfFW2h81j4h8uD9vX1z/cS4bbYb6Y2cs5mZazULKsrjiNa5HlHuUY9b7tZK2SfNnxJdkt
kwdupPWEWlqCC5B5iZtz4nVEPWWmxfD8mSVBnUi54f/zyu249FUQdvg9J1aJjoiSzsZd8kT8M/tI
dPI0Q5310toniUSA2QIFk/jBfhyhFWvqeuJJSxSEUPPJpZL0FhQhNEfIPZaTDdKOW861e3rRvYl1
t2yWpoTngz2vNKO1SteJbO7o9esLLsKM/GzkbWCWjApfis7KsHOIoYJB916lPdCrlRob/CQkIlIt
ei0uE8SWrjMUpOx+O8CQwKpfcysHY7ofrOswn39SoVD83V9OB3HCVA+xk1H5/JCCPe1QYIOYgNL9
RczOcsxrZVM1fjmlX7NVC6E9RHHblEMbG78uyWbkUIGQraCE/+Cf9mNSguRiI7skxYPtp2Ha0GJV
dLZ4P96y/LEw24C+PbudXBbGXSe94eNWHhHvTOR64Dk8eMLUDT6kxIT91WVxku7kofNkTEp3oniY
mWjMFA/LoavNmE099WfSU6jZJLJKOHKZk90K00XFQJSZ+iiHZL4NcJu4isAajjqoKROZbuuddTex
uhBWUII6vn0Xi7fjGFBVi16oHomYTT4/c9PL+CHiFYrNWtM/XPY/aJphrLP3ldQ0cKwLmVcTtYVd
yHntc+/gJL+UbUjtM8cNXpvZHtWDRmrIZydqCl8vOuOrLXFJGDQ8BRk7vl9GxB70wPlzsFBqIb+V
TDUI4jYYzBm76bhMtkgJnKLn1DWS3gz1lZ9wXfyxFzka8sqIBPmJGz5ZI9yewDKMPBaj60qPyV3h
wqHZhs9jNGZY1MRMCPiJ+vyv1J+7S0lvlkUMirjD4SR2gLPlgs0U3DSbgeqO2eM4A5eP+Ve+AuDw
pt7qHxvOr3664vM+peMvGdxDA9nhxRINXYwmwieONsGrj8dmlvK+Cl9NPHaM+apE4wql4FK5J6L2
y0dBhs+jUj75BAVpjBfT3CRi3wSAtHk0aRhFe8TPktr4XkoRvcTQaGaw8JnqByXVKcXRg05ZXkBt
BhVA8d0NiDNqTtJGX/Yigj5BQuJUf8kpnsSJxOIhQgv2pgmkajtdGcNoUuhFLcIuMwwhBlN5j0d0
pWHVFzg6csG6seqdxzhCEhZFYym9XoAV/qtRwRWmUIVTDgmNKIbJRWw+E6vp8XIxxxuV3ziKzXZi
7Tj2mBUxrELZt38DKnLBGOTVT25w0gQgF1UNn2nzmeogREdgkziwWReoopJ7x+YQf96qkav27ZWY
ESNcqJkdAEaTSk5ood5HU1zxwtf66ZlISuQf/kofbvYuWru+DpWco9Mi1vlwe17fpv6P74FMrPA5
ZA9r9yTmU2V/BI/sP5uBTCyYm01KbzelaXgCJMVdlYiNSJQH0FlujWJ+3fpd5RWU0PCLho04F8ft
cfNNd+Njf+cnR+sPsu37usaZTxox5jb/FNwxBOQCzp3tXu4c3jRtzZayUfZw4WKvk1/Suy2O2CmK
lYemhVi/kEJbj47ysCdtlhi9ctu71GwVG2z5AnXiUuUThMoFI2UzZwrtCr84dIEqTxMzOHA+cLk1
kW0sYJUQp+OFqffQywtUsXxy1Q/nv1tUFMFAZM50dYj7Kq9XXT1DZCISP5zaTNyR486IFEbLfJ6t
3Yga3zpi5LRNnHr1t6qZ8WGpfdOTW2/fsa7N8LyF8DNpUuijldkdk1EF/QCt7J+ikExvDVZBa5tu
IV0GTLerSQD8BP5HFBJcOOSiItwMoIbqWGiadR17UngrwRGRom+hC1gEHl7kGu8xhA+5H6bhzWzC
O2ZbokxzVxvVH8qARvYZ2xGhlJpNwJ6VArW8ArpLjA3W+6ceppKhTb5m5A6zLBQSHmv0X+JcrVq4
HM227PklWvnX+top0MsRmbk/ac45MlOy10okqX2KWDic7I+EQRnpygxRSyc9ksUH/fhcO6gn0BUY
QxvFICyNmf9Xk5kYYpP5RhKoNK+QErCPmGhryF3Wil+Bpe5qW5Wq5774regbiEcgTrCYMLYdgIbG
ShFgYRb4tvCfW/N7Lp9gLh2O6edI/enbksmIbSfjAJMs0NpnmbRvSQeRnnrCX1szv/XrSD4nEP55
nEA9Ew1kbvXd3VWE/YWrjA6X9pJwJE8cWRpOPk9iDkBmk8Iw7gAwjDG/Rl7RRF0JBrBEpEIv9xFw
YHAVAi89DUKxD4pVMNS8kS52CkRDhMQ3+OIdQc5HQ9UXuwX/bWxTN7yOO3/N1P8RZKkjgZqJf+Vv
KrSpPF1aeGfRsckbsYvQRUgSqW8iNpGFO4KUG+3XusoQIPjwBCgc8N9va6cMNmpONAEVBwlRALBv
w2y6NYsF/5mIjfdzNNICCbWAL8BbyqSM2LyCG+lC3Bvb3pAT9PZWAKfaVWGWgj1AHiebnILPD+TG
5HIePJlO38aGK+4U5mIuBWx6axNZYuk5VkMSQEg0FChSn9+W4x/OMzAfhaL5+qmn8w8y5V5gk7V5
nESc/w2xpQLzCrn7JC57TJFUg7naKw7Al3rUEdYTqqZoqOv2R+yHkdU++PRqdrJNkW7x8EL1ydXc
ntY6KxbaYIHNSnuw6uq6FAK9ocaL/u9EGSvxstIf83xHvzUR0p7kUMo1njTczYI1DV+EsqtQmybz
0R67dn3FL2fJ4iqw1YyaTWfmu+g1hdJ1/i99sVY12ElCwTa9M+0c6Di7xYi6+O09AmJSV65XBWxM
MsjAzORBdCAOUknlO4tQg0VE6iRaZlLvA1Y1T1JEXAstmU2odPHIuIXTvz2wyrV37mnFAyGny3p6
kZOl9vfFpC2WzrnIYzJaJc+WTae9rBMxz1G5KJyMs4oAy0p6JP3Fp9b9Z2WZ7L1KKX78emHToqhr
wk2sJRCwbwshC79J7XpwozTi/mFePJV7jkDI74NRkszcJFlps4wnCVn9XnVvR5zVzH2G6yIqtfLL
+Q0Dv6NJ/590lPr5SaV8KgxZ3HDKj5U8TUvy5WHsmswlL5rTlH3SBirFr8PMH6UIc+o5vMfIXRfb
vuVIxXYQoACx9e2cCNyPXL6vDWnVQKyxyZsiX6rF3o8+urqZjziiXunwvNFtZIgOdOc0F7dpXWWD
GOSngS5t2XsSZolPY+ozaok4bA3ik6jF/Cht1yhU6n1hWfqddqGYCArD1bMLlIHBG2Fs65cBofhA
dc0LwzbAG65iuSnXercb9mJ3pgqYXbsuxUAExQesk2jIUOp7W60mkBU3Y1RwkzhFx/GmNtxiBS91
GRhtsWOHailFeMWsd5uisCG6D35s+I3xQ9d9mblSzbPtADzMrH00GYQmnzLy7/Rjy02HAfvCgLeu
jRA+w4Cc49KmryOre8iEidOL4fESSvzQA3ogDJfkvf1Ph8pGdAnLcFFzZAhHHrzNqX4PBLNzb7xO
NWia5YDnFvvkqOob6iIr+Nrh9aAWhdS6t7/NJC5hwsvrlc+GIDuBCRutrBmANsJZHFjtOa0+b2vb
vyeq0JGMUVs3KgnDuNYSpuRCbFFRJWGfvt5IIwyF4LO0NPUiPHQ/O6Hixc1MTct6eZhPE3Fbv61T
JmFx24m42IZzRAPXuY3D4YVG7zgUJ12orq/4uJh7d/0UL98JCNthd+ZeaDEqLYEfsFGfKRnBrkJI
eyWI2aaOR8j8dsvo2UJYMii3EmvFGQwKONdaPG1HmRcKXs2qGwQpzom8xP34Z+2LhdBE3JfU+D+o
YVVwPfjK8rbetwEvb+kw6V3zZexHW6LAXfNVEmRuYmUgouulZ2qD/t662tzTwXcge24CljCJC/wf
Htk6xHIKWnMHNWLwyCtUheFe9CigjN1bCAcu64grpfheNcdRRLuk4ml1aXHE9UDH+7DZ5ngd7IGt
SF2JpRIkPXHQnIU1KOK3lr9IvTh1wkpr5n2DkU8lJUnt5sF9Q9SVVFoUWfqwG+/MydOafZD7oExY
18qh+2CvD7qeOKqSJI1P7IBsfN8OvfqBtoVP8lb/lWun2XH8/C05j6XOOvaCcYYO9JGnnlX0HaDz
FrOoCcTUdfAgZDs3I9BG77C494UxBzaM2klAtbmgc2P64Zr+yu2rjsR0pBPl5i1mojragzIC88VI
XeIIwK4Zd82xRBBChSiVTaq4arsPNi1cosrxkPqF8UD/S4Qy84OIIL7WZeDxj9jjN58eervLrlxQ
MpLNCtfe8Ji8Gw5O15jc+hraurdpjO1GiqECat0Wzk8m/JSzkCXBxCbnYoN4DKaWpAzFd7WcewTP
z7Oh1bYxbK376ocuzdOMv8hHaphZBlObND8jiwSew1RXEPfe9VyaJiFgyRY5asvLiO513g4N1upX
jfL2Oxw+Al0ZQHgGNGhfkN3NsPwjQ6z+agpmO5KFE2k8cdQfNiqsXhlzsY9Cn8YH5hrjiAW3yX+F
g+tNxHVeiH056B7qKZ4D/LlvRQgCIBYWvp2+a+JoUIu/dU9Sq+pV3MFUcLsErwLSYqhJfwZqMdIW
/r9folzrhJqHSZATO6OtJuUHXH8aW+RCgOFtMk6s0h/a3upKp6rSsBqHBpZiIukSajHq4aAMbWDo
ZhR571uVROeNwXaFyYcWKc/uToUp5FRFWq1qrfNNkUt241QGr99BWa9UPsIInd8Sa421gtE7pcZN
H58jsNOtnJKyOanl8IKRCJl97OSe69+YWxGaSMPSf+m2lx3+lQfpsKy+D22lYA7ReJZW+oVHlCg+
xzDJ50WBuD8V1OkSX1d6zeRsprPeZH5OWKu9F+wt9XQeL0QoWYNx90C2hLqJ1VV+u6Vh+TH/18me
sSg0BjvqHuvn7yKsAIE+7BS9odKjH7bafO//ThPVFA+4/pxvFfrbHsoLp4n4ydHWEGO8ih1Dici6
N2M4KTKdxUpoSuWYq3qCJFrz9qWvshOu4KnCB3OfV0z7s+l5o+O+w6Ajv4Oj/O0DfmBFx+SZvMuK
OdWuMlRyHSp74G4dHm4rsabuED5i/8vU0xXY6Dhsy/sFdVinsWtPZcCkWCD84fdDEN60Jq860aDU
N0q7qgPXDxq7zuPqHYBW7GwhkIuzaWy+vmfqiO7FI5SKoN6FM6bvaUC1anEi9ZgwRcFYgYNGMF40
niro0/JDOWB/tivWWDzTNNpx0TUvFbxZxaJOGg1zxfTRBT7774HEXa4onWyHrmkfI+CBifKUboAy
8c47Ia+vcW+NHhaC/O+krMJEjpb+KyHQBfCQ7/4h5IQg3M7/YaIOoKpBgOmDDYqj32wLTlsAuEbh
7d4l3cbJf0MqH4s0gVXIHVrHMDfHMophhQr71+l22DqNshjifqlvgyPrMSH4PmQaemF/Xa8t4ycF
AUhyzCGPTjafSevLCm/O5jcFd9vL0/1QLhWIB371I3vy6KNQUBfxrygw1swOi23//4VuLIgcqFeX
q+RZtN5poR0xvF9R93cTaqFuIpzssjVsrR2Ik4RpOKU6ojgN9URoDFzmRtCJVY00HudZHYVgunjJ
A72aLdUR7dXyx+5uyp9BzQ92HgiwfhOvMlPaIcTZW5PwTT8KNkvXQJs6/Je8fbpg/9mqtB0qxsJm
6KzdPA7tAY+yxA7/6NbJdnBekvX6aq7j62xkPn8Cjuj2D5evrgU9BSlP6DtH2hCwH/DKS/RQ3jje
IbtiH1AiDZJ2wZcmTpp1cvUgpgbeRWZJD4iMQMN09YChe9PL8fLF9ZGu+ebFlxK+8Ezs95aagnR8
ZNgwFE7LL+YdPyuMUadK9jh3kmjdgmmLF/Nhnbrh/0BU2qCJcwmBfRz+T0A+sI+WNkWQ4cTnBrAG
JERasoUGPeNA6JfA2kgHyz4RtIHFtYxsxzc8EqWxYrnIwzBPtT1XBfGWyrZgNuH2zhJjiuNX8J+s
zAsdXa9HynrZHbFXB7nHy6no50Dz51PYZk1ZFJ/a+/48PXYqwRDr2xB0b9zQ3oYxUNy5NW/dyKwe
faSQiY0gQBDuDnmfm6VvwGbR8TwEE8bBa2Y3CSoaIH9BhaDhu+d/GMJN9n5oDEIzCfctb1It6+5M
GJnix1sLRtX2f0+Hhbi3O9rsNcw4zJcaB/P+MTuYl+oPBOulTb8zrSdjxZdxD5r3DkVdz2pU/UXb
wwSMbdfDp/IAm5drbULyz0FdB2EmL8+t0Dw8Ffy4S4Vx3ROARqmw9Sp2RdnhhpH2ODixJAG4FA9m
ifoTFyKhek7nltSxdNJh2XPQkfbkeWnkX4eTuFVF4emjKPLOP0BfKK6M6SojVxZ54hRman9Mnz24
g6iDgpytYGeMkOVWDBs37NaVXF9N0xObNQ1rR0CAaH5D/O80n3NDQaP3yRqQvrimRyZojq54OBxR
lDhKKqDnDY6KXqiTbULT+OVrPXcFDanz6YZ8Y6P2MhSyZyESCZPSn+YyKYToYLGFAlWcXrpOCKmc
SEt2GZhu20O9/Ntch16/mM8GVJFmyp1ELtmN66Lt7f24feWa9q0/HGxRGLZ6czXrCm8Hh6NOP9qA
7GouInjHOcVH9e0i+5Nm+j6zAwXF1JLNfED27VyFeMSlAz3U4q0+F00ud4I+BfQpAMaPcD7Ja1vy
MKd83SGj0I6ns59Q8HX6Ko6HoEUhpQWgJ7jxSDJ98abRUJSm6yNDayH+rbQqJ+njaTa1Nz/fsFYR
IADTXRbNCynGcvOWka7LZQZIlzCOm62swNx0ZVJzosDjUclhjAa71kNT7dXrn4O6DTNGOFBtc/Y4
rbQd4UB4g61eYxVW0OxbdGlurdUW1t3vkzhnylptgajwyjsSkpx5WYjUID2RIUUkLZ31ya4yEO3/
LVyb+1W1A7yLjG/K1gvA12eQzkigN8TUf2y0Q0GM2Bj/BFjtszyOINVRcia+Bj8Kd5GYZ+inMd/Z
Fc+34yK9Ai5xFEKv/PNqDeAeyubGfNDji/XC7xGD7+DvKHDf2FbeCWQbinisxMSmzxGe9brrxGXC
d+apqNxric56ZQt9p8CqAubpoxyQVLe7H1QDCrZMBhTZvcm15VBs8cMkNW/qwNSdvqf26IedAQN4
4iPIY/OCo7BKSzC23WKOR9vzEDjDwIdtzoKd171/dITimJqkFNMLRzw64nvZxVEW6eN8cNq+zsEX
CKAzqBOZtDAJzcfEYb0Bbu9JvsGIhkLsOFVfrNsPg+0TC577xkMFOD2oVJqkwLjJM6FMFswnibBM
9RKHhDuAYnl30D4eu0JUTeFYgkJPiFeI1VouatEPMtt5l77MZElyRZSX3zEFfNcK3jeRA4oWJDSv
pMgNU+icvUXcKoyTKQZDeWq4VzaBQouLdUk+iqkPzcctSU/7+uvWf6FQZDMvn2JHrn5cvW9vy8jb
Hp/zTH1au8NHDEfS/DvV7qOcymfEOwjcd/oyMoUfJaXl2qsvrnP88lNs1QkVJa/yrr1wlyDow/O0
cjtWN5AVuWg+CEn1ELi/zNCIkpcmytsOD8Hqj8Cs5UMqAUqwFJx03P59/XjGdyvlUwVlMGZhgD80
gdQLVEG2MdyDvNjKXGVDvfIKNSsn7KOHjt1FsapAxVq/lj5R5c3qY+ARg5VfRHvGqkr8Ja0mf9Da
xZ9S/1PetfjUho7EXX26rYseIniBRmfMd3818OrXUsHdt3jKatc5eUg/gqmGjUW2S7QciT5UH2I6
GEQsg/kF15qbrqsMcAcPwnfKxSnjUHdWXYAXlMmXBPoj75r7geWgGA9evY0zlhWRVOfrwC4X9XON
kg3wGLUvjy/PTZV6t4QXKRw3V+nxXLIhDrRLWN7bQk4tMzLna21jwPuOrcMokEMyP/HtxKLwsw8H
Ss+FZAtyTrxjoSYsWDxktnBkxZrJ1k/+M+aZOp+XXzN9mvR8uS9mdUSU6Lg//nJD6XrFi3i0FUwO
mQJ8j5d2qTH1r9JpQXEEPo3BfWxUAb6IDMOLw+xLrlapGl6id4ZDR4o/BmSfjkdcksuba2ZWHK5p
MqKXVXsPGqedyiikyzu8sDkzsTRJCSJaGUnxCEMpoa2eU92PTpXKJPvPEgbNerBIjUf87FxncQ9J
GYaG2koN2uoyykEHwq8lD1QYZQfH8vyCaYOjHJ9+Vp1diCNgr0UN/cOHyZVPTgfZEhmGCD4OEGcE
0AW22jdhdnS+pITMbkMkUDnDtXdvF88ZH5JPJBKo4imw1bTgE0k6hgbtXNernrsMIhrBaloI4+cH
ctP10f2lrYX7sPOtoGF4JpXyNS6bzj9CrYRNpPFL155TDzqaBogAed03IVLf+mD73WM7yokwwCSI
MUurFwYcSh91p9xC3HuQ6Gnu22o0ZHGjA/W80kHL+xFFJrc66JlrVgFWTDM5kKhFFkn+uFxsSe0B
44sBpMhTgT8daZmSifvhlruRMkmUn6ht+jHT8qYBZbpdHkxo2kUZM8DO05qCWWUZkVxOXeu3HKyi
wDKgcAlnwWi+vICeHvUwZRAfgZmRkSmqJ49svi3xduN/AirV/9lQw3VUtdFBOb0ri489BvE5tgPm
3gLweeB2Mf/QzzT0KHDP4j5uj0lUIypm/yGetdWHuJCsNV7ZXCE6BpuiIkkAWnGSNl8yKB29xSP4
p5QmAvgExnX6lVpjjK7sAj2oGg8YIy/cnqHcFciX3YZvW1b2R5akdDRhaDuC5RxTfeG2Ynudl9aJ
GmBM1qPFZWEMqa6PFeQl/RF+JyrhFvOkKRGlY2BfkCt0hh2nZRN1fvxsUbMKcvILFB1ih0jUemiu
smsuoO3U6GUeJfYWnXHqLznOR8RTo5tjShrxBxE7rfAfbTK8Y1shShlh9GmPQXUwIn7DA1hGmEnR
RyU9Klhij1inNNw3YJYDtjuklwvxHFytU3sFBj1nLrQqdoW4jsDGT1PTVN73dPEXhV7KjzU9H9jC
OmMjMWJcEBS//TutM8XYmwvl+Y7hV5bm48mWIZYbLkP0fYTPV+DV+H/Lvh0Eg4jDBMUdZkFjg9bY
H2yNNY9llLtrufCUrFZg+ueMFoAISeAp8rR8tq46vF5nOyRZHmWsxqMJqMERFgB/OGv6M2IdrNXn
q7gWnko765D2K+bRMynWNrqn+mqepOzuG9HoQzXcg2M2Ty8Pl+4tD7istl1ceS7A3U07rkOLcYL/
FO7A8vFXMrofYKpBntwSJPivKljX8vs0Xj7lsLLTMpW7e8rjrsYPk8aNSeQ9BPUrXqW+ftv6jSv5
iIe3833V0loLVJXHJjkVLmi5cHsjfSLM44ND/3/nXORpPbU4QMHs1Vyfq72dYsphd/IsWEpM6EIm
TYKFOc174lUN7h5szKOqaNTgrcKmlxtBkbyPN10aYjlK3zZaYBWZun5Alu/0Tx+Bvby5G+kfeHxb
mw1ihHJ6bvArmKY+oRPVuWf9qZig+cl7inReZqXBDooVRXiRPmAsOYzP4qlVr6PqgjrbwXCCrJ/B
w0J6xrx8mL/SP/Cz9LpDoUBhs5kqfcqCqUOvRe4/9r4Pm7Fs6Ea+ZktGTt78l0m3hsUoqklcNClp
sAwfm5fwXRZXThbkKa8sqftzT8Xf5DflFu+E1Tq9jaxFqEAUtlOwSQsIuOP3JA/q9e7iVldSsnp9
tuF8GtbZwjlBEBRoj/LtZ7PluW0NZb0jGsYuUyKxU58rGcKHUhV5JsJxBfiz3ZmybUR0PmAOI7nc
MMxSi3EY2PvQnoWnDpi2pdb49k2lVvRTGffSUhHnfwrYRLC9hu+R77HSrjrOPFGcSngAhfguSaro
zwdrYVPxbSp0dg3zy3sfAgO/ySCCdemtWz9JAIg7ecpLM5wyLkfsRA8prtl6olqbyZc97G6FpRHz
em6bwsrvRjiASiDFUyze7COPO1LoN75SmjGzLeoLmEzVWXprGp1tyoRRTOlH8mYKWJZfVDkr97We
cnQCXsBvjOecKLhfcMnOL+qofWq47qaoC+Osa15CqZguAXj9FJbNal8JvLz49S0Z9Nkm/31oSp5H
0qsSLIVx+e2zGAr9Ndus+Rl/iUVONX3VfeKaOk7+rRpJi/oyLXB3iifrRmSRtj1Su7yhOhiOTUBB
fWqNjqkXVPVZIezYL4DaAoNsieFaCyS6Tji8NEQYS6OOOBSM/1LozxEsrOB04fMcjP3gMoCWuj5r
dKfl6UKqjIKYLlYPerclOboXbgKnyz+ohXDgGxCYzjnTZ3sAGPDnOKOsLofag7ZV6DIRQbsHfI8U
ibtn/efSYhjSDm70XJkBzxarCSuPPf27377QxXD0KywDasfAhqaavUdlPqojPOkL0xRqkAGFoBpq
8BhhF7VCaBW0NoVkBGtRsCfZVAUXlviu5xUZb/8MWuu2cjGQdrNug/mRjWyU7YHOYR4kaecG8Soq
mSOIblRpCCu/8i/RVBfcHH/KvlClg4pP8NThqzlykJNvT7KGkwRHr0ai7kRtUjx0X5F97AQNoQHr
WnjLdHMg4bIOPRJ6JDKj2W482w8uoo/THVEGVA/hJRqWFkPkeZ3NHLYjLZrieRfi6EX+X7CZLPhM
OKKYSj6pg3ci+c/1C/nRqg8E3356MV0Wk2EYghBkPWenVXdC0eXdQxQa0SRAuS1mdCB9UqPZpgXH
YN80zFHTd9MhQmopkFESOTsIgDbQ7/V1Hnhz7Z0NuAagTshwmludLxIILefo+UYFLINoSkbMEhBc
M5J/7pVbjeeNt/Xkmw0vBpYMKSFsilyAZ1INdIrGTNDp+TWqfZ5Vc+I/Ry+CQ8ta/vuYjCGdLpIb
VIVcQ5vg461v/UHNW9kLcCHlfaPeBlfUu1VGSBDrOmlxeJTLRuWiqSYYpjIe6HmIMj19CoSLbH1R
9cb7aNmBQfDHSHgMLsvQR0sBleHECgbdoO+7M49sKA97ijiYMzDWx/ruBFV0fvaBfTV0SKtvmlDB
Bi8vewb2tnxZGwNRrq6Ikyd/18OG/H2UJsEYrnOuETxHo7rqJhnN60mYwgJVPCsCqO/kkvp7JiKr
zq29j0hTjdMsKRMXNhH3qKYZ+ytiiceLPbib6YWDT8Qvbt4ghxucTaPBb2suA+T81eH4AApzZbko
4aJxipw174ETelhwVUZhfV5Ce+ErdOprPSZrzlt/Gn6qwC3nqNmPZfZORhVTgv/bAaAwYbctyRwQ
J5w3IwZdYODVs9sR/BOxt/kWBll+KXTJLf3AVUXlxohwokaPCtTfPcqHdOIKI/0Q4QWdg1PmMysb
STUkdd2rjt3/819RKBXJb6maq+kBKj9TZ4sRrEN06PUF0Q+IcVKvRJpTwvqayZxEeOVRhpRQWfKl
aKzUMObdTOjS/5YV314JdFxfnOVGuaMzHQSiFo0UG/tnbfKia79uzTmdkxvztyxYu7tm5karADl2
cEPqV/Cww0aIWZp93oXdNMf7PfzQgr/BnhBItrJyHCt1oaUD2zxPESRitCX5rhXjpZJS4UTO5Yiw
HlV2l0O1CNlFy7npIIyxneV3ZEu2Zl4yhrPizS2+Kn9ylg1dbYaqGuqNG3DR3NodMVmz1E/lqCRG
6ZPYkgWHWy8FTnKvymHi4hbOujDLFyF+l31FiXbQjtxhafcL6oOh+XvZXrVrNOhTyOunjcq6UnfC
rJT4fex1tFHdBVuX8YI2Ox21QPKMtHAR3AO+25gc7YV94fAGSahPFUkqRKTGn34p5UQNmDqnlkC0
BVVfub8tl1AepA113ROOmstCEzCAlsDehSIZsgH3G8wgGd3fUFnsarIpkfsS3LpygqruWlm37HpF
o4PaVf1jGd+UVGGjHp/E4daNXL2ZRvTgAEY8zkhzb7FUUQCKP5dJKHTOy+S5ehNjDJfBNzuSdtq0
3KnWlRXatkCutj/AvQM6iShKHjj1fyUVgiPUHHMglnACIlTrATOIKzjirjwDef+/l1lzwgLWYNoe
K5uqR1Z8ewwktxAfPq37qf0fbY6oUyq2nayfpsyfpI2t3DuFwYUl+63WY6eh7326Rp+Mp96NK3C/
/3luzV8wetHD0qQzSStAWVYQxl9G9Ta678VMudc5Nkfih54PB6iTR0IkvDxF/00sPh+55y1g6NcZ
CjgulT8WT76TLiLadwVzbOxiDDXyNIJsXfVlMcub4yPGWXB4cJKAd0scxfY4MhHekX9LVgF/tBLc
vsoUd/xA8zd3uAT3VubyZFrCNT8bRryu4/fD7EC/ndFUGyaEnNqXSUMhKixFvtHEm/lUkA+9ATO5
rCn54WM5FL/tc8XqWzOCwNIM6w16yeU0W+YoLNPKHdvnKwH+r9emdyIrIln5J6h7XLXsm3vtxKCq
sEy9K366EU+MPGt80LDHZAlSX8RuRgydqu4x/QiswnCgdKV8EPk9FFGA1GcPWGiaqSocX1D/sqAZ
Hka3KqVWDOovuaQ4OH4fd4RZBS9nGLnT2F4L2z1euDkN83nDUzH4r0ucwHf0pFVf8MV3XMzRV4N4
EF6Cr408VleIReXzRAPJCmTK/bIra9SCfalyUizs1TvtL4+vhmJpIbI/d7bHoktubqc5Ct6zUN7h
jbG/uaYuq98f8+OBUJQKL7e0wi1+PV42zxoxJNtp2bExVsU5id4Lib6npFvYQKI19TQAJm/BJsdt
nRi4O72Yfj5Z4BDhYfz+RxxVVGnahzOxKB6MfvF2cu1Kx+f/iVnlTPV9E9IK9l0VHZw7WICiZ/6U
rVvJiwjrqf4ci9ffR23iUIaTDSHCafhrfraoxRdwwjrd0hthAcOGbvd2S0PxyrM9U2SQFqN0Et9+
7TiTefJM3dsMIxxzRZXKpwKcQpRfosTK5f6I61aJ/F14pC9OIPpzhF2h+iRD46YDDqpeoON6Rfd+
l/isoBNNH6lzP+t4E3T3r47hbqLDBpqSCzEvMsEIoy0YwjJXn5OJSHW3tXImvJYdQGE1hJy98kvm
/1ayyH8fr4iUqF6BmpVrhsOwcRF9EG6QuXOZGJOHjSYHZ8llkVQocr5/JJgOKAb5flf7BgYsBKBV
qILAJvoknPBGBpyveT9EiWr8q6n+hqBreiY2WfaY4Cy6kaalQd4pLXBMqJSfw2UVK5FJn1VlnMjF
uQfbX+MZQTr1eX/hvSpbZvvcRtBCj9+5szMEovnlCLGVgv7jJJa0m3ilZpyxtJWk4jUexIRwoyep
CHl9E92H1ttUXgkqe1+LsYOnTFd6sC1FYkpzL0JExIsOqJbIF+ioLmltKdXjUdk0sJNhnjH9oN97
awb5KmppUvEdBOoksSv6a+zv2guAO/nfJr67PCxvX/J+a5IwKEer8l3Mio+AuWoyAhisX10PQk+m
EutwYBONwc3Oyh+/1H7NXqSD7Ldm7T21cUCnFvdJhgcHYme6lXP7gAfImyGkt85nSBdS3bcG/i92
Nyasc19ZSHB8RMwMvYfplhpBwz0czOWax1jau7NYenoEQ3dejsQMpzz90mLDeLpVF/hprfWJ4NLK
dIP67k6zCzzB+7sn46Exm2p2Uda7LS+qZPsZ3Sob+QK16n76vP9EmTXcNUwJyFG43WnOl2kE3joP
wWv3l0s8qmcGLhdRkWv3xm6MRtn3RlFsS/4K1Hyu1pGZYHnwaMvbTj6lmsjotZx6g82yeJqfJn1W
+gQ7TcooU3sFKFHZXdLdwBtl58Y5V7q3IvJGlejANiMfpJkZ7+WYzRY29dGvZaRoD6yWt+2i4IbI
DsBef7gVbJGmE2oX2hXiX/o9AIleb9qPkPh77//4LENxod4ZhMkOTgMeCY7n376OAzQlgIFZMXEa
719fKCMaOVjxpZ1tIE90EvRR9VpCg3M7rGLk27pz4k3GYmbsd425A0VTsOCQP7qOSfqxZ7BU0vyg
7IWIFA4uKB5GYtfJUEaa50spcWobsjc6MsvbFjQPUxla4NTyyDm93vnn2wZ9c54mz+Fu9Js+Ctwz
ZuVl20jG8J4jNklUEnW1FYiWH3eucQsDudz9G2L439m14xij4SQ0/NowmDcLMmoBUM/wHbVzX1PF
UjPc2qAjgWmiZOe4HLqTSJyydqvR68vzagNZKDu1Cmfkn5S1hXJS2Q3WiuP7U7BrBU5ZX4pO7rm+
WoTwhBVnLlX4H3Y6R5dKTNrMQm3PnPVI/hxMm6MxBZYW+wkb3L4XuIn82SIt+jB37ibSNvtYrHdr
NSAZUaohtlJT0qieSaUHugmUndjL3QYkg/D+6UNy/KGl1eL04gRJhtRnUPhqDoVB8TshxV3x/tLq
Og9AoAVBFhKXysBmk2h54WPLMFvm6xx1Pg2VHE3bavdwVE7tTthHqvwjjgfpqKHeopZGQjZNqn2c
Udinh0tKC+Fw/Ul12p4CVNf3OJp4CD2JzM50NaqvDU9PRPAl4jcJte1UmK1yJVBO4JfbBlpNSSyv
2MVKxm0MXmn2fLak+smT+NS4hJqwpbnx0xQ7EmXotLC5VNhywR3gChD7vU/X2rTUbvqa746Hoj8X
nrionCIRtT66JL3Pfw+Dlueb9XNmvNL+VFjw2acXbxsvWijxhsq8LKlosQXdnW8mMJBtytC79DF7
/S4ZA7EOqnNuqkRqr83CvM6ck9zQpkymE2EYfIyX6aq34BTCt626Q6Aoqh8nid3W+X+yKpAv48mi
VmmBugtX6LuesX8XWQAEvJaqPE2EDr5tkhNPFAmEqr6x9d38b2ZkP/d82KXYAJfFTSp/gwcs8tVL
zUFzkbq4ULCGKnS9/OjOlXLFf9eI4b+MbzYE2eLtW6e/U+9CUjHl/gPSve+uPQbr2miG6e/oibNz
/GGNNB13QEsRCfKdLXkWFWUrycEyjVt8pnvpu2uwDtZh7womk2S98ujqo6Cvi6p72AxoiZ0lv/d0
RFxtzaZ0OlOw5stL57Y4qnHd+lmXtii7ribMmFt+XaZN58Elv2cFF6+n1bAIg2T/3HnUVcY+q6jg
GBRjYSpqVnfnutl9QJvdsmyABYEcXwtrCeWfY6u66BJyEWryEp6LVJ6ykU31yji7y5kWuaTklHVE
xf4DgFhB/F+O/QdANrv2ntSpgOhc0ZB9jlJfBGQQxAzsd7Zb6cM2X6Mhaq8TFjcRtHVKVyoRvmj0
wX5uUgJeTndqnAUcIe9oCfCGwUc3IakCNqnL7UhApTBCOUF/gPpw4vk7uUVScrvACIgnWUHddHYb
tJLpdkMAGasURBg5M4Z2Qrzd1tE9ZPbo0lT/ntxXR1npTH36ePwNRa0TiMOR5SQnyBrR6UXxedIS
I8+MX/AI3vw5bR08y+02cmdK63Y59eOa585eHhXqinvdcXn7wE3SjA4Qh36uscaw8Q+QXK+ktPn4
b+D/hFczF+bt9mwyJSLvxIUfDL8eJY11JpR7/WLUTfJpj3KWagGco+0PnxQNv6+3fa03N7GXBAqH
duRlYUkezAcPgrmNaOBLjQR/5p24m5DIfA/u4cii/S76gSOY2rUHck1NkX9ERjKW6xofLPStxMeB
TPYoKyGOy9WSCG0DRGxUI6SAnXnDmerHJywuNDgp2hk0MVgpqV8zjtSZ+/tFSBbDV4P288GGwHUX
JL/epyW60B0+tnoPmj3jqiK6qJcV+T0K5G+Hu6t8Zkl6GJXxE5MdwQeiDdEERdJ5ZPhX4+8TTPuI
k6sdntf1VWHgro4I9z3axbSAiPZHJf+vZ88UsLycmXHPVrmniEYYOJNAt19kBSj5qMgJ3d03yu4c
iITzfkiPUMSNuahKEI3RhHQivZEyGh5UALKrpzLdAHFjiYO6Ra6TiA1BaJCYqE3Uhw0gDavimG1s
auikaujwd/HMPTfbud8LFOdNoE6MMOeD8L2OfCPt9GSy7WrUGoIplI7445EIPucI0OBFC2HXBgY9
BMfppMn6rd2WKo8ydiJQKxZAeFHdisUawzPsYjnwdUCuxeDBDzfi6PwP8/gwwEbov2Was5flEi/h
2TMfapBAn23QWbo5a6XyUes7dfSLogFeR3jcuIilT0NCDKZvg9AhsBUaFN+kAE+zjiS5xWhdiI4B
oeiyHpCXfqBvvGww/2PJMvcdqZP5AicJmbbLr/VdTuG0kwQeZOfVmimgmz3elFv8/1ChbyUkqEWI
3AZL2vKzfkxSr39jx8F2ROrz2WZ5ZPCAEOhhCudrI1jgN6DsUd5xtpRBXiSMBKNNqbaANbdmXCPO
iOGHOs6UF1e6QdFt03prkatwKw73UqQm5vMrX1Xv4l1fVMawvck/2kf2cNGGyEGheoTb00Z4cvo+
ojgalWHapsFIvfmv1tU6jyXuf/e5S2ytXgoB2I44qo+q6fRAFF3W4buypxf8wshXPGXExvDJ7eRC
CecLuMx0Ibvw15+w8nyvpo6PCKjtcfZ/H4E9qQVzugjQdvSBgfjxx2Wg1uNckPAjzOp4f5Qzo5Vm
ZQO/ijU0jC6nCXBMtecZxjv6bR66h3ivUA+CZ3q3zieE7qjfrWjyIduCtDPEgFwmv6//PaJdNJJY
tkT98f5PNGkVOtNOerTomFHGPHusTZty9CD8jOlCeUWR6zyaeSQm02TH5tcFZbTanyF8d0LfIviA
gQty2ZMQDNxCXSAS8DnuqUNgxcqnChWuVFW9nq7LyFLJ8fJLwHkuWcQoje0jQl9HODrjPuV0pBMN
4nPQZky2udCwdcb8NYmIadqANZSkMAiLMFMmIYKc4F3dh/YFA/cmE/snOgfU2BoEBz5491XQn6AT
OUApJwjihIWHajTrPVTmw0S/0acB8cDtakxNjNvXDzRVB9tjElaEj33X4ZfSKLQjTHTtXxPXP3mq
JN6oYcTA+xUfIzM4cRW9t3ZU8QTxwFDeCdTTENqp0OMMWObb/RmNlk2NRHfKnb7XJQqyDH7GSYTd
FYP/++RwVlYGxEoawmJNklbD+MCO54EhgR1FLTunCx+6tfnz4JT4XeSLy7EhKYtyUGULU1xcBIas
5yMBrtJwqiGB0FLZlfj92Dlh1vqensLB1g+pmFjJozyYPt8ZAIfDpiNwlIpPVXZGsF2/YPPv0n+M
OxWpScBTmYTr0tY3XoyPHhKNkKWuvvX8Gqt0YWuHBLcx19i+e4nwN7PCD0LpiXWZqK+PekAXz8iE
75qY/o/ZQWZMwOUXe29TzObEE+VOnMMXQXcTSI0IFWZJ67/Ml15WQjtazS0WeX6Nw6FlsCQdJyfy
bOJW7rsv0vMW1nZ0w0W/UojHo7+K4iGqo9fjShROJZq/giL/T4QpQbAE9cBBxvP+3HjkFx5jiMQP
vc57PUNCKSGZWEtMY5QgHR9pP6LmiT37bIG/4ao9LeVIEWguY4pNyF0sTZ08zJ4JMWxnOds8O0Ki
2XKMd52wkcxfUjGsTysNfomhgruj3H3Ure12R0puAgLYG44HdGuVXbjfXOxx9+jg5HsqrpD8NXpG
iDWh0njNQK/rxtcSUoVzCGA0PGLE/kv59ATaJQvNECaRCcjPFRVYtlbe1IbOc3qZSsR/kRjdE1fw
pY2VExocAdX3nhv+ObpEsf/USg5HZjyrV5RfetQoAUeDEh9XwExnJ6Cpmsz/gkLigGrhCxFWga5R
+uawa1CPRb8+/jj6MrKC1IQme46JzZfSELtMO5mQ7CnnvwB8Lufx5kBcCw4CzrYipARjr4mWoK3M
5u5HxSzeUW3jUX4vJiVsMzcrEeaUVTUAVtFv4Mnn/oPKAyqgK8BVnT9lqUQeI+emcPdkDbI9JARJ
MBZoN0rg7vpuyrXWQzK8KH2sfnFEIxO71OU54vQAZjjnuCpHD4JrhyYYynao4v0FVghgyGlw0dPS
9PALea5xj0ZumzThOQC8B5lx1mmPdB3JoiGEJLIYttc1tknG3N4hspSuDa1aE7ork83Smbzdf+O7
gAuN6lYI7zeyguyW5Ync9/w864lCEP/Am/AFhWpY3s3yDUwyyCk4mNd5v5ejipA0SI6m283H6Bls
ycJM03OxKQpJp/Vpvi/Kgx80kwxPfMRdxp+G79eJ36K8gocuQoAtdKsGKFXXK42tM6u5S/q+EL4D
sX0ALDDqkPxuTl/+B5SAeKa19aYkPr95fuv1TFIV8NuTMDOuxDuqf9THgQmkXiTl5TkPATlrMK/C
kGSWwc9FuFm9I//xE5uYrmjF8poUZA+QQyoqiY/fcCTnGZtAIqCwvNJRHeIgVEsCawDSz6pJQ7qZ
5o+wBki9Dpl3jtnVtRlYuUoS4HO4LU0na6bsFhgV9Xy0WSVs5FZ7oKOollIzeWsyJWHQhChO+yO3
JoDKf5WHDliSjEZEwS+22dloYYweR+RRTAjMZS8sP064yaZPqfJ9UMqI4r7YPFzm1raZmLBIRY/q
W09zu5eFLTPXe19DfTnh2g8iFjT4gNQlHV9tBadeL8sOiFjcRi17MG3cZCxDdYvnUmKUHXa5O2Ga
RdnSerdkr91w7e+4ukIZl+/IEjlC9Zo502TwCFglnG1ZCLA5746H0S6CLq+K2yWXV14BAkdzRbr4
qQUBHijFUlDNmw7lMFmO3u7ZSZpCFzTrLm3LHYRhByVjCuZ0JvzTiF9jjdOWgrDuq2pfvRxnOlC3
oCv6NHAUYwib3jedTBQB7jjIaiKvh5cyA5O7ykl4bs7j+wKzrMAQpGWf2BKRoUQhAgoAyQjhoTXD
4VTP92liawJUAEHbHsr+bs9jYah97g+pzlfTmjuYTUuIulYEsbVsRfEbqQYF8QVVkMW9qVZ3sflw
dBM+5JpoyDAd5+MEzBo+ISK33Fy0GZdstllDfSB69lUHzyQc1l+At55AUdKZ9+VRTqyx1zeRWuh6
Y3vmhUPS5Hs3z3Gaoujcm6lK2ed+6gjRWFhq2j0XUu4U4zY1hKClrFR2ao4g/h91keHROpq7BimK
Z8FPl2QG9wxzvlzOKHlgXVQZJutiMI55IRvud+FiFrKceHqbU+Hu7qcSfbdoWWQnhaJBYwxTFkt8
lU/Vp4AYjzy6Q6vysul1qUnyJECyEJld86NCPO87+qigDQKzcMgLdJ2qCg/zJa9XiLdDL7jelZU/
jON8rHLzDu569sVI6V6F0JXoz2N9W2ja6EmMTrtA3FhW66sRC7hNxSz9UlfJhKRe2dQS1QC7ylQY
E4tiwuPeTbLJNHr3rBe4lBLoSqe5qHcysFoGRiM91CTpRHbdOp8HnqL+WKZzYdiDMm8peAcPQK6E
OJmWVuOIWXAqa3Skh4vf9bMJvOTb6Ey5PBgg5UtnbRX+N733qmNssRWfRem2BqrCZmr4t3VM7oaP
iqihqJSGifY+NMV3KsBUFqlBApfUsRCKJSE/VKp3uvWiqXB0uJgoBxNcUVFDjql2mxRcR2IWdnV8
CFHt977zcDfXwuJZwa0nr9psb4KbDLEnPL02QTZ97i5sZRJGjH9dFHtZHliIc6KT5ykVDRb5qw0r
JvVmUcLxlLynAE1Ku+KgZgIkiGjR8JHvNBcKbynuh8YryFLg9WnZpPRkiQ1I4AZ8C7tSnkPVKD3W
zjhKAa4s8m7hqg64RDJgyIBkl5BrsveLOkzjc2U5pFUx9u7Jqr3xYBarU96qHVDmNpo9CIXG3SQv
JWwS7IqPZ/Vf1I4kN27FElAsKk0S1jTLeBDYpVwNfIAHvKVnyjmmJAEfTtCESZOugF3CDPNeKwQh
3LZ/Woz8LSpdv3WUu8mvfV0hcml+L5pfSBZA4bf7ToAI+ovocquAZFX77wx6rRVvjMrL82uQVGaV
5MndJfG4r1DtiFyHdLJi8Mmk7oiiNCER/eJTuoJnwHekrNyCzOMzyPTtCNuyt6tOjV7wyNavJdJM
4m7ju5UZ93SGXPYbWMEzxoqevhMfS7CNg8OgUEw+TWa65YAPS7P3BlcdGAjRXuEtxgBQh1HlU3bz
quZxQrKPImc1oSUW5TmLpddPLM8qp5VZ/7embF3j730r02SDr6zuwywaFomv2Xzvi0sUrCKBEbWa
fM+RmKjov64WwKPWjkb18p+1yhs6bipqYgMR/W8NmOIH3hTd1fv7IwlC/HbKNCKwMxW6d8We7a/p
RsFOjeQNIzeo/bG6iOTn33LgD9mMxUJK0hK1ctF3FBvJw/lwR6eFcGGpz3PUn1DtkU2z+HhtUedD
iSs5uTHaLDtXdsF6tnKsccwLyYivsAutnA9pGedetYv9pwdcDqaT6w6zMZhcMOhY/ICJdiiIszTY
Ojywa5yUUIc1YLq/Efxs1T/ub/a6UTWtKeG34YEhdTGpah1wOOTVVOB09Jsl/gOFg+zkO8Li79Wy
zEMtsaS8IjhlYIoCLq2TzMd9ukilT/xhABhAJgHXQWWJAbMbFv77ZxWc5Pnwy1jVi+R1qt8ceCqK
ug4tARc+3lQaHbGf7MbEDCyZar0kBNzzlT9mj7N9k++yVUOmPaRaolhHrmUFAp9x8JFa2WEOZj0f
lJhj5tZWgVYxNyD+z2AqlNJ4M2tvZtN6/S176znKaiiDfsOoZGpaDKNCYHsCj7KIh8efCgECNyuA
lTVLb2ZbcdnTvaD+JXGk+JGK1HiNPEkZC2jEylUBkWIHjQnHq2xSix7y3Tkres1NKWskt2MOBZ+9
+4/xFqTbnV5tuq8YCjV3ViQs+YZ9Bqfg50qBTuqfXny2EiiwqcpSzF2zVkGg+EX8hm2RBkyKo/qg
+Hh/CRSEV/prlmBuF+uKPp0HQN5STde4FuVp2QDJQAot803aEvBQVbGKe+AqiwDNIZWh98cV4snx
rh8UNWUjGUcwEjAaXT5rfYSARRhNpNaP2ODsaxkXmPcc3TYh2M7jMCoKFPK81kXGQ7t2ZGLEaM+O
SF88g27sBe/gc4kXTiHXf4AHR/ZSDpBSFPOsF5we5FZPJwqpvVxD3ZwaE9JEoaOiatO/4Vg77y9u
91mout2Ea06o/nCUftgCk08pDM8EBinm665dJHtRSN/IQoGKLkk2OjrTxI9JSztikwXghBgVvCFF
IXL0dL3RS/fD0VoWWRaMiujD4Nc+3E73VyEq4Q946BpY2LIrk6bBK4XjWZdKX1TrjqVhuM1xXO98
MObrRFbQazwqiCVjCg8p4o7B09CeWnpKaDhcBlf0GjW47IYJ9KNdaUMEcfXeTb3G+VHBjN3Bj4a4
V3rgGADpEYOd7gR/50umTL1dUmcppuhg5LwAqc10YUGFPi5VTK72cFzInser+xy7IiXzcQcn9686
9bRd1WllIYyHsBKZK7gi34aA6UM0bjquXWgJEVNQhwVFg/s+DzHqArx7oIBVkA2DvY9uuIOBe+pa
H9DAtR+t2enECKg5QScH6kCEQ1xGyo/gN2nKCjJWgFiVoYVu6meaMqm4myXTOBXhSkKNow0f43TM
HHdZEBneZgcH+eOkySVSfX35JazzA/Pldl7BHI7vmhAmFCYiiDUp4DZ7BAzhvox8/vvfFl5Rl6Lr
bojjSvhKUe2/JFfTbIgZIbFhZGF15zD4D4VfvSlGloF1dGUL9pzUodq2wMqjIHl473vDFNrcFvki
PRKRV75sLVAg3ePix6oWISt+4NavsG4tg9ux0JQbjz0NmXrNOkMEergUSyTiDYaeLSbOG4AxgsMg
JXj/PwjltStKw+GMTbcaDl9k9cjGUfkE4O1NSOM4vGP4UbGuOyfNw9fFKMuQcaRHUm1AKXcrYav/
PwPzq7QMDS0FpUMDcky9OVb+6JU7Vh/nken3EVC3OQDq+h4K6U2JDapzRq1v5GHH6VsFotgN3ywt
liHVAwDt44jEGDIutgNj1RW4Hbxq7wBwVM6qSAghIV1msPP+h3j3ZANQGLu/iBv+Y+y7tMhUyQY5
dTzd5lvYRXwr4zIr6L1mi1yZ9hMN1vXxs3nNlCg7ChbujL+IKxWNa4mXFC1GHIpn9CYCXq1KiRQc
Mt0oUXstjb++OmGDcIcWu8NSkY4e/fdIPC8ITilGo7Dz6mUaCR9iaHCVs3EkmAsVA0b1Z53zaGQn
QMlzvXRqbzJlVyycnLVPQkPFLbtN52MSQGJ4G+y3dbxmjtLc44X3Y+8BtK4QqxyYuzLQckfH7qT6
qXiH+Ggkh012UWCmLyQzlQqGHBaxg/TrrYmQIc+v21TdzJy/OgpQ+yd66n5McSGv+TmPdvs7zbWY
FSToP+Fid3dL8dFA8hgEc4P4OB4hcxawZYHIgw1iK+tMKu039ycPNw1gYINRqJ4CpzPv4pHQBLPN
bpQzQKKYBR64wdKNWJBBlv6H8ZlptbauDptNSyodLf7pqznkKtsheY0MClZ/foKL2ZK8FF3Q7sH9
9Twsd3QrsTEn/W96EFb077BX7CZ0SUu/ljod6OeRN47Pi1jYOhDVJ92yj+eTsLL9EdUhvxRg03n+
0Ek1CxUYPl0tfg1LrYG0XOYeumQ6w7USZmttcrM/TpHjo+lpBhy9xvXTQFkgZCbBmCth38Pgp60j
vniV7invbMtqqnGZquSrYdx/hWeVNFaHfTFbV2qLyjYuU4vwCcMHf1ElvxgQqfK3vx6tUYIGDIio
S8RIyCOlaFaWnsYkSlIOkWWuhGtRSWe149LBBAGl8wHr9gy79eSSI1wzuRF1O6lk8W8K3OLRc1pU
mf8PUafEvCjjCFcZoLvm+lg8ogKBrX4zuMEs23YVeI0FfI+rr4bvzCzhKz9idw8NADb3u/9ZTck5
eXmY6Sa/IzvZ23q3AtJBP76Vjk/OPJDprYXywXMmGySFa8YmWABbZ+BoQ7fTVOFb3YWgZOZ+r6u2
ff0FfV43TSzmd2U30NPe/SBCSvUS2pcN6RDflYm/XJ6xu7XMX4xPCddblQWa9xA25p8pbUah/HmI
XO1wP41zvTtmNJ0ubiiOqqE0XQGYtKuY6sNJ1DCXJrY3kbuVqcZuLtzs1hCbybvkfih5/GdGBhAi
1g/TwP61sU337T9XL4IftDu9EgGcWk6OTvb+1XSb5b9QpbqnO/Xta1CDchBJiuP7lz7E/dVAoyzI
NUBE02QSwoYnBpbHgF++YvxduvXoJuBwdMme5PPomueVVarLEHCDwkFa38dKXpW4VxwTdsfryiQ0
x+xGvbFVRfSBsfTO2f7UnRKIRyriZ/TKjweg0CTLKKcCqW+yKOzcjEmd8h46To7sS5xzRRi/w0nz
5tR5jloVfAqBX/CkkVh/dJ4uIMO0hNvu7Xky0g6kGHLhdTkYnAtQ+YjShc5rVfNDjYBkFoMhYxft
9KxeBFKBJYq0k6R0JVsRBCIduu3mkFW6pFctb6NtKwAmbfg3v/TKzgLK1kBhYxpdwmv+9Y6FPWVA
5ovtvKrmsXkingIB5jEARr2Bs6vGPWf0s/8YQuGvekw/8OzkPvpvudA29UnhDcvXJu3Kk1pJoy7s
gy/hoL75RtG8THLuW28fCpHwXdQoJZXWVKMpI3VNDxk/+g6Y06ytjIWNQYfDurqssJSFZ2dwJUh3
1nNbiaArghjk5K2YKfR8YueqCJwEqtBkoet+mvNQVPAYhNNOXriI+j4JHt3bxu+b2z+tT7sY3htt
E6vC4PT6vR+u0QG9QUABraIfKKTYSeAMNwOZa3UbSrDVmRjxQExugyODr2OBONbPKJw5uCgETfpF
sdr3gJ+DGWLDu4hsu9x/O+qYaMhJRqlTbhvb6rWgsgM/1IHE31QyoCxydzHKg+QKQ1PZ12g48k2j
xWYqKJ5nPlN5vxaNYHc/9+s1m6SCyLRD1t4nzbxasYVDUgn34eGbWtgr4SeX68hVUyhaev9Vod+p
SLMMuSGvrIxf7Lb7vjkir3pmWqH6AfdHRuE7yVuB6T9kMVpA81WDwkF3I0XdYo+WIrZG/+s8M/df
bkr0N36q7ELmkFhh5RkOCdrPR37uxyLJRv/DgFmxzlY702PgKw513rM+bCB39kwzHCM+avakCcTJ
oeNxD5DSP1KejWnBalawySh+zdzOf2PGBTRND4/XZWOBpUiNmDNbtxbtYzcEfk61TzVi4LadrVfV
KwG+x/rWt5tJ2P7FzHY09jJYGjAfo6aB+qRfu+S0JK2oTuWj3emxPfruEcAOuFWaIzIl9HWoRyRc
nEWQNFOhmRNMmeL4mmf2QA5oH+QIznSfBAmbwB40Ovk10/ta0wBtQKVnd38kIJ9Wys+eOFTCIqyO
ZrjJGfbaesBKalgyqscb3vQi6AHgMLjVzANLMlxveynvqMcpivrGQ2Dz4YtHvVpDhy5ZpxgpRqbj
MAvCZ1n/Sn0v6HT+E9I7mOVnMFVqn8itIL6JudGa9ILBruJ9w7jg0NuGuIzzXy3S9Euyla5YeEb4
esDnr/RimDgeG9iiu+SeR6obBjNZMDJtuyjetfHkS2h8XZ80QDZP+G7uTrSDbe252cZLZmAhunon
kfURRv+MCoy+CVwRirWl8I7CcPsWjNAtVrwWXqgaUWcXKr73MN6MjQVbdPWr72dCpABr8+4maUoW
2j5OfUKwRz8IbfRdnPY50bl0fiNcx0KHHt2/+EUS+I5582hOJoVHkNGzXV6QagQL43/U2wE4bJKR
8KiLmi13TTniaS+BwhP5rKxGEY2TE6C0E0Btn7m+sOlkjFx6NLrUDlr9IhXH2MHF9B6cEKosoqqg
teF9Xd31TSSRtZ/r0BQ/GmlJYTX9sLAmIUF0S1hcYDOQp/4g/iR4njIb7/lEOfbphOdItVqq/NPh
kvvwLy9rWsZVXtLZnCcVYJoZJWBmMn5CpN+WspcfzoQGZ8FbiQ3FYPZ1g5joD8Ufiby7Z+kgrE4d
CbwjOlH2aNhcyJaEerW2UqKtoZ+3ZfUKDWLq0eFCXU9+mS+bXS7vGxzEwskFXtnZHD0411tEJx4W
UUjJLGFrnmlWCepVkMu4UM/f4f7OpkD0p8u1b2Q7lOGIOFWtVpbfcqathQ4A/D/0zRslCQKEZx92
dZT0UhenKwe8fSbWzudlmKRT8xrv+nsVAhRSWWrPW2RFIu1rVopJUGFEDDWiokuRAHb0AtvHDu3P
fzPMhf1rxuOJPuldwRW1Rl7iTdR0rmD/DBU44POtU7dhg4TRMyyzq0Ewlgnn07XH/kcNlesxQAgt
5GZvrrNN18j0w1bMii8ozvW4BWApLsqNnR52yM5UmW6FyxDdmt8E5WdCIAqP9h1fSnSCoqPpR8Kg
8Q2QDQP5msJtUZSjVC4Ciltn/6stIqTsri+6q/GO79E3CVqL0UOdqsuJVCm8qJ7dc+qeJI8UluiI
376WFMYPzLEyc3FBqAVUQSM009OCBLHRtWNasNX7QkLXP66SC2kYFwSLPimMxgiJxjllgsG7HGqs
yFZFhKQFdedUuIE9d9ZLeUzyseeclcvU+ldolJTu0upbAN2C9Utef8vBz/urnh8W5bJYaITDTaYa
oZzIl1ecwetLsLft9wsv7bU5k5vTG3H0BPt13NURcZ6FiFQtPm+k7gjwP18WJEea5PvFj8TdcMn4
ONlWaYq/4aripkECyQmOKsWM8PqvbCDZywYaMlwvQImb6+aOT7Me22t6rzjKDwHAS614n3G8M4Fl
uO4tsS8+Y0OIYg8sUmcyhtBalYg7cSExjgBJFT7rTVUmThTbZbrnVJTav+M8hXR3505gZs0fz/gl
WzCYqwkkBdEJWC0x/ByygoSpAGXlHU9mk3ipZQOSd3Lr0dV/BvDIwNnJIDsH060monESL8wYw9s3
iiy1UHVgUtSK55hFJvitLugjNnnKvTtBAIUUVnfyQbB4NPvRn0hDVKxAcI8UOUUuU33aWETf+5Y4
rc30p1S5CgOW/1Cg3buqsLBj4aliYztZb976nbaVpr57hF13L0bfleo1AT8tfRfRiFBz2QkEx8+J
TOAZLeAlHoLgidNCl/v9MI7Ed2rlbVLPro09FnEeA/ELTLr5lveFrQjfmt9/Q+wya6f3v8IDG/NO
5FdZs58LJ5nxfvQo2dErJpY+QeChmV55PRl6/yMfxaBm/PAG9Pwc+hGWPPH2cjIXnc1TpbVzVQoL
FNwFftDqAqgaMrmgMseZTftv2LhK3TjFXi/ch6+4GIPCRazY8U6qI9x//poK9pUFMBc2QT5bdllb
4fxjxMLUy+4QrE8+LoKkmReFDndBhsVtb8HGedaiQzdo7WUFZy4ufqn9n/hVMn7vxUAmxsGE8irX
VIlHVUPzd29hdlzf3RG73syB6i0H7XaJWGospKPR9H4qwTqGof33wt25Je7LYnmKndezie8cc4P5
RO0pu6MmRlbqojotK5Rxm5Sxmnt5fQBsS5sHPUxd2ZXLSJzqarFEHivURZ9dc2R3qLFAfCWPKKLg
vwp+FcuqC6i1mHbu/79RUmeYiOp4VwN4VychSFIWJ5LNsoqEqjHGFjbYEUDDaGhof9YxcKrJgsXK
Gtaj41ty0QhmMW9pQMSg0uWdmL7AnbcnPHQmYnRc//9NzCPCCYoQbNyQDF9VHpf1AQpSVkdD2OGn
cvRZr3FbzifHmBqfeSN76wx1AF7yeb0mbaxiUzDy3EKkSpy/oliyFSBBAFo2KUCgtfuIuKvkhrVE
YCOjKz0BC65xe2uzPjjkyNnx3ytY2BDaEL+0uyR1obFpyyZon7Kf+LIOFZKpvpy1Hm1pUp3rbtd2
HO2PGZmOEOOwlhppQm+TXYaR6fU8emUTshk6VrfwO9Ibfc4FaMKvFt+0I3UGEOouAc8CEiGMjVod
SV+O7fA1Uh7bcwZ7aVFyo7EtNOw+4TulgkWb2WRpPUbZ1ucbiC2peIDsFFD3YLSACQSLpZ8AvKtO
7AAdKoQq4NBKd8t7u+dH019nZ3R5vy10kRGRlCK0j2J+pX6Kcce3MK2HvPiIYgg/qMK1A78v++mJ
2JI+7YzVfFg77kuM2idTId9Rk0W+S63lVuSRtTTIUhKpNkcCRJMwieeNn4OgqQeeqqbQT1IFKQwp
gLacv7dTHpdJ8IwA4GczAo7nHbA1/TFy/Da06xuD++s/4O/hlWmkzsJiD+szvIMzsl0p2geNSdbG
RHMBcPAVBPDMbApThdsdHWkvhHhFWSLTdERHFGIHHzS/3Bbp3+TSERPTSpEVpWaO2JUDRn/qdtc+
PW9FJbjvk7FRvEb4IVpbaN8a8tJshpiCxvEYqmmUEvWr7F4zwYBXrp3WmxtmVtTu22UWtA2NTLZM
qlz0S6XQ2BM5X27+iUEnDHTkBn7PKKVtky0AS2eXF6Wy2S1hnbLX4w9sansvJ4hixMi9drkcxUro
wyRWZlrzhGH0zEHFAd6X7D+fUi0vySJ1+05/Dv8ZatFmKHiWoYwNTBgiSC/sUolMo3AgCHgT15A6
zEekh+h3GNTXQGLXuIf/mfOc+4ct2O9P36Hbsmy1i3r+zNYEElpfPeOmvrPtO1BGfmfA0KzF39q0
Dl/6p7lRnZjw7/WKUC4om+FXTF8P+qakmnxzhkFTwci2AfXdN4ozCJNpm7S8PMrKEvvAApzpyDz4
TS94luD+GlSgIePwFfNTeOanbRolyGPys9ZoxWiFbYjP+fJTxMb3WsDuFA7zYRCNf4zbm/jOuLwg
zsxrI17AWrXXukPcU0ODdc7I7PaOIik2VnxJiM7NjnWooaALGyvDCmns2AjSiXfp38qlBHw9PknO
B03KV4kJ/Nh52joA/GM34yTW0pwOKFPwIVd9lVKGpdVUJbDrS7Iy7jddDehA84YdW2p11pSbe66i
01WEXK/7bhFWVu5qbok+qw9oAy6jJAYcY14wjTl4AaLMs5+Te2Cf+iG+IBFa8bmpZkSTNoz8hcHh
nN7nUoECImoSOInNrWnjP/6zGFZB7Fp/eXB2z8DFd8wTh+HQIfvy0PDX6dzxc5MgxqYUTxiHcXyL
+h/2A3TqHDR70WyBAjZWheK2dIBro1koOu7jW3mPZ1sU5Jx5sAkUTwlWhM2xlFvkcdLJQWm34Vmo
nMeMku896qbx6ATwFpN83a0o2/q0HkLKGPEikEUU1sDcnMU9XIpr9zzZD4Mg/HzkkBjkBd74RaxH
dbZODzB6+rAR/FjmFctQfZAcaFTDFZjyZAwu+Gwbz1adJ4wLvfF4t4UTwmDhgZEe9rPD8wabqOVN
uASNPr5RAMFUTxCC3/ySG5U0im2mJLAHLsOKUx1Hr7kZU1FKUaNtQphna2gYvJHXT4x2OTH8IyYz
R1o36CUIVlUD2n4uLpkcUkneXjz5IUWSTmB2/YEaZHylz5PshXGdxW9IfBOaQpBnFqd3U6xnzBef
eGDPd9HTolTKk8btDL7NwA9YXuBPrfynDuYCWHT5Wi0KgfcCjUK4VOA3afOdOYiiKyO/hjLGEzQD
UrznLg7mmQOMZ4FT7Gd/LRaqxesBm07Yzfid8dO0zQVW9IpKb8dboJZOQMzxWyOkJWw0GI2HPr/8
39wDa5OvDa+ZlI/5uNFNH/EnrWOCDaUzQekrrzEgqkJDTYkiRfxCOH5nV8Vf2tq2G88fJKydOHZb
2dqaH8Hbshh7YXnx92jJMcr93MWXmTfi4iNKW6f2uQ+zRnlQ3NCXB6ktVGKAvtfRu+uRdZ+Oo/Wb
Ikm8CSQ2vYvnX7r3rDAsIXabKK0Mak/vKS+CdHm47UjmywuY5kcboupJR3JF2OmFl5JmSlOPtKrL
YCHSGRLQlvi83bRmpD0/ilitP/n9VpGpt+qk1DWN2Bl1LqZ/R8VJdIJEx99M7E+ne46l+bd8dGw+
EUjWOQPtKhiO1BNmghj7SGvWqmcXFjIJsF0ZRxFUJxUTbccm/SOoGV22Xury0DRxqpmL6WXn+0/N
jYU3MAPgx8pSHtKdq4SlRGNvMOK7EKXwhsEP6RQLq7qFHflSJvPhu6yA9gno1LdUBNfRe4IQ/bsJ
uq0ZIpkXNQG6kwnv2/FYFFIZoFRSpy4InKPt+aUOBRFejLZIgCKSb7fhSfaZzdFCa1TLSnK9pAsP
Grq8gL4E31aRlRX3uQ7vi8N8Dm3++AEvsbvZZ132h1KwaUl0RPwh89jYhCKYerP4/KINNoIhz+LP
PMM/nPcCpcELAZdsVYGChwmrGjI9lHES57PPhcbp+qciLUcS9P5wuH/h+Tp2jXzaSpW7pEu45S0q
HFdyw0sRRz4Y7Xz70PxDdZpli326GNq4rg+Vf7ay2km5blIsk3HNGSHhTHx0LsDujQDFdFiXVqva
n6XqmrayuYQ1Ohavo0YIHe0HzAaBvADqhz2pb+P06xrdskhYvZqF8z0qHIR4cho2R3AJeYygI5h7
s53nB2LqhSfiHMUtUfUtQEvEsWwVMk7MPlPt8R5T+1A4tO2a2bUD/4YF0TbDDxYi2MVsvmbG0gq4
YqVzi9x1Rn3Cj3TjYwWZZHnDER5PcvJD463bO+8wFQ0MZTDJS2tnx5MJERBkyJtX0nLDztOvk0uj
8uHnLB7RMZ0fxyen/SGp+hk4yIrwe/rn7p0Eeg2OCQQSKfvxzioHMcOULk15A1Hr44FPyXoixoqT
znU3pwSJ+GRGbCf61XnU+GqXE5x5PiEMRE4YOUbys/TUKVVlDoXm7l6tT83zwBTgN+FEh6oO6MT+
NcZefv6X6vNjoa0nWSdziX9sbyfmf6AZfMZDgkOXs3h/Uxt/VLjBPY/4u7IBHW3aT0s0UisgBudO
VAug9/L+CtrAqvtP3Opwpm8NEM/uI8Iz/GSH6WOGQcvWhcI2Biwan4pCEfBPNg8jHyiXty5rVMcU
oMrfPchbq+3EWqNo7NgzzkkePDQukpobn56uzMwAKD1cBErCZYGmKjKtAFDKjQYFHXFdPjtMUY7E
0/4OjwtYaKHOkeXuRrunJXHH4qbYM7EiZXtNEwgTstmI2ZpSgG2SXwe31Fhs3N8u80nMrVIjIyOD
nXGZSF5RqAAxeKivRtQB+Ze/1NXBYEj6GNxlGzdvKF4uiYTntRv/FcsYAYriYmTPrl/j8fb+CjhP
GZRRAZuX4WmycIqm84RJyBOhl6K0f4DgtEx+XNe3XqufrSlvIlhGZ4CyZ3oPr8KvlSjwMu1xRzYh
6MAeUGI17NX+I3n2i2livp0JCZCnOZSgNfHMmvp8O8YyGmyvuvrWPtDuVhi+u4ubDbi98hBYozK0
84grHYAHuNadlTpr+sqHWbcx/m17rYUt+bAIfmvJHXVUJEhhI3HmqIwWlohceOXN3qMaaLPJxMXL
opDKpgpOOFkmSJ9Iy7UUnA1g0Rqb5vQpJ8LRieeJEtBi0EdU4Tmi0YUDY4xfxs9f1rJVvG2cq9bC
Ak+odwroYdW3u+P8NmpmyrXg9iT4HCkVM+D5Fsap/wa7nzYhdJGUM/wV7fFgMl33kQO3Bj/O7FQ3
D+AXbIFPiRTyiJmI28mUfUe8lRBsD268AKUPIV23vfLLhE70vCY2YDuOiUtKRQfRcnEdUXuQPUN4
6yrcM4KJzG8d+ND+sxQxIEYMvmBi/BCrqumk1ygTt9GcGLYh3nYNzN3taO4alC3H3S+ZNALFcrX2
ZFO/a/BZLrlf9K/W4eKZFRZctG/xGrQiPPtGpVyyQtKcOEb1VDtLn/9GzRLxVGUt+m14J5eqJsJK
Q9qn7vehuZqpsvK2FiMZ/DppNQHmJVFKZl8hmDymCsrvRavRHcuyBB5U6/edsAEc16RjI3MsfFsb
VircpmcydYEeVlUhk6h7OJVothnE0VouBaEm5phSHnmbRN4hjmu/VGe0dqiD6sBzlfsAB0GoS9uO
SZtdXkjvq0uDiKFW7/c3MC01z2ddd8heIiVNLO4WYBjrBzzCqufkHdo+7NEjCoeKyIeW8F8Hky5L
LYFw1vPPyr3agPeg9yV341x8fMIaM2K/kznIBexs40AI/5lYCGDjAFensVtCR8yqeKr8Paa3w5fF
2sPDdGk4Su7RtBTWz0O6syEqBOVTKesoP9Wqfyv+Yv/AQxfpDGZBUsQ6KxsssADRAbKlwO966kjO
uMgqr3p4TXI0Ed3Fy7exKZ3GlYUayYPvkEMjxtI6S1sbHFzp8XXridPMWI+4ED8DOIjAxuA8qk1g
UggIpJxN4riJV9zfa+5ICMBG0bOmMI1apXhiu2GSuA+X5M1xNjgptw/bxI6hCQAwF8mUHZA5Xlnd
Rg8xG7bDyWX0TZkoH2HwquWxr/N9XunnIvdSy6rjSdiAMNITCxxeYdYNJyfD4RTxMdbpLDJe1dLP
82PjP8gRqreB2mwOQUXbVbbDrkkQb+wzePFwEmN/kVc9nDn8yKItZLcGwGAsh81KrqJtBOsX04v0
Cyx/TxCmO/ALDoy9rXiI4JVcjWQWdafuMF0DtUVQ/gfhRsETV1LkpAg1/q5PCKrl+OqGAgLL1EO5
ohcWPVrVuXSus1BETdrh3GCKVIlRKAhqB7XRhPqHat1gcRvCtWvYiNl6np6j2U96UIRJzBLF7dLG
6jI8pLqVlzVPqwy4fwAW/kkPBK3g8w+hJCXAcmV3108RO3wWrW3beOdP4y3cIlmS2QJwxtc1PUZL
C/4huYVLCfK6zHVYRVfdfBDm/fglzsGCAtMU2Uouf8zjuuM1j9VASlpk5dAJ9arA9hOEO6xUkNtJ
aHVG90mNv3RgTePgBeA3yFtvobpxHY6RnUIB61WqrFWdwC6T0OqkPUmau47xzONj3lxwNZJCdxrE
Th62+aJXBJPZTZTo1n0qHRD6QoN1lIjj6665yRoz8uwUafzNcKbOy7uamJbBn8WneeD0WUFIv2Sr
CLEDjooeutrlCuJFe8lSXlUh5AKrIVT32O2DT9v7aaL49tVyxkYFiH5yX3Gpie/5VQt0BRwUTBKV
xvxbPe9bYAc0QcXaF9FINGJ9zh3j5UcQhPLlHiijRKodj7LB+njGk/V/xLkaHWF9noXi33hrHbST
cCHGWvTH8XTtWwWaba3sbOieXM7AurWZvkUewnuARjt7whCe3oSoJrGpbcFfzF4FG+qftDXX8adw
UPOlbC26+V9VcM1wgJP2kV4KdtyiL4CbPw9su0EuV8FEBQ+Rd6jubfzNdCGs7jD5u3c7OGsAYItu
VemaJpZXODo3mAO8+rgDTTUFn3J0ax8b03CzYZO/WYFEcNya9gRLrCXG7skvQ+XPaI4E+Ko8x6kU
ZhlOnGoG/+Rn3SQUJ+Jt1WcqfethvdIsKg3IUmqasgrlBRSe3CiB5QSLjyeZ1pcB5WGqjG49cheH
7b9AQxQcQHmfkNsAKhNxmOpkrU1ZFRsl/ea6JE20V5JOYtBljxKfUXw9onm8AVhRLo4mmTTnIhdy
pbZxJPPe2t0548Ds3+k7xoHDJxTBpuAOAkw9MxPud/LJqdV1ghloM5cNcS54Qm1+7R7wI1LVP3VE
G9I/lYG8NYBV8bbtQ3KYpSSbHl+GKKWwWyFfVXbBVFu8uAvX1TESquPWHEWAP+JfdvyIg4slsop5
Q3awNNPoQT85h+UwUx4HN72/Q6d5cLUO0ou+V5kgfH4wLj0vdMfg82KFjUkbrFy+BPgFpfyZh8ZP
xrjpRfnENACUK5eB6L+FDDdQZUzIr/zo4v2FbPgm8OSTq9r4V+ZsqY216kh+2j9k/zkxFtpY/5L8
mvppqwlhQKF7NdZGeMiiSIvXttXQhnVF3OJJP/qaiSc5ua8djTfGWDC0B0BfZPnc+eiiXZnP+QFh
62lxQLSUd9YfYVY2y9oB+NiHulhtMIKNmRU5lCrRaH+Ygvk0PxOYbe7BfKBhw4pqao2KZd601Pq4
nXbd5s2TrDYocy7P+fYa2Jo6po1IRFxEBoCR5vB+5WVcQ5AplQAg0C3SuBpdWjI+CtViXq507CcC
ZZdpWPm6XKDyi4J7nYhnMjBhjyiBrQRNikaOajPVhnCuiJ0S0+SrAsygNycuX8JkfHnNumkaBQ8A
h7FVDYTF6iwHdBtHD2xQsgGG2rHoNJk5fBCNwAqh9eQ4L7RB/BwxeYeOd62SgtijCySW7Kwl8+B5
LbP9NzRK0lOZt5lJWbztNuqNO/mLDsVOytqCOi62iQerCYMNJzdVlU2Wvu9VWw+nLguBXpfTDo5f
WpameXJQBKjaoBZ9lKY5LK6ZN2vCDOWvL34HWKuZE5jHuTnsLCDo/2ngJkkQYQwKldUp2OGzjEBf
b1RB9sy2gw8AcsvWHilRmh0UeDK3QeN/uV4X0NRA9rhd+2FalkK/TJo7w05BiYJHkwtePwf2zDU4
giBrbX87jSJNVgdh5Fpxds2+bDMHQC0dmIZsMF+KB1qD39lwOhXjxRfbFVcMF9B0FBuVVqg84OHV
0HKoWAKyxQKJqhri0X1h13n8DZx399vxGfeJvamixDr3aHcg2zxd3icZg8/0RwNtHhNllonrf94A
aAXfrVSsODCRbK/Cm8fy2LaBteuBSP/MuhqFcPkbrgzx/t8jWCMTt5hY1/xMDiNt641CUa+eZo6V
MKNUeslAg4OF1A7DaO6JNrj5j0DMSBg/8szgEh2ar0CykK3PCncEywI9G/hFjDrGkFxYUzl5Vn/+
eBPM68p3EH4a4XJLSuyzlsBOESD75u9jc7SoPewRo+XAKGRa04oYzUV4X8IZzwE+FcJC0ZqYsawY
+9b+Ju9WZS53YEt+Ap3ektpKCLldM7wfFWpLBi8Ypvxrdy6LZtnBoh2i3P+ReGQR2HBrIzwjCoYj
G6Sc8P9pFAxg2uJk3W7mWJrndQDZUqFCjZkuJJUW74dQO77vKpdkY53CVpyRGad3qUccr0VOa91a
BHx2p7L4A0JsDS84GeyeAdm/PJHN6PkX3VaJXsSinpd0ZGeeT2pybqbIBIeopTl2Gu3kst6gKnOZ
uYRwG9PKyhEJX8YgIepg22Djavxwxt4O9W2Z5H3Bh+lxmWvg0JYLYGnQRVH37zZ/qb3GwSRrQKtN
5GHz30xSn148+7jYmgW4w3vF8Dm2NcKh9xJlNuf8M3VbcwSShVzdIbaA9vHvZv3zg1BghLwWnFDp
gkdibQDKmuyh5JAf6sl55ybJKcPHPVrKZ6HuexLGkxsUtNHj4DbsKcsLLMvvQvBbXkQtqSGjtvkH
v70YT4QMa9uVMlXwx26dXxAJHQQ4dXjGUyiBjZaUCHxuDzp7Xmewdejq7v/6N5GOhkszrfMDbFVl
X3uC8RiYYphDeS8YLoWiim996Vj+l2Rr+oNXDvZtRPUDHeCnkA21gJCk+dVNhqt2gWgb/gw0KdCV
07ZZVCjbk7m0Q2wzHpgirKvdEc8JM/RtH3PbvES8szKqW63izBdMzHlw0e/Hqtky25SAihcTXPfA
SbWypOkxH/1PoYd/5Tu2b+S5NyAsc6v9ZrBkDRSVYFDDtFG67liZQqhV9HHllUoOx+1KLXM3vSPA
gMt0BDn7KnLYOIyzRLoIGYBUYYgtbKqwmSEGJoQ4OfVdSLLButHgsDOalZSx3ESElOmUdxZuZOzu
cybuM0hBygLFcWZULFfPq2myFdTlxGJv5ZUY4hcuuROfvB8OmF292yu42b6sfRkk84OZTnV6cwkX
dZIkP6oAsMzGcqKT8EBpFqsCSxvVZkQofuaMSHsUO1Mbd3fyoXVChNo6QWysM8Gb5JIdNJf/ZZsy
T12M69V8rJjDVn9++ATzxa2yaXxQAI3MKEaFxcmRtzwMiPD6pBOK7AdkpQH7yioIq8C+ztYVIVQg
pXvMsM56xdVEif8QaSqAgowjI0RtG6N98siWXtcBF52ge2sTnrTob/UOnszX0aWqAVJDcgbxPXwb
wc6izUk+iXWndwQGCucxJSASGO60lhIviDjuV87X++K5OoI5guwIJjbPn6BWOPSvBfZIiKx59EKg
WYacVmXhpjz8VdE4NrDDHWmPuw63hg87KKjgxhh6EtY49DFuwqUgMpscrFkQ+3rMGE2Dl4WNVj5S
LoMTDf1C7EjNBIJILy4wH/ouhMH64Ao1rDOI+kdm1LYrl8zhrb6vAysGUGwSK9UtBFIbAtxQINnw
TroKqsAmJaUbJngOA/alzwu5Ds0pysSU9NYmOvnwHOQcrGNlacme17V0EPxQjdI3LpfZornPpAwK
5AXLeOdwgrMGYhC84sEQxYIZSfoiinqnJ55ztH64zysxAs1OYYN0MXXkQUbag/GlkL6dsJ6zQzD/
+3ZBsFK1vyYh7oXlGxlVX4x2I/cxqCoiI48yiewHQCORDZQorC386/aJo0LFBKq0Cpmw0a9Bvk7h
qk9gSCm7BNfn3VaxB+R1kzogf7bWu9K1uFPPcdLx/L/t9r20HJ+FgFDaIBtm4yxt9WqirjhB3BCo
tuZaJqOkxPFmxaFI5Yu922NnG+fmb+Q7VhjF/eHVmYkVNpcErqCe2YcEq8IJVgJv0FMxyOU2A8TU
DQHrFT5LEZLTRIjqvug4O2S8WY+SzSyidFreuRrzBbFO7tCHFeVftqceWv9K7r6C+L1Hpg+0XlMP
HG44HWqsCjpOuUN23nXlGDD+xoeGY9pwe+EKgHBst71V10xS/cK2lindDVvxBpQ9DnqlXC58wG0r
Iy/zsXhTHChQdXE0uC6mYN8XA7pPEr7WcPYZHMlreCw+zcSth5Od32wy/owRJ+g/tz6gtr7PUtjf
MdfF4Vn8kAF7H+aHF1SmUHfvMcaJOPEs216wu8GNjn9LcphXhq6CIRqSfVsIVUb1pse36jDBCEHV
APw/gJPo4OVNgiLDFr2X545rf+1HrTP+70Ah69H4U2p76VSkV8NFDLfn8tK+uvHSzkwBi/Qlu3h/
f4MPy3BliAs6dvdgHPmq10BotNZNrVtCTyTHWbzSqgllGNS6saKtT/yq1FXj/ZpG6mcPwynHsbyj
KxRynngG3vsrjK6f1bs4qoZ4wrDo+hx+OTZRMy753f20CpsnARAram0ZvSmf3Ll3xUfQw2yLqFI0
d3gILkgI3AwNKX5z0bVfEUb+lhnWg/NWyZ6X6SLwhys6sc7EIEqOoe4w8ZstapdF01uHTfZBWLhs
UFtLNRdIZYWwJ5Bhma8wHZKEoP8A6bqdQyvVgRuIJc16+L1CYxjw/jncsmVQr1Rub6xU5M138sKG
FM2btnwS+8qQi8VFhUoPAzdIQXjL0EfPks1U+zm1WfehOoKendRY51oBwqw8OlE5cf1Q5WX/9rZi
2S18ElrjRpMa/DPK0lcqh6UhKEC34n3h1zwiitKcD8oCRnPryK1XMtB0g5DBaO4jTvujtLDx6fg9
/WFc6gWYS1qJDRF0mo0ZAaGATVfFIOXDMpTWsLBO3Z+hVSu1h/LqN6hXHqXy4/6POz1RdgX4YzbZ
IKS2cQe8s9DHSted1Olxvb7gyhrj02iz21i+0USj5PF52c9LzdIc38NZBL13F4HqLV7h5MqwFqrS
irzaDIPzzgvaCxsE/nGS+kFUauz4eCSkqopzCGuUUJQ4SEXwJhsSe9gb/Gdq15xNz1hGEdZfa9nK
XVxQwtja9b6Rc9QAwLqzQVSa7xSVMF7lFyszEqmLK8vA1IlktFLBugzFxCfU9txvGIEzBCQHKSFi
wy3vrhjw6ZHmmiwUH1uU6Ge7V4fh9NO7aKgd5ZOaesXN21GHU5z9x3U8JFazGAAN7Yo923+hY3uy
K/ksNIbL3XvFKldKpWqXSs2sYaLs9W++8zqHyFLIJHNC7XYjqImt1KqRQV/JebHOYgKYnKBEqGcI
T4G6V3K0Ci4COcz/xoiUdjkMlXQh+DQPXjboyth2W8OdDSWDqS0e+BbLqmYs4HV9cb6Gbegohw5a
W3KuwgKe5Nz5gD49jc9zCYSMaD/HWC6uNsYiy/jNKf8fuzq74vVxdTZ+zuJr8yCLMbQDEBhp+CfI
V7sosNkidwdDrTaBcKJYbJFGv+D5Su42BDluiBYaa0YUs7WtJtiFqWpVjIcmFGoT8p/6/d9Y8J5z
hi78413551LnZURk7mF2UomDXFifM6/8oLzu+7pkHsqjfud3CDeAlbfr5Z/GQc2KC1RQIWKLSfG+
wquWBx0zYvESr8P3ZgF9gx3uO7Yd4VXh7LGquW7tBJ/blfJPku70mtzP25/5oytkFL4ylMK+bbQn
9MxkNX/PatbZ8aJBn9Ry0/38yXjuGSjPLhNIcuVIQp4NILLFCjYBmiXJwlngTgpHkenGcNbJYB5J
YBcyz5j13Zx5IuVXRsOv8AO8uQdPX3UjAc586gwlJmUSGn+yDKs81n/nSYwtBLNTOuQHpE73ZohN
wJyFmqYj5L18pci8nNy7kzO7tSv7ZYgkzMHxAI3JPY4fkECBFyN2CuEuFGnIoyaJUKbmWnKejGHm
2Z2Nj3A4axLuKcikbC+w4STkAU3M+XMdsx3YmS5o3DDMjqZH3M93RVjLaKrk9S35WWmGke9vIwO5
010sc4bn/d06u5VHWr1k9b5zpjErAFN9iyTBV+NgyZSCEynRGYETDymZSYHOCIumAkfPi19dxiCF
z4M/c66KKDSFrZcHvoJTWnCDuBZecwjrH1DwHLUaFYprBRGkkLmMx8HUlcLI7yLIfpdkulVlNos/
xpvJM6yoxCunie6ZWwvyIB9PqUZfs5kON1g36LBi80NuZHi6BWbUMqB8bYt+wv81CSDDbeU1tbC/
NlPpiAk7PfvQ7UkapFYYiLwQwbHVZzOvV7E8hz6WzkogMg6fA6advKikkFo9s7U7AaYc7aQKYYDc
J5GWIr2jhAv3j5D+CpEHebsTdoQRsFcmkKeqRNR7JSXcFhQ6MkZPNB3SUQQiWu4H+Mem/bA/WkB7
qskIMLaB6j0CsSOet5iBgg+vMcg+DPzp7Wzt4owuMOsXIrIfjsDNgSrvmQqcDXTt1jzXH0qVsUHY
zdwuN+o/bh8MhwFk7S6FwNd7FK9fSa+ZtwPPTUBdeqayQws/LN8ZnMMbZ9cwThxpCgXuVivKOk3u
P+t7WuoGBtvVg25WQ99BM2M5Pqg3KjiXavG0oDbA0l32f6GuRNZhO5IyAC2eV+sbdDjl/NqofFVg
/MQIcZeyBhOPq/xMbJ2Ig0jxx3tKI+BNjbsCFs5YCxvE14R+bE6EgOH6FRQoXOgGViwuxqJ7kOqo
maXI6pb3qAAmqDFldhjbmnDW0RFTPrbmt1xeQX2EAaJGvMRJkXYv88UOXgk+gtwzuqjPsqmjFxtQ
DBXsRpWC579ij87bNRMYpu3BVhRaOGB4QnxK+owZkzh0Nw2HQsALUXvUvs6/l9WjoibGv65wnbHo
9CeccZryufumXtPxJezQ6xeb80guq3Ck+wvDgVGzemqQrEr3cKYRnPf3397eylp8yBqpIdPneWeU
6WmxKA7qufvd4NQSOOE5CT1zeJzaXf5v/be1QEBtEYzTWjM3QtcoQmpnZKeeDYMATvH0VIFpMf4s
rg4yh5U9FsMnUml4J2yW4desTylz2WnM9bFhx3WzloPjqDl6YCZsNnnRxeLRpa2RwJrLYDzbjJGM
sVvyB5SDNIi2rFpIjzZDRSrImqQ4A14OPPpazw0k0bLnxt7vdD6pRnnomQ4/TOL4AgIAAIa2RirL
0rN2il2dt9p3+ZIZuI1wXPmrV2ujB95GyLIMxToCy7tWoifCUJ2db1lgcGMOUnoHWcGcr8TweSVs
qbJg0aHw84TVcUcw2zV09iM/4JVSyJZXWqce9TZenYUW+BV520sGbVwUcDE8vn2Sl2YpulnhAITH
aj3lKmS4uYayWQVpIoxxRTbSoBaa6ivoFgGec11GLlRydK/l6mevrUrMWjav3ESQYWqCQRFdUEab
+74aibCAN02DlbqE6VZzplLM9O9UT0T9NdDaZOWbOwqOSloH7Jbd5TN45lJyX4kgsWsE/8XFD3uT
BlVjE1I/LbhBo7orlNH7PdR1PinwFqNw173WVEYtihkUNxfDY98jFuV1vZJLc0UV71MP2FWCUY4t
R2hIfZ10gOO1qgcdw54rcndYaVerRdfhakpuphlK4jQTWkK3ZPPjRkiSbkCEfGxYd8jfhrrjd7dR
wwN2+0gUizfRsiju7yPpiq3ABiHV7vSafYJcIwgOrimuZZGgmgnybLsaaKjlslcqpGzwllSYux0a
2HpfU5ySNK781JIxOpLZtmeGih3G/8P5TR2ZvFzhinkaVdjawz1B/awZsAJ6cs7U5XA+yYaSo9I9
KdyfPHRSk4TgZNB4pKAeCXdB672v3ez3XHHkHQyVu96BQEhQ1jpYATa7NzXSJA4b5hzkBlxbLwiX
5Bg9dnyUCL+0wZrykoLqVPw1Y30CEtQ+dZsa7qc328Vh6+O0jqkMfSbrPq7nXsg1m3hg67IZnaDI
rkabUnI+mMi2SLYyoNsOb+vG4r3Qh5WBukfy+42DeVFk+eJ9QGZhdvyRTUkaw86nAJPoIsGY5psF
YQfZVkagaHFTOpCeZH3y4uzNG4u1JuvNC2GBUxZXOwYjpX0zmOEOI0isNiWeJDbT+E+X6Nd3FsrH
vT1XRrfMJz+3B9BvoFzgL19NHD1o5ufgrqAed4uMbtx2dkLUbLbSqBIXM4J5QUxUC/KGMy6ENLol
CJ/RkblB/v8onEc28EdQ1STDYMKktD2V64w6vqqyIpa3ZMq8TYqrwg2ktcMSbXK7sBQfN0n0ooh3
MZr0ss7v/z3kf5FXNasibu1DYXMAbIo1bQsqdOsRlDjROC+BYGiFlZeZYILY4CjZlAJjdmPCM4H1
q3Wl5uXndEFZvgSP3LKVTnpXTt9S9OkRr0XasLVkJfHUDK6CQvSDZKUaNGEJYhurv53JtgiSSsdY
T79CXapUFeW2W/Wox6PGdjSsNdNcL5DBUxTBMfP2OflFPlYAs2XdQ2zYkY1Wps5jZd6vIT9Km8es
AVGpGZzlxRTn1xzZxylhoZMpuxn+t7RL93552v/GdMMejOTBbjSIwp0ewMMUSR0aiuAWPLHrA/a2
Oty5QZYZC7yNZ3rW8l/6QSuY4LWZamHa3Gkz3MVcqL99c3hmLgdyHsS4jQfHOo4uV06JCcw89i3B
JYFxidzeen/1Lyjb3mmuLGDW1a4vBdMlL0VFcMwIra+GEOvBO/KlXXcF5dZYIUtIeZIKYkE/XzB/
mYQcjw6718Bp7pc6X1/+OeDmJHNIEqXxtgp8Ks4avvaRsQ+yLlOY1zPtrFWsnF3l0roldQ6TiBPp
efOoMGzKJ6l48nqg1FQLKX9j7y+5J/UllsrRvNU0uJTFBDJVcVObfNUZVxZCBNGWP18d7M5bNKDf
mEB1yXuVHn+f5ZZPbPPeMGgq3PbQ/jxngxHaYNZBlTdPSF6DA163Y1XEt2vCiCO7maou8Y6gFRJx
Zrz/6/dAAGzyEQVrITE+vIRl7bDIMbO0unB2bzFQJrHe/nssuCHohjLjmdeuaIvwwfT8tzzZ1s0Z
BCGCwhPgP9p9LgSwbNtbMLqN2q6aeRVXFcTSakdLL5haciNUkx3u/ZnDMt959dZf5Fj1PU80CBYV
BHqynPTpgejrkjjCH9rjbsX6vgWyKiOif2oMZW1+2kZFeYRVxjrgoqfb/bAL1wRP9n1mAkQ2GgMt
dGzdv2gmjg/4zVevX7C7qX1R7w8Fgr8nHonO/yfGZzQgNMYPOmflE/71D0rn7u/ga3ARJjfMFKTq
+vnY0/wAmDMk34yF0fBw24QNDQ2BdX5LjDwdhaJEHkKclbpcHgZoKA11OT4oIB6FKVmsmfTDTR3O
+GBpyOs4fThcziHA+/wrgv0mmOkjoMaNPcxldiPf/82IZ+7xfBzhK0RUmy4mR9IZjy3q1M5m1PBf
rk4TuasBH7auv1TacSKlqGZynPHT1tZGOrqAzm7eqJSel1pVtVbcsOSDPEXWvdJhAd8bgUySZ8jV
e2s7ilXmDYKMo7JN6zw1gV+kWbnZoThGzSp4Grl9iN5yziAr5Op3TuFTj8t1J/fmAK2Oivxam3AA
Yl01Fx2X/rC7pQVZieR62RrPHefcYYatiTN0MVGazcF8euXgPAn+t/xQ1ZHrgHAT00LjSiccNq1F
riF+hc6ja7ehlVZ1mZeyc/MaO8R0qHzqWOwBTgJuHy4ykXcZ5Stdj/shoEci0AMH5pxxwLfEqKmI
bcBnZcn+/vStzOIoyIGWsWhMqq4nkDJDubIzf3fcYl72g2NFP4Cb30Su5EkQgyhxu6SxLvIMC2FP
Dd/z0SlLXOgpnu8XJZNZLwbnKWVCqHJEyR3vDblYVZyjZyH/4KWJx1Fjq96fbvh2WULMJsG8RlhL
4YWV/LjWDPNfGq5oDmVAPxa8DPG5bkio98k56MQL9NtoUIoRmuGw9vG2IOpZXCKbM7pJIP/f+Fjf
yg0+fvMKbbcqjiXlrmp2sgxqvRwu9WhpoYI7/sqnhw9iqLdpchmZ8ILo+layt1ckm6exv9cIYrck
c3j9z3mWyjzkHxEWqFJjvCWHc2Mw2FrPlzL3n9DU9+ayC3G8XI/D8x8fDpTquagCdlHJkIp80g6G
EV/YIK8UaYsyHortkX4R/0uVNPJjM78lUQr7PQpdkkERTpS8O6yypZo4Zxfy6hV4X4Uc9euaE5qx
RvOTA3sGNWf5Y4QGgnl/K85JTsbUZ92/tjtb3X7+kWGaaT25758FcFnAsWAvsua00r6IP+ud2VJu
IzM1xbDYEQXK0UJP27aE95H4Y2zUFCI671ojg8yQmqVYI0Iy72LBvnbV6pYXtEG2J9x9GKTpz0M6
WJF5f9UPkSXBwjL6snRte37CznXRpMXiWSnecevCpK9M58S5ljJAVn+SPXqCBn0SVqUsMRTafwKB
eKxYboLjNSAlZ4Nh8KPbY8pcY+jw0LEovTf59YfTDowMtZZuT8FOLFULMutlWyHiR4Prc4rdO3AJ
c5s0Xz7tGbRBUd6P+9D4t/vqlPJl4Ox2emzzmHNP6TZgKzBlqd1oHbtryAciWN76aD3m9BX6cd3F
ezO5ljy/e6gA4FFPd9xSFReWeCUq2Tq86BglpkP8CldSoiD11sa9mFsT0MR2Az2NuYrpiGkRQ+vZ
KNbt/f4S65nDFcgHuKFWzA/+3nGM2e8hO9VNpA0tH0NiNB8m4sjg8YqKP5koS6E53grDQzoL4dvN
sTozZ26XAaONNANjW0+o7Afs8D9a8odFEYgw9z42zSvRn8sN3DCmKYTJaW/UFPiIf/eejSd8aDaj
WhhtRu1ocWTtdM75Ca/ylYDf1CW0CsOd6IdkGJPwUnG7Fn+NIlgeVr848ac6Jxl4aXUL0V2uiOid
qyY8IVMFm+OoBnJ2P3Ti2uIlvfgR9nI/6A82bUycG6zALZc1CtWmDVNWRqwgGxXI2PxRqghigX1/
cG9O2j8h4WZDXs2s4b5dL3JobQ4DfNwJOsBMZMIij6ebBxjoZTl4ndqqnEBUiTSqbovG1nUBU20t
AXoqU761VlBD8Kj6aLqUrJjWP4CSs+fjcBbt8oboZOVQoV6mZUwECJp1b7EB77eaQBPp8p53GzHi
ylDL+MgpwH86kvdhbqGS/ZU/VKrvrbJsS0vHfpSfV0gLgh/qB8vVrE2q79dHOg4A1vqDBkZiBUma
fCPjZ7IP7E69U7T6fhkJy9+z2JZ56i9frOKdvFEvrtVbpoFjsVZhqrQ2olVlqZJzB0F1qnoyeuc4
3+iOdPgmwRvU06p5mIsQ5H69WNrurRMcbJIv1YUENSfF48PnkcQhig/kkabN84O6w6OfUw4pBl2k
x5QBPSjzM+Lg7feA99tQYkkut4OQRp1fqHd3FzwANR869BUfnDNnL2y9mpVofsZo+qo1z465kSuj
GV8NukBSuwTgW3mC/Z7NvciKsmwyywPvhb17f/aLsS12o5YjEhZ3h5ACgSijc3ebhXpakZKck/un
caE3pLj1CVES0LrFPxqEjLU7R27tgSsFRhc4KJR+sLvH6IZL2eaRx/z31Z79qZvvpd5elmdGX8en
eH43nh1OB3e28+StPNxPy6Vhma0gqbct4UTAC6rrx2MaT49i4aOO0efgTIRMxyPvFVLcvHWI8oOw
m09ZbPonicHMspdE/Xpy3H7See6YfBtT8uide4XGXH3ord+I5sMog707I+h+MmVNlDOa9CFIJ53n
Xqo9ipj88/jiiwWvYF0i3A8qX9OJAG43Pzmfx+0fhKaR5darz5rV7WxqB6eL2KBROqOv6bIIPLs5
WsxcN3/S44ZixgsgVstL+NtcLKuJtzBa0uDHmbnpngZKJ8iyOUZEuByZgBMW0RBOqHza65j7kfkl
JL9ARP18mFDcRSwrh6UbuFIU4tOXl0Was51vvNgPJ2/meQ1a0A4qKFLMxc1A2vg9LvBOXwa1cDWK
h9mkWRD5yaCsDHYmIIUcwB4gyZzxUun5twM704lS+5fxgZm020ggdBzR7YEce1ewAEt12Al79yR5
5JTLZZzqvkkI+7C7RktBdKpehb7PYDeiIg/2YIhbjgrb2B1HieUBRAWQBcwsY/cmgR+77aitjlU3
O2r+Q3X8EtzaXcaualwVhvOEAuZnpaHG6x4ogWx72mRFAO06RxXlbhfoIi/lbmFp/y/evKSLkMIO
pHlTReORgu8yYhPpMRbYyN5t+lsjD3MDIqNlf6sK8FJK5JvbWxH5YwchoMjKGj0nVdHiHBWjGKqy
7edBt15bd6aZMUESkGyyOGRlzSJoA9lYEivmkPwNy5rk5qUngoOa6hjQ9g49LUAKSSyrvUlI7kEp
ONLzinJ797/yQtezOhTmFFgDziA7kEFtacAVyRrx7lRDIYCagmlFaDyT6jKoqAsCweOqkpcrfQHK
ZPEHf2+c1eHKs/azIzbOt1Cev+g27IU6h3tjBHTWk295SG0H8cgJAwSDilr/CmMVz8Lv/MUWO7zL
gdYGrJ8jjjJmdG1iWCqCpKIwvpdsuipDNBtFk13Qn24Urh0bXWkpb2GtlLQNIpdvzH/Y0eoypgHx
FoRIVV+VHHK4s4EW0kMs3q6yFZ9uiRPclpDd672mXP5+GdSugKQFUxHmzbssy4umIn3ZULG1hNNZ
n9H1a9rLXhPFK887KFfrfeBgHlbJaI16gr779QqesUr0FKRaW9tbx6SNcRFetNcuRtkXAdY2y+2Y
8sHnPN13FwJoSAtqQ0VT4C/BukvS9Ya306Qmx3RpNBYv+ad7CqIuF4nLnHckYC5zUyeiHlc4HcdZ
ddA9RdaMWMSKqHunMx1is6Giz8tteeA9C439WqT7+OOdd9oOdXf0OCCdULBftzqeCfzVXvofBhYl
ppfAF7DvL16+/EcTeLzYB+QQgRFPQIOyQUK6OsU1p6hHShrJM3t8k0CXLpy+/ln9mmAtQ6sXklZ3
DoQci9F3f44cfmIAKOB4Bsd4TgC8V9FWTCp6DSykQLdk5CNDt/lHVGWsnUOwwq3gXeeq9v9sHVAk
5O0XHU9ijIVoHoySynfEJawgTXSNXon+2YDAZsO+a3cajNe7gLTknYANOQOtRg1iT81CJRuysWhP
/OGtf7SF8piXMVeBuCJbYnt5Fbj/O8h2HDkmqrl5CBaswYm00hurDvKo5AaVob4ioVKmWHbB6WKJ
3HoZduKsUQXkSbLZAkPknepwIgoGA+cK5346mBUzlQJ8nf4Ja/QRiP371AlbuHnycU4ztxq+tSXF
n1xnKWMA9nKyHe0iRyzJ1F+wIMUl7coSIFrWAARRugYlIifmbpTZEfJA7syXJQYJsDRZXZQrE7HA
/rHHjrVw3PqNtqcHhVc4XJCI1eygWdioTM8KR4PkdPOPxFkI1az8sGc3o32LfmTqtAMg8GHzwsrL
odOeg15pf4QmNOfXfgRq+G7Hqiyzbz5i7aRlXynQrAA73ZVLn0+gcETnPR7y1KtLRBARAlZlaO3z
CYZrlxzSxY9pvlVvQUE4FDbQOx8/wElGquCeGfsyaeLiv0bJthP+vptlfKspC5lX2dEfbtfBvJEE
/rhXnSypgWV+YpqghBgq9hRW0DWUN3QZ9fJRcuyS58pqVJzxJ++PsgQv4zUZTXPyNNYt0Mfc4VAm
nvBUlo0mJFd/joZIdP5XQSiEznli54dHf+0Gu+Nv3Wx18OFTPJuRKK1B4znv8y9z2vTei9HNitD0
W/Z+g76RKgQbGpqvvw/Ml4pJE73bdS7BulNuEVXPilwe7FCV8N8DSW8LrhzJ1FhY8DVa4z38RwIN
JjPmFarZwUGA+Ehw/om+k+aEamNB0/dpptXFtG8OnYmfITAnnDSv6gvokrKimDHDvkMXw01SUWZf
ry42HcmqByFgYCvKSWffH+7+Mryx0Y6zElUdo5mz9Cnk1IeymFlJegX/XzkmAppqkseACFWTqPVu
zrXRVtAHuzjrOu+15RyfkFDwm5Q+4AL7HohPPTOaTxDF7saJvOSpY6j0YRNJws1lfmfY3Z+1vUQU
Lv5C7lHvFRgIJRHLRPQBhI9cXeR7szR0SLzsycnwLr/YVGrhMhLk43nws8/HWDN1J6L5hoXJMhZr
u1EwQsOnJXJpLEBefKxz6i0yyKVr86cmjBW/bqiH7vkC45lWVg13L5JkBKU748rQe1wWl5ykV9JP
1roCzzpLSLOPrFwEVFAplsX+ZqfAxBOaWDFZnCVVyHtrq1chUDmETkeHb1oigEwxMDUrgOc2ZUl2
n0ehrKUjQ5NsCua2cEDFXCBz6oyJgijxEwao6HSS3B1wFs9MTS4PkrqLHKR2VeP+NIuVOx4v5g5o
wFSY3/i2GEJgbyA+mJUw/cC5tiOkJ/HjndVkgasIso8AOYzDVBk6ngALPY58sG9V0GB1vNWMKbN9
rdOZz9+BICJ8esXwtLFeoNSD/Ma81U/JdPtDWkeRdulSP5N8Y6dNJ6nLipxZzuImNKUtw78WPZjd
gNzCcTTjSgZ1oDuGtG7CDZ4KN/Tb/9JjANi1EYBOXP7sxykDoN881/D+p9osYffIw0hoy5KlIuXw
XbkOs1Ukf7jtWXP2AWc6er/rRIZWSB/53hjw1Qd1wzEPKCD/VqULwP4TpF+77z+xsN4xzyp1MTSE
xHmwij94gAbA5aAmYds6vW7hcep7ErnbzdQVgFhsfzjYtz4SPvGpX/Y1g5loN6zbu64D0gGnSlmQ
QPe8PUQUz4Zkfxk8KiHWGa1FMI2/T/ZdhyEWkir3zGSxWvganmDokS6jPVbBxcfKWahqLqbiE+Bj
MNqQhzMdj7yzABuQdfzYHtpyXY1zQfnm9N/IAq2oukqjqYJOorzTSY73DBleDhzoSpq1jslT9vy3
pCQma+qUqInQZPNsnJKO2psCBgHe8rrbQGHA3dXn5MzdOduYEvcJqk9NbWZ1NIS1lU1P5HOLDgMj
C7Eg1T0KGuNxnQVp7c59pD2iEY4+vU82OqKIozRQEP+49wP5c6P8BJ9tTJ2by+jwDWzYJKfBcL1F
o8Fj3Yq6+J1ldVZOCJ1zyJdJ8Vz29wZjK2K08tXY+0lbynOQhLAqtlNGznGWhqmk4IGcl8LeiIKo
sH+Xfg0FndtejmR9HW2FOevQ8aXOgD7Wewz+SfccdKb6eTF90gRCWkK7rek1GcIJksOZKnL224bh
S6Yltw022KpF724XIgEUnwG5ad8nDCFiltsMMxFn3ryNZSp7b4GA2MdgWc7gvXOC4BWqAKU7/K2X
MA82wp1O/H753E8UppRM7mDqV85WZpgnn1n2v9PQFRgbInuYyGY/1msR10vmyQAzOeNtfAH7H6tZ
cTmVKV2gODe9t4mxSDNMceYtPuyCTVHJ0kArYfg633THAt3HaitWbEcPkhFhBx4FwseEdbnF+hnT
lT7PStzZgJtgV7+9B+1gz9buCLFc+OhtmRry76MfS4oAh1A78C5OKZELMdVIUym3OJDWBdc7L4ww
BPK4zyVwQK0yYjUCHDJ8aC6EDciN+l/wFtSrRz72Mf0IraJP6xzOaDI/LAXpfrGFnFnCiNe8H8y0
4Rzu6i5YfeStShhDEmUQ4kxdf2gVbBB8MOkWqoLMC23S4KRGV9BtEADZIL1QQtxwiJ32HL1ZpVqm
fp2ocFazmMt+pTnH6vGdRWhW8v/y14xQWKvZYP3QQJiHrEz1hbmFxbTW/8L+MGJyycd44AszWGQ4
benXubxDhzIXRuwo+8Zgwha7f3joLyLZYuHw40cSDHs/uVZXdNZFxHzJ/zlWqMga3Sj923cz4o6h
xIKQdQQE4SVFzntkGHs7Dhd/w0FLMBmOIt/0b2peT9YnRqGXOn1VHq9CgQLCyt4bLsq9HRarOTI4
SdxTj3TTaawTDzjnLnC3j6E1SKJZkCJotOtbw4KnfPztgn8EidFLdQqFOSIPKIpxBPwDMr2pVdnQ
Ts2tJAEtmxeFlZogXMdC8woHXWNhgC9ceQDIK3Etu1ao8dHOc35KCFlR1Xnoxvr25LcGZOWOxIOl
EmGMS/AP9DGc1iH53iuDN0TDT0KpezV0ytVBbCnQOR57X4n8plnn7FbL/Bv8uglR7aFzQTCWQifa
eXlVVg45b6O6K+H1IJjeuq+LPOuDLaEbQW/Z8+fM2gRxfSDjhmeL3FLPemxH01iZpKe21wIR/YCT
QgWzh5FyuXFsIFKdQKGwhko+wLM16jQTqVdYKmhMUS63P6VT/PEbagh2HGPj+G2QO1ajSb/+9NBn
wyR7IeJ9dpMBAscNbJaZvN9K3d0oLYHJcPT5f3sx1tWsw94q6/OMl9wuKTtAAAvoYBLtUxOd9IMt
2VWQbQa59ASnTFqYcVOUJBTSDzo1Rh84mNKGtcKg+XUq30FMCIlyizMNLZgosEBcXdMynQmiaN0s
OxaMwd68iDux5JvxpNATAl2YZyzCxQwQh72Hh7db/ucfHSKe/jL0oOt+hFMNmzx+EzhVjHNoAqHl
SoMQbDpUe/Wogj2vqUwrSlmnestrIifB2eyCXTcAxu5U/3T3j8Q2UQL5dDlQdVKAOuoVVHtd5FRQ
csRjdFhjQoPkJG/gbRHIes/KMrE+h8tSIlZhtX2D8g7SAXL/hn/HVI9mvd/Gh9F+uVEDXUy7q/sg
VIYZhT5Czd3M0wPcVoxvew13xMbVXyDdLziN6aAvASIKKCvSi7qgS479aSzz22kEU/s3xhuNoBn+
0o+9isGqVqv5UlverJ2SLED4F/wla/iu9z1/ieUQQ2bXhSjm26Uww8L+wjn2B9CyFWsjibBMPnrG
nQDI86JmhhMVKkD069Oo0zQZ907ClDaw39BtJiiyH7EQ8DZJbT/x33hXPGyex6LvsZQCXOVykMjA
71mCm7HsALd/3/D9bzmCcH9+rhH8Pwoa2fpS6ftxhL3UBjdzugjzzKDu9azbXIKF2ADu7RFyxZM6
VAXLAGGnebzMDSHpL0qIuZanJHdNZptl7OowkxIDO/GG+V9iB9MaYQ72Ok6TOQYmp2eYTQGHz5qZ
NT48AxZKNRpc4bdd7K4pGRM9WHuMbkbU/5ViFeXqpvuJG3GyhmTBY428pkDRZzXo5fGHoh1pyPmj
nAb1MCQKran6hMGA69JDdQQKH2thlYauA7kEXzqOvYwqmJokvLevGsBx61c2hJ+RQVVWlhTQUTH1
PnWU9fwhmUyy+VXTxEOkFX04hiNz/wZUlpg94ldF1DYc+BlTYxVAjlv//XQ8raNrPP+NS/0DNXzr
WewgKDBMPY/w3VNIBE7k01a9zEDZwxLkzUJCS3At9PBIO99of334v68nTTTpvDR2fHD5ygSfzh2Z
bCfxj3EPndL2KuovOT0qzE7pacdEQ9BjDzY7afKugFDTKM2Uy7PPN6TT4igu1ixTAQKnwH0hDvY6
13sold1FYX9iP6U9Y+m/kUN1v2w1gXSDksEzdJWOJb+e4Jm5VwnVHam1Ax4fM9dea6cVjKGL1b0v
deG7ol6QtXJfZzEIWNbfXiUFjqv/fo+cqOHXK8S33ADSm0veg1cPb4KAX9KA6gYjRH8713+FNk/W
ipdwYx3CMUiDaTBSXJE0+wuV6PXPeznynIYnlAFV2CeSGvejIfjpDoJK6ZAVFnqK9zkISOWXkGUY
/ZEVjIszj1KOv+QJb2wF9E1265PBxJCwySEZfk1ucz1prnuQxNC+BPbbtVSyfwR+1POfWWz3U2El
ngFQIuaeOpoT98qgYjDDXcUjKUFlKq+C81kOkUPzN6BPgZGOKQtaw5TU7VyoTGPnoexVub9yw81r
zKCQliHluX+jZ+G4O5TlTv0DazeXQhHdYkI2UVDWheR3jY9d26kUqcpieFsgOL8H1DvxXHlomNP8
p7+OZpcS6oeQ/KeLzK5krpXyqT/7z+ol/uAyjGkhmA7GVK9J4ovxMlRojeorph2LZzDK3ahSPQ3v
GPaAnDOU33uJHUDwS65o4ovqMtG5xmyRuewh4pME7IpYaD/5Rio6UvXDypwIk8unaklmZivgdyDX
AJZnblpwPmc7KipfK0Vk8ncLBQP+G4tosxkN4Te8LvtE+JTy2gq6DobMHYrjFCFwY0PJ4IqW1p//
73TcKYUW8feZAmZO4TG//nHK1Zx/O0N6JO/RKW4Zv0LqzTRqW+sUC2Ux98PszfG7RjVRMRGPY0fA
jNyxsZqx8KNz8f+ujpjz45016+S1kNzjvZfVMbUmASDHjNgzWzZ0iyLkiEjEWgeqyWgrhX7bGZOE
EGnEhCBNeyQUlO2r3aEtyhv6rXCXR4Ctdiz0ZSvPBN4huuuLTPnr7Immpt/S9HdAoM671pEOkkn2
y+IgNS4jTD7eWw7saJynKYKY71dK3sRmH4K/Mq5Gw49WSJLJ0b7zZq3i+ZNv+NeHrHJVePFCA17Z
JAIaReUeDB1sRnVBOOKIkRKsTaHjtX8FJfQ+sCBgCvX2ehKsAWY2qVupNVSOpMR3t50+Iv7ru4gR
3GOMI1aICqg+O12fQFBmDMRjOLT1qeQURKEJBt2QW+tlzh4+L11tQ+9mqdQBwku5l1x/8H1BOdVl
zU0Xh2nPO0S3Qdpkpk7wQG1CSsrE7h4KCRtE2mys1LR2gyVdeTDuhi0GpmHh6XIU2k8iv6GYNdBO
+/bEUsUJEm3721g/zGjlMOB13bR9+KdmjJYwx/fscuIAXI0ejjxXpUMwPT5WxvDaMP5OTXKUYS4Z
s9gCORo37SLskhpNPP9bvSH1ZblPBeDmLUFRIzOBVR9SJqanpsPgGKBodG6Ea3b/aZiaPVbbXUDR
2uUDJSW7O9MPpjAfR+reWOOZbJ/8Y3zZIp0zWGWfymxWq1Uvo0ZdhYc7hiVNW/kUBnDvghdtYgz6
O8fN9HjWTSTsTLYTXNcrB9sC8Q/r2gITkfA5l/1O7wTs6SVu+X5jTVT7bHu9rtdcTTrS/nz0qJP2
/cNMbyNNRjFEYBaJLLsrusz1EHX34BpKKnezCWDrzUxwgNaaOgDNZMg5UmPHFW2TxRB5dl9CQlSC
Ndiu4rJG8t+ycYPhW84G+pBOeRpECpbiA7FeMwcweaUkxuEYy6QjHogCzn07PKO2E92XCpuVigAs
bCV83KKuoJUUb7+iAzYlMtdNu0ExgxJ7lfcTITYRaL+YOOTau6z9PHXT4pm8I9d0vxcyGjQD/LpM
x5Lxva1demoprqbPn81aQD0lbR2S/6eF07uorZuki5GJpip+wmx3uNhtQZAB+iLLFWJ7rJ58uxLe
5+C+jcwlZlbF2tVHzhCaiWPZTuGikezE1TFt4Ph2yCSEVxFDQRDCV5xegVe6GcaQcLMXzYGwmVGG
Zh3NSBPPe+ztbv8QZWoL1wXVzhb0GBQqaPzVGcIBLHWKhstKSKfRmFAxlC/sZ1Vy/ato7CPfj0xc
WVzScKsefr+3HHwKuuMS7MdFnnDlv/VT3erY1bLoXPpEU6Rk46svyjxLkajBYkjkSRCx6Pu7AO9d
1PPdzf5WjdXZwxAtl5rzeHOGTL5QcPFFGQYQhT5KWhz9KW/6TZsa5ZjOUtR5kyGxrdwSb1YFLdJq
Luw1Eu2XW3KeNumrLzxUYMzq9mNoB7aJpCHFNZlg96gNL+WHoPcZAkM3ITpmcnFuKg+Y/2W1vW8n
bCF+Jk0QKHC3UYfyqe8ptRFwHubZN2dzK3dRhBX8uN7L8z9elpuwa3mXDymQuh/+YHf950fruUDQ
WOysW98i1vn8tiL+6HgnIT50dZTjnaE0IeOBn921BE7fQWmBSfF1zZHEDfQDv47qbFQb130HOZe0
RDx0VTGFZLm8LCGHmbPc8/6qzXp80Na2SugxA8C+wz5rtf0D4Qj91k6asrNGk4F1MNCiJTEaRV50
cvEKWyAviIPoczU38PQSKe9zrrqrtnvqULOhubv/ba0rlR7exLUj5pq4sHA0nlf1wH04NtjNBlCj
4v4VRVy9GlmKCisg3mzoF+jiSos/ioFp7jd901nXBfF5Q20lX+0GDeZCLWRyWG5Utznshw6k69XU
7IzH3tlNf1WYFc9fcd8Zr4cAG2gxTVBO9mfGJzlUE6C1QKSoaoLcV7EQAh2BJg2AH5jsLgXA5grd
i2xzLmfMmwB4ZmuFHsPbksB9KoWmpLtfPj8MCfrO6x87kFZnjPJzCILcZoJD4OU2lA3rJd5cp+VA
7Icpe2DjAywcWmYONUOar8LYojvLAp847wa2a3QRzehcvMdu+ERc9trRaUFBmfeqTruCmsa82Rt2
lPwV8K71HF9ih9TBPpHH5aMtu31Eo+J3mVh3Wm4u3SsH0DbrEBI4Saco4uKHqzlGB+g5cHvW42/u
OPdV7DpuBLThXfpzGTG13AZY+Ezy/vH1kk22wdADHxDV4GqDDrmo85+R96t325VNmNo/B65hxzHg
+13KG4Q+dQ3hRDAQHWFVHQPrP312ZANQWLc0z6aWMLIV+r177N+GxyQA+HUTJJZFdFyPOBlj9EE/
UwUcWJz1zdaJSUXezelB+xDdFeZW+usxTCZv+rw397xp9E5O7E8n8FoH8+Dt/KtSZUULgqzA02X/
fdXPMU/34/CWpTFmII5QfQmrxtGEdkezijTKCv1n+a5h46epJRgzKcVhjkpKd4Sh/2bLh8NvJqK0
kyBRWFQ0ajxPOXHOmXpUiE5sGGmG79Cq/hCSKs40ne6zn32u/LiPmTB8YIQxEYWXx/YsQmlrfvNv
hKw2HxgWa3Ec4CqIMhM1NW+ryTcaK8mTlrhM9iSYXt1xb0ALFRD1iz6SiuYscqrKKC7l7kchOBrg
aqdu9L9r20rwIwFKfeeQqfsiSv04/flLQNHb/5eW8G54FTxdFURK5X805/YCy3UzvSUgKR4IwD/i
6FajqGPIraqIUcpUj8A+7pwUjIL2m4lPqAjFH1TtRtDqzkudQiK/6CDSrPPJ87m6/+qTj3BLPh0+
sC/bJVC2mLRccrXLQoiMCDgC/6pDByGw9Y7YYFFgeYgGAyy4Q0V8/oFcg4kL94lD9VfUDRsN2HaX
SPT52VUL/RC7+zXx9Ee9I3qw4V/w4afxVnV07SYaaToWaRTBj/UknG/W9FqVuVnlsJjc7PwQmU4I
ZFK6Sfj5HlbtRUoMYI5gwfxTLNluh4CrOjJfMTYlxK8iF4P5d6TAutJrGBkIOWE3xT3GV/R8IJqV
bxnQEfI0YVJ1lWVjyPy7T4XjOAG/RKF9fO8lFgqqbHFYl9RfHUgLzqrg2KsxLJsrwTDiQvE6UQMZ
Ws2Hmspe5xvSYHLqF4jwvkQDJ6ZotSjiIm9OW8Vsmu9X0AGYmTUAdrJSzLoLpMeUA7tI/m2px8HH
DksQiMUdZ4IyJi8u9FV47zkJkFKTK2Zq5HfcpkzdzD32W9WsbwWpwlnQyMGXnihck+Y2AKRuh9Ks
pCDEjy9z4XM3ggguenK/hmZOBSlnpgwQtbKLZOb0hihPXttHB6/wyBur2mpJjnUaG+CL7IycSSte
iWE8V7NvwM17r4ZLGoeD6dc6qeqfCvBR03PovkZ+evo3Vk4XVv6Sl/W8D3wwjviWZQ/NbliPwp/H
2gcLNg99Lzd/5yDfzJPlYWH+cxm8wyMM47ROQl1mG3Uwvpqssi31bJGYQX0o8XIRJ6c6i9TXlWZi
wwlgfKSitViDzDc+IGbkYuqnqTf03D6YRH6sHZ51Fm54ab1xQEBHM6icm57Zk1HaXjFhenQC0I2i
tGy06f713hVbPkaWI5YnVr16HWp9xrsDnnCtnYHeSwlu/0kIFiBunL55R+Z6S6baZse09/OQs7w4
LdKVa4QFZAU2JhNxydJcAqQL1xmDjpZddGyViWOvPx5HHAwOvNE4R5+EUZBHLTFc12tIDuqNOMRY
2IF/WE+Nnx8gHvrFx+rTxDP5LuUW2Jq07++P/YniPNK/fVNgOvAgPobPZ6Dgg+LenjBEOHdg7LsS
3XNX6sKKyRGl3ZmOZzcT5F+/Gnaj5RDrIX1aQpAunwMn58IftBcH2QMiMALHfZNiqiiL8S5QFGEo
GsfX/opPC4H9uMKAd23Awbt7cCnfkNxS2C1l82OuI6DEBfNLH+YfJGoq4IY2ncAvPpNNT3y9VuVa
s3wzHg66HNgmQzZZ41+psZLUGMKdTHtn94ro3XYJgg2GQ9ngiYr2w2erFMvH/LxTP6RiC5YM0LCr
yE4wKS+Vognaqpt1cH4msVbTv33Glns6McwB48yX8AWa+GTo14fROh0YhXGCkXA5O0OCvaAGrVkO
bq5Bn6Hh0JaIqA2VbOhluLnqcpn4JaSPK1AKMCUbx9IQs7qVRLa827OQGURQJqJ4kaS7dtRIkcCZ
6FszoAm+kuYxeWyqRQeyWVyvNzOr7QvzNK1rf4P4IkauVBYchlWUNTZ4r+QD3gr3b/jbeJdA9j4o
jETSJZ5BYrvEV7sfJxGZeQ5chGsZdP2sUewHB/DFepPEVV46HR34+n/q6oXoj9JZsThGJnJ1emOr
kdX3Sbuyb5i+f86/qTc53QG+cjp7WWcfxJGIgv72AGf1GzpxebfB3l0+k+cNeD1ODOWpz14lX7sT
6o3zjNC/DPtA87d5FCDrdFra4qcBHLJgObCzyRUyIMUXqiVdNvB/HD1euQwgocxLcSDjvGvB87cc
vjqATe0jjFLTrXevswGFPECBjeiChp9BAH1oHLqy/9fcLTRyTkkg+BEK4BkoWmj9LpnnRhdgl8Ly
UNq4R4Y2nlVpo8D3p9LZNypTrddbyNJ4DINlCD8RIg6PTXwGKXswYNSFYl3KdalJJPzecxQjiYL7
aZa4AP6aGN/03vscRndDNwJWk15QXGsVVBgpDzsuCjMJg33Pp8OoSufrRxUkCyr438AXw665O7UL
QxF3Ww0hhmJpVaQc7uHexUdMa1LTzTE/yXzvTGtVusqFs4pT8hs2FY2Js6DHiOttrD88f/5Pb/7W
COB0tWAwKt/q2MiX2jlJprBn15MiH/f7CjxKnYfr3tVtCY1OP6shm6L4GXaku9o0cEa2O8uQbWi5
IycKNj7wTdMevo/lf6Y+FPgrEXvb3KQtDEwwtYabYcsMXA5/CvDxftDNIzzZc2EqzmU/gzT+i9Jw
jL6Wy5Mk//AkHsXenpV8SiXkqIz61yo3BPAvhp4LQZB4bY5QOa2Zm73cDX8eFEc9OjWegXPQ+rre
bkkuH5Tn64kxB1ZPwrJqwWXPQ7f3YMyMk/+YcEOI9nP3uX7WXEJW/wRgna8jJ7p9QHQnEYuFqD4d
10j3IXl1ksVVunf124CAUb0I5TkEkeVb4PZSS3xWDa1Ldl08awIQ4/8aOOKOrkdJoWXV3hQpHDIj
Awb+/dMGa4tiZzUCDbnLoEeCLA6/RktJ6j+ThdARqTzJi6VHLJMU+b/dQg5Q7ZR4M+s3eUwZ+nPp
JSEqN1C0OYLttQFJWfFTkqhXKQz2xDlygMS/zLevFDCNa6M0eP3agYnHnbAS/X+NAdlxmacaJTt7
wBTw3Q8TgYYtcjx9vt5SHdsGNP5BcAK6cOf6e4qMOOvSCykKMdrUeMns9INFLsX04xfduBdOvv7/
qnBslFOIG0n2u0Et+kPrT5Dl4T4Y5rbnz2J1fspQ8/s2YSYLvR4MTRyS1uoUsG9VdOaPA3W7LEfp
lXcFKxSxpWrwkOnS+MP5G6nWBHN/RJliycN6mTIkJ9IeG2re4GUrvEbr96jg/S+ZO9/9UZLlpJiW
1d9Fk65dqUreXZY6FX0YQsPoRq5PCPqClBylwHRIeynPLLl/3b7SkEjKZN5WyvhvAv/tAos1WWW1
+BIPmWLwNtQ0bGvIWoOF4fQQJrRGJdythLEq8WPsbbkwHP5xIeZSYy9XG2NzlTsIzYdH/JZNbEjs
CP3LdzzcRcmT2qcOpMII+rnQa/yuz8SSZhUMScIvBWHJ9OPT/+DuOBUDpsIRYSHSyc8VsepVArBn
6KIpXK90fzl+KqbgHBqdTZy8S5kcfEfJ3RMrd5sqBL5h+jvXsQG2wJ+tWe7Cm3hlcq4xsFrmvTmK
rzwaRho5dGNFmRuoyGSPVGWXgQbQERvLcvm+evQbDMbbJQLoDcuopSIlffdoB5A9xb7sNXg6xAn6
Auvyj9/OmZaexhXSV3bYkWnL9EsHomd+BwhyMVl5pC9gM+sw2U4Y4AlRwzyryLv/FXFB8PiHJ+2O
r1umBVb+6Ft3Qm9nDYHujfXeZeO1iwUUX1PmFiKW2K/fnkb/X9A+6Ofbl/CR6IYIEPU3p3lC+0z+
2xjYNXft4pthLas+8IUICQwI/y9RoIHRDiNmWxQ55r5/hK5h0ykv/C6kSeO24xccUcMMDKnLxHsy
cLaK65M8NPyS9AiSWfgdYqfg40RxXz32UoZQ8RpJecR4Pk8WhxwCFLFKNco3pglIpRf/2bXs4/F5
9RQIuZEfHBTz+u1b/LrPSbtM9Vh0tQX0oeeXUbAn/mfQrzETGglxFo/0fn//RGAZ8vQFDjHPbz8J
/rB94b/Vbf1Sf3PJu3lnyl8ZuZPllrIKDzmfwOeBEpoZ9Kbudw+1CcZMQi+hrq6mhyt12ZCrv1Rf
PuVsoIUQ6Nem7A385H5MieQrPlLmjqi0K8YyOZwh63nPZPEO4rf0dDQnDMdwzexJiHqgW+8g1pdS
8T7IV0VxTCFe5XonluM8yCicUpePjrd4g+FD72eil7ir+t1rSdqJynjj7i1vUA3WdTDp8XDvsQvN
ZwTm66jU2P3nGO3Xs12Euji4InBPvRq01ttd0cd6wshgFHQa8ot92iE95zKC/lfwSQiqjV3NZsvf
9Tg9EwPAjcJSEHnwE3bqjpdP+UxK3hWnU6OC87CeEUR8r8sty8/7vcfCugANXinw/zRa+h+si9Gv
EMSQIJ1cOxwbHWCKvgkjalAcJAeg+q0G/Hf+z1U7zR/NPMBs1vIYxMGWFSeCA/EQ2kh7jzpBI3js
VFHzCZBWTAiy4zcCYris4nW24RhYgXXRNkfWNLmmDPtNDbQMLnaT5JvieAH0rufFaVkiMkCQF6l8
BOsFuVkvFLji+w59n9HB3pCjxBZNE4tKqDI6Gp9fX65CZCpqja9uZsz4SvYnIPkdtbdwmgpvk8t+
cOxe/RzDZJ4fJD6KslrVNo5sj1Lh7WuSkjI+ppB8Pfxm7hpB53wSE6ltBqMAm25AACVAM8+8Lg/3
hpSAIlTQy7UMLFeW6tQDFkGfqwLPYbGc5YpOVwHORoiC65B6vIcvhRgcFsT6RFaYvylwyEeKXP8O
fa9HItgDS/ehTHB9naZpM4kWC3ij0mT1z99D04QXmldsZ8RBQa5Ktt0xFqaYZIhUsbmEBufwIA0G
RdIv9T3VCwAGMhwE8yapAlzN+jI2ZJkD2BSj9b+7mqRsI+B99Qk9RB7Jmiyf8cawHieBeIU3cFkQ
hCg/1XS2eYMI8VSJCRWI0atwiG8bIkZq4PoZh7gcC+7cXQHRfgIrqyJxXsXCaloVX5cxZoa1Wy8C
Ptu4IaLZyO9KNCFR/HxB36qsuCZLc3repi7MLr94wztaJU2rdf9SbsuWw+4ORcmNyVIln06M1bkv
17w6SwO4Bc3DSeSnpIsABAtbnzSN6NVy1WhKs2Z6gbsa5a6pUe2MeLLWD64K0eFGa4DOpqTftahe
ekXKECXwJVLC1z4FlKtrW7GIbKts+/01WH3gztX6ibBSRzMT8exqQ9hwoEDpsHpD1c0gnryNBK7l
8DNBMTxHoaHcZvv3IC7xiDMmneLoUgvqW35lY8yx5pUMMxXZCHY4Uo7gSUJbMXMj0TLV99cevDnE
bPEvwLEvwgcasJNsEFSUkxw8G7i1dNahbqCMHZdHOFZQGqIDnyi3ar5mKX3/pv4F9NXnNKeMj7Yv
ylizkg9JRX7JzDyZ6bqdF+M20qYZ9wTURBNzf1Tpe649Vsvv1ocugLFO0ktU8jWjAb9H4kigutky
sjRwAoBeDhd1iIWeAbpY9Pu8ohsG2lyqaTL2FI4fvHAywpUcV5IEoj18nlpLMqYd7fH7vXGnuCHu
KC4ZoU26D9xIo3bukXAeotRViu75M3g1eu1gbPqAspbGB17H8+Kwu+0OipXajaTEK+XP3SI5Zotc
Ot1UiZ6ihkcldYrKomAhKR6JzbFQvBGUaezCLN1cBcKfIuVCZCCMy8ZbNuLMyBnEOktGlIgZ9xUN
Vj7weEnwtLxvIVqbwCFZqZpd3+q5LN+htM6RFvmNOng2GFHTJ2VUbxR89Z/VPsuUVOv6yr6MID15
uFC2bgYEbbNxGmCLjv0wQqazAuplQDyR8eRheh5ZDJVaYgqU+uEyqJ8LtKsNu4rLDlwQurorh/uW
49RFfAyW4Y7mQDTMipjwGVy47hpB4BU9IXi7bvqRuhNhcnTlAXvFiObjArZqGXpA4edacVTboA2x
3gOaEhMRRxH3++NkeM8sbJktxcFPj/vRPez7FfwmYdEZOEAkN50lKgCKZ+IC3jAgD1Lhl+mLgo/+
JNo8NkPDuJ6TuO++oDdG4nmTFsIxhS5VW5OdHhLuL6hcS/VSBD0hGczLXBMsvzqlx6yuGEh6dHNR
VkoCTqzSo/VvSnB/VdLiByvEDtLIo6eeTpc8BXtmAv1ctTEZFIKBN6SV1sl2mVDWdbMoZM0Auikm
x0xpWAeKN8LOF+lTRBbyevKlskixXE1t2gbpifSJfsmyxHq6NxGthbToyo6fZR5iL4rMOxyghgsB
mSsK6kUjQPAfth8TUowlLjLzapQkYhla9WJf8g8uU1jtnJM/DKju0btxN+VXXPktzUlNv/QuTjkD
H4+UNzkgKHUiYJFcugwItsTU2NTqe878NhaP+CHSnN83ruEOfLbqG5sLX3U8PjL9T26gCh1pcTiK
xj43/IOxLL4R1EwMpG3Psf2Q3qKdsV2lheKdlP/Pge4wNxYWhws9NibtKHoT1767Puajdc7KdT1q
6sBGGzUf7G8cQVHZD+6D/evILNjIImWZv+l+C+9GuxmztRfb74kP1+adKjAYmQaHalRwui8G/kLs
YThG9GdXhW8Kx3lmsdlfQ0mX/+2DLinpeYjbvL2Rso7aHBH4AvU2rYtegVSbXQtD2N37C1Bv6fdB
ZRl7XbiksPO2oKvexRX6YGCHjOP53icc/xvEgn6SHIQbQlPY2ePVAwrelrN/8GUtzLkElXzwJfIG
6nxrWhDRWlZdGmoOFMa0zpOB4zV30pvaPza8Vg5FmW9bY7KEBOG8FaVo/yULz/BPS4Pr7SmYCHue
yjL0BhMetRsvZrpFtSZSR1X9oLYKd+p/oRS2IMBbEn6uQm7kJEFsYNH9nmMvRJjPxmHUzcSDpaO5
IDaIqBKcjZ1jmm3iPnjxUgDLyV17ub8rfnQXzeTCZPXxdwWiS5FM6UlAOe7yCXzh9ste6DTHaGTM
sRGNWqgKgwbajQndRveh/xfdBndKaEkx+tmkkZxk8F4wGrxA1jMuD2iw+1xfAF7e//29zMFq4Su+
UDclNpSSK5nCrdrvbdyX2PEuGnWyQvoimGdR3aKXE4dmJUtJQxPJ8haVc8cVsLYZPZL/YU6ibEvE
pV1Co/S7Fy3QcnXte+ENc+kE+dP2Zk4zj++YThOglWzcOSdFhJSKSWfQuS058VP9MrpdNZNREHB7
ohH3N7Ri6mswrqlszc+040FPc2MDEC9Nzu3Sg+D3uUfHdF/PD/Z0PXrrnyioiAKH7RLOzeCxGOSE
n02lXxMdJtPq0RxQtqEtGkujVM8zAZmetw6JM6YzwJQLRl6ONhmBJrn+9OU9p9CfvkLtvDF8aYpN
p+FQtfxd9Na0D6ZpfS0VmKSq+UuPLw7/+zdNstWNMYGvqIWAJu/H4euNVh5pwW7OZ2kt4Q3bNYh7
mOOB/IMJh3LGrypPuZpGv1P16WRruQ+p15qzX6qQdprX00C4ra0QGELqVHvHPwrYx8Tu/ps6gRDv
q8VoOSLnclhakrxN5Gz1ExLUwe9sbxcvfa4VQaM35JX/kpBAkBj4sn0ApHNxJhM0KslIfgQtEcRc
T0W/qlWzX/dhr7kHECxEevzAXAIJg77uuhZUs/pBNqD+20CX63FPar9pz0yPhmyOm/egldJna3iq
ZkQg0Kv8iRmo0QzYNdXVMO5fGZ75ZgU5fWC2c+BzmdQxcLIqOv03PvItiROM0E8GWzGhhqbeZDL0
KxoWi2j4GpGzyfZiri2Tb0LiVav7gbyc8uvvjZuBnDc/mC256gocNE8Sf2M/M+beZCq6FJewbe8J
1v4n1nxHPE4yUo/JUO4vDv6bGLzSyeDa6Kj9njl8hjJ3lGLOQj1Aco7nQSYdW/17rJuGF2EJRZXX
ncROQOack7hxFifg8GlcrCE51Y9nTwCzrWbVHqtvvKW5TIH0i6hQtRG1+IDBGV2MdfrIM9ESQd7D
4Wv/PwtrLZrl9hotB0lD634TjfT5WUQX/9cwhWOMuyYRp2fToo8bVa68Ts3nALi+67IVIOL40XGd
MyNUOGHR0b543WD83g0eqrGpMjnaK35N+1Zug2K1lATzu4Wegm6rcA0vJAwP0oBOYa5Ng1DYMZF2
pkxgftBawUIXMCxDLpqOqBngwyi1rrQghcL35045w+n/JYbatum1FU44JFJebM4k3SIxtzV7z45H
lNTW7qBSnr5PyFRx0kKVulQZVKpqN9mmdOK5sCIvnsB+wlObXDGkFjaDh30Y8wWzCFgO3WFfey/N
obiUx7zHh20Ka1DALEur5WMdVMK7NMksqZZ0pl1lhsHvOgk8Q3vO0J8rjibRC5LsytGjWJx7k9Jq
TJfdlDJ4MF5tDXhlsj+gXzYiiGI7Jz9c+J3Sdihtauv42zJgNcEU+IU9mGbON9BIrGjtXatts5XX
mWHJTIuRVU6DW7qNOHh7/HVYfVLRf/0bFirZG5gcDiegwQVRLFXHygfzi5d8gtGKyEFY+Jq+uagW
8NAvUTy5dCLKlNTK/YUqbE9rauyBqBiF3Da9moR+QZweJ9UtctjNcGm+b8XHKIAZG5ByOtkB2Bnd
i4lAb7+L4pccTxDLOR6k7QlVHWcq/UIrJRe+7ItNgFr1QZlxQBaM+Tyoxf39uIO23QO/b3pcAe+n
edCcz3qdPS0JR0/OUhP2/9bfT20CKxnNVxdtjUVKO5SHPG49XX/RczODCiuErSGfvy/K7BIpH3QJ
kCdhoN1UelROyWOf+eFU+SszmZcSC3AFm1Q/82O525vGihtQJ8Bomx9FA474/mjndeCyjRJF1Dps
YTc1k92c+N6/+uNGRG7qvb4aPgsZgtAUdf6aC8Qmk0oq4xqkTwIcFcajHheHbTBv2bERRhiAJHd7
p4DeKQaxXqOWvuGj2u0Ika82Q0uUlSZW4CcrAYMZNe+a37b0vz5QMwPtI9CsYB/2HF1sqwldNU5E
EyEGmvYeQoHNCq2kRcY3BprKdTLobJ0zGt2yAHMq4YLrFTH+cAcoVEu/ez6grEGq1xc5j8KCc3AE
Xdtbl0kKqcA9iuVWcgB/xWuT8nH9b7FIu+xIxZ9WTS1oJMjQYj8IBiEfysxLAkYtRsKw7CInNcc9
vqpEQaWhoMpOe3RhhBkgUPxgrjDpThOqJ8Di9SmJyrKlixe7TxkPt3nMfz/Zu2VTB/u54iqg26kr
zW+0hnhDOf+hMAv4s2cjI30s4Zg7+md5AA7XZYcHDAf1VtE8njCo82AhoydN/uKSVqzejztvAopo
wisbnBHabuU6Tn90d3xSwQhZ3x7bw/5ja6OIh6en94EDWL75tGmHUW3U5RsUoTm9R5UiYx+gYaAl
UsjBJla2Fn5dqZ8D1NJWE2nuSp3Y+h0pOkj0VOvD5OsRjEF2lCXooA7eePcCvGlZv86UxPD5Bs07
CcVZEzkgoTc6IjuF1GYif7Bb+U7edJKhJ3eQ4pO0IXzAcOach8Ew9pT5StnQDq4NHQG8powd4SqW
oC80MMTAc2evCtvMCvnftMgmjAWKs/H5RJBTutNOW8D8ty0RQYH83xNOkZWI9rDh4aCfA2/V3sqH
37VEk5iy1vMj9kJzwBBm3Sw4UH6eFQB2xTGBd9fhztw9nweS0pXxIXaUOo0kIloTwW4LmYWRotf0
TE3aQyYDppDjfVf/GdPV+Qf9ocKBWb7IFbpldkl/u3/JG3gg2qcnFXa+5uH21wR157unYhEHQa4M
A2Watd0NMncmdZ0hx3LSdv+UgqgQmValMOruVOmYUL6WPWnUozg+erbU1UzemdrhB0H8iqqrqqro
/G+wIcd2oRAnZSYgffaEgN7l+pcJERpl8hvomyBGyAtaDYrHBhwM+P3hAZ47ST1zo0qOrLWAtQNY
fy0D3Aut6puJ2c02e0jGwh8a2m8x/80BET9Kg9vZQek4XsYZzS73sP4KhICElV6Z8n50ZSEMLwdf
F3fwD8J8eidmMdiktK3f6OH6VqHR6SP02daq6CtxmxblkQvdo0AUnl4qE52stu+9oqOd/W6gFPqD
kJ7vEl3hty3cCjGIP5WjdLOxAuph2Ihu2xR9LxO7ljJzon4KdvnIHkY0nxI/WOEZg8kLAnmXqOyk
l4OIqf00S6uKrJH5E8H1JbeeMood0kZlEVQHRGrREpwF0d14jE1YVJ1Wbxx0DP3CktR+Dw6Rnk2b
KRiFXqDJqoQppF86EHCurgyBICSIKGVUEyG1VvmRy00AUlX0WvJ1s5qUNF/nyZDgaApIu+Nqqtqk
hGOdzk00IWoCE0012cvHyN7Y1nQl4vvT7ICUnqL8NnQPkgOdTQdOmQILcQCzeKKeN0vhNAoOVnjw
2wGXXJgl7BAa1DyILUJMr3NuNvAiiUTmkKVI8tUZDdzsp19ZKf7ry36MeL+YsvirUgJk2x5OIZox
l6Ff5tyBQxL0MWS9INviqJzNu9mFkGztRIKIX1Y1CIl8I4Ali7YUMYI34rr/tt5/a6OVuuzVj/JV
/JZr/lZRVmWT7BeGKgDYeipxaNxaxKEXOnQ8FDc9KH4SrLSRTTMI2mDrZFxPQ6SLSHe/gho4PtAU
I/Yr3T3MtjazGBT+B0vGqSjKqxa1ZUb6NQ9Q+799oHfP1QvesSFBpeE0nNaWyjK5ADQsft+PC9q8
rVS92ayVoCnyYMxpWupRXIib39OCJ2rOVjoxESTxyLT3hYI8csQ+I5mG7WV8pI7vULb1khlui3d6
7JmrT1pzUweRX9IpwfdDmiCXAmaaA2E69zcaZgt+vCcKC70KDwFuSl2wCtPghSwKbYpYZgeIn0lM
dQvJTO2MGI/RJA9wZCaqWkELSpAyLx64YZEzocgXVnAmUvfs5rWND3oEeacbWXO9uCdCUnnvWsLa
Xqn7t1dOM3BDNIR5Jb+hW3oEdPkRIfJ3bPRDOH53wHJMgajsgbp5iVXxUw58ECesTJKilTj08U7M
Efp99Euc8qp98DMLnY9wh0UPybOKjxuESiq3wmTFosmgOeoHA16HfaiI1xPSqBv0VhskCnhPfq6y
M2C63H4Ec3E4GwqRv/ZUlzlYBadrnpwWGi8JbZgoB/RIBCdfCtbCybLB4yI3GCJZ08eftLWF/ddj
/u9SvzKMlUslXgO/5IDZDhvae7WCFpijcZHI73uGQjgakdFPLKXIl6KS0QLZokVN2fp/w83B0SBI
voaO+Dzf+M1d2NiARVnJiO3H7rkSQb8Ns0zxK/Yg6jCstvMOULM/BoP90TX6V4wXOxrnH3iV/lvU
ZRHAZXdo7mafeT1Q/ojvk6fBlYublDIuFmlt1kkItvOUSrvccj7VFIaohXrXjXIsH9+JhguX8F1I
7dm1Gx4Nc4e8CeA/qs4m+gEbo9Iy3z9Bx48yEzHPYkGI0/UYIbOmjmfc76RYHwrjYJ6+CW9AasRD
DuLCDHQHYaFSY5YrFCfLItcvzxGGJESGgfxp69esEMc2VJS1b3vwC1ctn2cVJw9C9CJmYpyOoyVp
dB4iHA5VXE/H8/MxHRMHt0DnASptgUrjLG3KviTLnpEpANUbdnlqlpWfa0NhLIHz1718oAWFiyQa
msEX5sjTISzU+hNo2WIAvX1yte/BsjQjstaKtyzLkVEQZDXJo+L+vr8alH7HDQiZZAXd7Sl+VlfJ
g9OaDbqW8ZKTnq2Y8Kop+8kZg7AwrDcWYyhkJNPnoA9VSAeVGpS7MMBFSqz+eC+RnrQevSE1jU8z
5OKQ4XryEJwbHQN/Ww1f+t1iCWju16r8qeJ12C+75jnZujKYwLdueNawwlRMkuL9AH0D4ESU1au/
uFQPG1EdPpcpzQRdm3DXXX3JV2j+PfVrsU6vqVMkwkLJ8vo12BgJgCQTSpVoHnxsQ5Qbv/9jDsVd
A8bOYZ7Nt87ugEEuyArJAkXtvx+8fpzH6PrrvYbdmA1CMFnLIf1So/3QmJYYj8SXnnF7xOGICm8I
wNlPi3wK48LG+XQeyHJDcinKUSv7l58vMf+/S4qvWpdWD/lCACj3Gh4yUCDcACkw8VA+H4gixHqu
dXwL7g0KtH2gZxSyhbT1YaqJI2KA6hIXkyvo2jiBaAe0nE4BLaZJrupnrbu8g19KmV/eeYMd9fQY
rR4uFfzixqrfDxEuDTe1/eKGibNDamfs9fI8Vfpxo+hqnGuOn7UkwIprykYch/jwyUmcupNYURtg
8QAYdK2Jp3EI1gMOjqJptewjKuenlTo7e7uAd1hJINj9SIxL8LZTsSJxVlI3BTdnDzUgcpIaBqBi
UjrMK+mZm3z6l+ePAIdm3rrrh9Fm80aHgfQbKm+tIboU3uSgkk/OxYydD5LLBDvo1lyB2dHKWcRZ
oFbFb9uL8uPlRJ7q84EdNh0d8KuWtnldR8fWvINX5uhLyk4J4goJLT++sAW6EmCDuTTtSTudJEAE
axaM8Zw47x0StfQESNTm1WiGNBdWWqtWjNzHogwUBOGm3dj/O+W5f/ocNJlUTtxGNdlCOciijfzH
L5kjm8lPkEE4PsPl4qpUNIIo5aN/v1DmslO7mzWKznuX4hQVEcIqO83gXE8P4uq7ZsVV2VuWocpq
qqSKcfPLe4d+D6X7JtGTHMmDNgczRfbSNJxEVbfsaZCqWUG+uaexzbOgF059CWzZUIz7lc19lMmI
0G+dJdQmXWwRieLMy4fpkgLSjPuN9cFGu9USV/gWlpEtrS4t56fcwtt+Z9oGGUM102QSDMG+ErbI
PdEA+dJ1i6/AMevHoQILAga111uLSUBZ3b+DnNqei72NYBxhf7Lwdv92yIIqhwZjDYikn0aCRPmO
H+cR7t0Y5/fHwOtkTk3g26cg8oq+2CmzjSKr5cfQHnfV2+MwAElJC+HMOFHg79lKnMj/88LYysfP
TIvWv6xlzc4zIGmUzT0GqQ6ur04m65jrTktjn48vXspOruVO4x6v1Kn7RbQJ0d/8cPp5MrzwfGBa
vuVjrqcGJUnUEaW6pZGUvgLxmKY300uwvKmpYLu9pmC4pVQfgPEg6jf9FpqahiinLU1IMvsuoTjC
uxQDPy+3MvL9WKn4K5kZGh+DXQwgdtxESQ31pnZbHdNETGMbpIiis4N9NhQY2EzMPFvAIshS82pi
boqgXu05QLh1J9a0YXdLIyKfTlkQFzh0G+hV2cEOXFSlDIH7ERMyM8EL7yjhLTNSE3teRAxlAgZW
Vsl1XCdgdIBbN49HYnvrurD8LNNDuMdSKoixtvoRqKtxx03Y6WftCEE7BZ7rl/86DoJc9XndlBvb
Gy56s0wfm/l7Mxr7yoDgdq0Rd0OFroSjlTmHmHLpCxZG/TANWtQpSTcdmkuiwCbTHXdKGDv+CWQ7
SreFMg6aQb2EyfXnt9/kdsky8v34SWXSnqPRVedzWVfQ+E1UuR/QaGtBt0jIPAHH3JEAxhKi4INw
VAXeDiooFcvtepOQaBHYC7B4LbxzKQOq2bBRY7MjQ0MpP1+zLRWErgxueXdUdC9tQpAu5zWdP2+t
XPrqtGYSlBqKyUaKOHfDVTBfhy1It8LeeQhVfD2tE0m+BL+Y9ds+/EDxoBVIxfJKswS2rMWuwJGr
sysXgpys+k1EeGYUPRh57N0NuaUFQ7eS6ISxdxnB9hsZMAOffPk4/BGk9RusW/Db08D6KQQ4j/2y
ii22D/mv7OvKzRj6G7KJJllyf2Uo/AnKaAldNAaD2iDr2dOEBVVJh96ZdkKJwCf2P/oAJDC/YK9K
yq7/K5ThV7/zj4pjDZxXxJC9ER2ongElxKqVGjCsAbUqRqViDJ8WyYk9T3uK3uHMrz2uexM0VCVQ
JyP6YZ8Dct5aG6tJGwKu5h5ixhziYRupk1PipLEi9wzayLzVPFxesL64JUeX8s6dxgQVNuFjuhDW
wkE3bdmAcC30IjoW7ymgJUx35+nuhs661aCN4j83XckW7vZSg94iaKPqaLmTpa6JF5g3GGS5Z0Kw
Ih+8ocvq+6ufJv57f0SsFQk6vbtujlwziF7UjJd7LzNberF6H10c3ev8Z9mOQrrpQkYuab/FvaQf
9PP2PUTQAQetz2AiYsjFdEBP5SJYBU1HcnH+ctDPodpFqs+pFZqnuJdanrKJjwHheL9xDPdZ2RoA
+ly37YOJnYTRde7eYXmSiAo4hQfVdPYqXo+FaNJhSxvF3uiQ9Zju3DCKxXH+v+fQ0GjcHdrIeGWv
LFCNM9PeOVc2TU9CYo3fk6zuEC2isNbZkSAu9OJUzQMwgblOTLrGvKzAIK0VwNFavbicDFfdzk0h
73h6/odDHxW8RNVsqBXpUvriBRL9J0lApYMX423WiJJ8eu+YRCNfPboWAf6dWzwwP57k4WckjcQE
wqXhjNsF2TCKz8gyo05Xg/CWaN+CtYp/ZEUGvvQD+MOkCbrEKWB0KHVCuhSG9H9Shtiu0G4v3pw7
p4rw4iRVARY9cdPjpVwSGylnDkypudE34vsDp8rT7JWEcHo5wCGSMDFEQXMJGModzL0zdvorqD9y
5XzSSt/hI9ECxkpWUioOaGrCc+pONOO8EWuUFSicO7HjHi7FxKFLwvjDJfk1IqZBpI+OsIpQMR3I
H84lThXINcX2AvfLmD7ZWjbXfXA07oclgrSHNFtoaEuNq50KhNMr9W6EKozHfv2fZCVOaERJL07z
VhtTfFIDgv5sRvlyFe4DnCDerYYLyW6BriH00Q7gjOUxE+o5x52s5/NTf1pv4gvC8bzE37YpKkvA
lad1hSMjFlxnshfRpUbe0SaYVnZLgE7w9uhSn4l5q0egdEe91GaUgB0KcXfdMGXC7g36u5ubu4/1
tEXbFbnXmGjxdJBFdT8K03xplTIQWTZMaG8o/HIv/0ZQM0ePU2/nZ3k4qtGNdXmHJnSiArt66jwt
IrJvkyXoWTmlAv9njmj37iufuu/OhcHF6smaZpv3Y0DW0eclIor1xs/crzLipeWyR8ZEhi/0O+g+
QyORfmZXC1TywXGlgCiHfsdPgQtYUe3LOYKr+VsJBHlSk2gIEWxf/+GH51Bwgv1dzYM+YF49a9Qa
WiQrIivCUYAejdTPmZzSdQU9SVTY9l6z4oFFvW1+dP78y3i1cLSeET+Vt9HycHWRPaslbuJlQ/o4
vEb2v3wId+UeM4NqyWX25r1nYG8GM4N3NK8bNGUwouDxw4j7URFXV3HbvzZNKKPu5nmTP8d9OFj4
CDJp//+wM0nNM8oWgkj3M8EXW2ZruGE3txGy0knOjp+xNgI9jm1gfJBYkLXOt6UekAWNQq34CoQ2
Bn8Rc4/dX89qtPUezylCjhzVm5NTPR2Cb2MRwbPycVWj1tbvTgwMhP5xo8b1JWzigYl3QOpW6MhJ
IJK5xNw9JWAwZ1TvlXZ2tZ/Abc8HYePqCsIr88WNkQKRYJg/uDxnFmccyajytvzj/N9I+l7aFQLi
wZwUkk3WlVIz8vtHx6yP5dTq69HdXYDMnDRdKFZKLe35cRASaqQyw8GmF5ZhkogWOrL2AJsXiMlg
4mj9wVGkT9h54W15JLAwFZ6+RL1W+5NKYpc1ZlNBLNvlRir15OLjx3BtOFb6LK+CuGVTjbyY2g2L
hqrEcWtYprvC/ZsdRWqouvwG4sj2JDKX0/eOkmFX8r4QNAVzYIFLf1gnmsI4CPuVRIAimuPB/gFO
YBEc9dT2w5TekKrRgt+9mzVV7058juk5rzHKrmQdaaTDvycFWk0Cah2PvDIlfGHhfFu1VWS4tR0L
t6s/PYp93mcm0QhoRKBXpGEHdi8mPotbYS6s2wHBDdu1tad6mv40WlWjV/XsXgz5g1LRu79++Cyj
LBcAvDNETvoEsF9whnnQGLgrb8be5iPgko4/QelBPUTYnEXZjjgfbc6iuxarN5JMFkif2hAWqe+K
Xe2zhmG5mmBiIaOBNn25UnFnzqZvhT8z4JTdTF4Op4i35t7xyTQMxCwuYx0zdPW/wpsX67oMznnr
y1cnuLpWmmU5N/w7GYbYRVxbgqQBUGmaq8htlqqWxOLNdtIZUzkrswK3C3XNgcDa7W4FHKWzbcz4
xVwgJWAyOhS37iXIGPNgEmQMG3ZQEb7Fc1TLYCka+fMp01qP8+7Tu89A3fV1cO005vJ06il43gBd
zkRqtdbYMPstO5EZjzAiAUB6hXcmzlXNVNLOqcFNkF1lh6+cKHI0WxFtxRjZr97CW6WsFIaoR8sk
xAZkI4fKCzDBEIDvM0ng16/2K7rECxc0YPg6q+PblzgUXDu/iQttR/7k4EMkZejGri4L3oR8vc68
PKZo2e5qXwXqaRE7Aslh8fy3cufWMHLLCKAdy7+VObdLsz+G1RSQ8OVmUV3SlO0UqfzVtl1qBBuC
FnmuF8jBmCngzIB/zq4KYC1Ape7PnKQn0qnBhbL8zBIJ9IoO7+VDNFcTU/7s76K37/p79Jp6E0Bz
QoniI4YLSQQz5I6GPvtpVOKLbjvOzuVMv0LjbQ7xIstPDyyQxYVwsW71Bg0C/psBar6W1hqCWOrd
Y+lPEf+FGtWhTXDISn/VX3HZwu6S7PBiK4ttlhAarewM8x6NsTpPm4AP3xRnqhFT8htYY5ToulEk
pGwL/a0mAnoML1acXERJAxJuZWTw5UXcB7b7RTOsa6ROJbV49+J5EaCXOI85c9CRJl9TB9yow2lQ
/+TpgMhgJkcDBvaJLce4tJdWS39ro10ZdA5cyohJizYc2bSyS//SY+NIk41tiS+1EC0BaGcYP7Xv
BPLDZNtptReGM2VDzCAg6UlSAwGIhYu4fttsIhCEACzeFtnugL7KcfQbQKfLU/eCAg7ACxZ6rv5a
0PpjqjbCq/jDzSuh7vCriiE4GWnwxg2JT8RGMLh1Vj1sRtTDjbHVTpGQkJwiI3PVh7lkBKQ40Dfw
+Y5UON4zr/NxYZRG4U96ufrARgucxFlSFKDny/i74k/nfyC27sK0iJmXI4pXrqGctUc8KeEP0pDG
U/TmtvLfGwVTwuioDoe/vEXMx9ULN/IUbZ9zKPj4ykf3quC6uJak+L8anAYAQQ0Lag8A0f+dkgXz
u8jIjvGBNP4+Bu+46DO94NKwBBbWOMYjXixZ+3asKxwe7yztHVyGEJktLSNFb8RZu7Fa5ChIMYbY
GAsUHM29R+uz9OIkX03o4J3G/qHpdxlm8YyMb/BaB48gBTGNy36sx2LsmsZ+3xsC9q/juZZTO8Gn
ghkS6DKciS/SwfS59Y+wWE6rd2+GiRywAoHk3kSmrJvpBtO4QbhafeiaBeBwx9lyBbGJu8hcpxgu
qWfhua9nKZCoZIj+YlR4RRHa25ZRp1AeaBLaD0KBo+5s2M1kFhMXHj8ogPgDoKA7SOoUJtp769nH
h/44f5XFlw1XMcAPnkcIib3iQqnSTLen+8V6Y4hq076/jBjxexnIBEXEdYUg/ZCpr51e/8H8VfO+
AckaoxU5RsPKtFzgkjGug71FPyL8hwPiWN5e/jhdRps9gi9fYom63xgbdMs99xXzYg5yt65gC4xP
98OHqLpOJIAHhpRkqKLErqC5qTLaztnu9JRLcq4sYcaugv7g/48cdfHZ48gdVe6RfUsLsKcLPQTH
OQLmYeOJXM6qwP98pvNDGtJot4vlQ9U9owtw3++Le2cUxFbeFdaS8rGHAeKJxyjCtxf+EJof0V5a
t0/RU/4qa1JU5k/awGqrCLif6vCpaMzH9bNFuVnyay9LzPsmC+Q7svq6A9l/cMpZVB86aQqDaQJf
znYT1kCSY8979hHUfTRiG7Y0FsbnP6GD23W/jmn64ptntszU+IovFJ7FQLo9zM6vTOk9joyL+XoE
jD35SwQ+TExLZKRgnjcHoU0VFjkuZtJffL/bFQ4OhF8Dhzy1zCgk7g6IKSmL1u7Y7EGnkgnCe6iT
HPbm7Y26CK9wHlJBko9e2TV1rloqhOGn5llcbBWecyqk9U4qeMnT/N9w0vH1WTwngud8wERUf8Vi
kQlEJ699VYipC1kCtMvjNQjEp+qN6Wc3ahqWdt9wog6FSeeqtG3SqRnu4lYhrR7Bp4KW/6oh9geW
wiDu1HuYwAt+o9a8jez0nbcb24TJCWhshWkAna4KgmomCechyZ0Yul1z3SyUbIfRe3zHgd9rSeVL
bH4FxZRYM9lx7oEn/A4ubtMOrxUU4lfbnFwwei/NqcWxxvwpdpaJmZiEG/UwfMZzPHJFdaZctr1E
CZquOEhSJVZvEDxf+9xvOQBwUQCmROof+zAaCQ7MN/+AM5fH/AFHQFRmFejsXkq6xBDFXupqjaSR
ANUzIPXv9wQGdgPpS7qWeRhw1ampYkFL5m3S5eASPAjeBl+8C3nBc+VAie3B2jqvA9fUaOFpjIFH
3wDv2ralegaZx8vdGXyBUUrdjv3WVrKCm6yzFc2wsryThdrqUEHQx4buW7tUNfELwbzIRm9ekBXN
acj+hJ/0ISbwWTZakcwZ1sq/hU1hCT5w3mcqzmFnHiK1pynQutq3tfIfV27zcoE7kxqExSk/Xu+p
SqjINcrUZkeoDJiAEZAli7w6kfqY73o9vmDuScNvE2Dz8vfdkDGl4O/bpFL4c/Ae/WeiYlUq/KQ4
d7HC03VA3G2df4WX85la/xGjPZy4dqCLlvkotXyJaeZzOmT/r91qrFdNJAHsBqMuUIy57SnENzvV
CZ7F7FYcD6fLAomRg8PUR3uHmQEsGhffI9pQMlgyK7qoZRs4nv79vPP+ezFR8+A9e8KLBpl/gOD1
16v0wWczTbu3YzPNywQG81D6rgDxNpfW5jarVW/qrdryRt8uVNvc71xddf87JB2XSvv3Rfll2COd
sp0W9f9y+LwIBkooyyj56psZZ4O/UaxaLswCklS4iG5eI71/Xz1Hi84Mx3FST3gq9G3AGCWyyY1j
gcY9FQkXj/PTuvHiT9JbJ0Wr4KjLN3LPbLR21n6aKzqhEo4ZwXzXqg6q1yMh0HoDznHLg/FlsB5L
JkAW51jvvSi1iABCEG9VFLSZVNRSEtMXDQwceQ+wRT81/njcKFx2KXOD5lcZPKAH3I/OLqGHP1/P
2ccHAorsmslNlOslRs1kgMKiCmUXGbgFl0Z4Mr/7WWEbFhuRsDglV/4kgcjbKB2cXOly6czf2GBg
WeKeOC97IMStCmC+PLMmLcFNLzg97UnXiw+XL5BCwvofANQPFZAF+I/X9D2t9CkXR++FMV5VTvSN
uCWSl7H4Dvvlz2w/Nys/g/FqqFVO8ZxI4eNtcccM6Lbd9GMBC8IEr1TJ3PI7NfL+koF3qLjbqF9U
vbTPr64bULtxHHTEP2ZA9TTrKYrvYiW1zyEOguMrschoVeXNPtfWTq4kB9M8GVLcR/Y8VOx81eMj
SpDGl3UMvLlq3kh7jU0+Jh1w5hSvHp0oXi8+r4vk0inFqSQbIyG2vzp1W9upGY0D1BPQmJk4oXzJ
lSmE2T3/ZA5c2+JEgWOzdeD3qYJ/kA+4hltUF7nOvAvGKjO5FSdBSXHaEnE5LjA4NIb3HTlCMdN8
XMo8Nw6JAGse7KWKDO2fbEgtXp98X/tkjEUUt2KyK3DgekYJLYnrIUBLYnb/W/LdAectnMwqJ+j7
mZxpKanYi6lqenOFQQVKYX2D6xKpZrPlvHLA0wO5WX3xq3FTb+BkVs8hPpG9G7eLvW8rWYuXUAT9
tAyu2gI19s73RVvRGgiL212NXdnCeQZwZPXOAufaGEF3MkmfL/y3UijmxwoPLdopHpRcYwqtLWc5
VeqFzG+mL5Cmdo9KqqhByfxajmANwks5GcZy/ze0Dr+mpPqJ3eDU3qE29/9+mfz4YoU1rZfP7j6c
LZEduSgYjmUO/TeQAjv3hapn/WkVRkJfVxLxGGGx8GJSbae6cHa8xkElNCk2N9gKNJ5KRp2mO8c4
fHdU/QESteWNvI13W5czaiAfp7ZKU1aK++lALwuBgg9PLFE8FWMZyFtToZ/ENcLNdTv+wGIc1Oyr
8htnUdCzqzxeqKupN6zv7SiOYN2S6aZpDoRoilCtOcZuhHqp1HcFoy3kJToWC9xIJnYVPnL5gBk9
qQR4+6ZYbYvmMMuZ2MOe24i7Aa5NGTpWMu5ES9io9qf6fZzQVYZgCJEBU58SbGiMgmkSa8bW4zY2
VRQV/2L5TaumIlNHN7RjbQFlv1yAx02J1FDVsjPsQD8lhJ2rrqq+8949ulchEIveCf1J2PdUQ6iJ
xRZXjjrgt6laki7MVNDKgApKhQqBpHFjSUC3OnsrF0UoOODvm5BziUHexRwvRIz8kRp8b1yMk/Yv
uau8yBx8xWUW/hdBtjJaE9JhOmRHgDt5yVL+tE4i4a7mVCWs1uOpTU1F0slLV8/SbAUkQKlo6tDf
bkMBRS2xd/QM0aBwW64GM71p6HOWwatCE20ENRH8jjUBcqyRLg+hY7YH0Ps0CRVrVPrRJhCNTety
/dmw3fKjDv8WNJd8cjsnbvY/CO/XqUbOBcUTfbcUfzKjZNj+XRRq52OkH+PJ73x3M9r2Yr1o+jov
ncbY4dsUnXN43O7jsFH48y/xngGDmWa7pO2p1OeWHx4hDX9iLb1igeOfDGfXILrRl5vdAg5KdeQA
vY2dzyPgd872v6nqpPCuHEBoJZGdj5ZNTX3gcIxXELkEMjL0uJQAssuGNv8C8+n95EKKorUomWL5
RfwGnr4b0VqyoXRKw/c7K+7YfPvtRJGzwiyp1KydJVxmKRurtL0Nw54dOXbRSizAZmYYZWH0dRlL
IdE2XhuimYAo/4eWhZeAC9o7FsMcr2xtGxO4EpNyJ2fBz+fDIvKQoSbEZpDFcgaqp/Cm5tCdWUUM
2vduERPps+o9nsxaS5JVY0Sj4cUiBpwpAoGlokQm6i3qZBa1/BIyLFZbcsDRjtrv/9G09Bq663q4
t07hW+BYJmQ6KwDcgsVbClMDmj8nrKasSxJLF41nMzeHPppTHwXDjld4RqYygh1fGBAj/wsSIALF
sRC+8X2y8BAXvBvvyIeSO17yFzXuSeHUxy4rSuFspHYZWabc6mJJTpoHv2TZiB5vE9jxPPdH0bG4
mlzMh2vZ4wUW8uvppDz/IDUJGPNZPsP1ZJdLZzKrsvU47KgpfOgNFaTFd2mV6Xi6InJ3Be4gU8vy
MVyU2YlhrvrTzwRw20jZgPn1TJRDN1Dw9KskYynul/ndIPLbusDzeungLiQ6FHKNBlOhwf8jFy+A
9SzfoEZFkVhykzzSyvp6K+Sn3NAVfHOFE+ma4dqS7P3/VLrLZALm7WtzNkMTd7GwdUV52WoikVrE
DbqKthUU8ks1wvvq1LJXAM+j0MEk/3NYaPtWuHoxPmoreyRi15AOC2QaZjASmlpM4nw6KDIRohH+
S4pdRPlGFqexrW8pKLfd1nIn4XVnfZnDYrlZCSFygisy/Vd2h07t7Xn0brXZyrIbZsdQ3lHpTMNI
66OXTwo7f8Vihj8lwAY1AGOgeRHl82SYUdq5WCd1LetjhSzGZA1rAo1uNn6snrnt5ezt2+UXUdNY
ONTgLyJjRk08fXHIGU5C7hF2aWX8tKZOnZJtwuirHUpp5wDZfdoCEJVcORCfgL8hos4uJNdC85LW
bquaXIPF1ZrCSc0GKVqAXxqgytfe4I5nSesFvH2HVLvhwEgBzBIIJ0nmhxlSS1xHsdPVcrorLLzv
dHr2/JTTlco2tgQzbalk2voKrVYrHW6e8EIhLxwAIfr70qGn8v9Spa/2lCoJqnPLdEZ/Pz68NnJr
OgdxuDbvy5k/H8nloqZ+BzrcjF3BSgRgFU+4Mu0zS62+GftvVnWymwp6pCI7ghkIjwO8JAUFXqAo
hYWOm24Idy9mn649E+dP/c5ESujoNBeswyeLVCieOPLa8+CYICAjFU1o9Qp1xw8l3wbyMJJqrgJQ
Z1Y3+a606bECqMqeeFx4u1MzAiJfqCRizmGxDnIjVyYEwzsEqNboNW/kqpbqwygmf6tOsC5IGo4A
1V4sjLP4sKbi/TgfqUGP2ATUgywMAztdmNkXvCc8MqqsaK+mFNAhsMWgPwyl+l02q8rXIpvxrhg0
3qIM2XiGobUCeouLEOq3aLd5eO0xL5N9wxaFS2xVcnQx+VodMy5ac8r7E1gvZqURBukOSntDVx1J
JarsK9Mna1kebj/fO2g1pegBNWuQluOZ5qxdabYoVAFxYYWeyYZ6WDIL4Etwo2dkdzWOF7FRK4vp
BHE6k4Re3q8VKxg7CJXHoIMT2WKktKVYQJdN7HWyJGJMILDQNmXVULGJBDcbDXF+kxxokYYeTY4v
JJrftJ5m9VK1Lw8XEXxoLMXQmlQrwtRTO4uo6lnDrcPHHQSHDBdKDne/F4ZikKaw40I8USUUw7y6
555cy/a5F0taUI0+fkNkjDHomThoQL2KEP73RE7a6uJaLsBmnKmDdgCPJXDZoxRhFdpdFFO099yi
06L0OCk92Fg4N0mEgJr5Otu9biRoxPod+WyJ7HlVrrW3nXQak+H8ZnJUg6A2knG7eYZZGbdwwBpa
1AYtLkFj0d0XWHdhp6so0UgVDKlrm68N+FgqtmaUCkrcaKlqSIxSMMFFPsQA3sNuQDbjthYox4zM
Qf+N9+aMnGzxvSTbx1/ViGlex4gsUbSsklRtYFmiVdxPSJJGsT3p7piMHwPaqvnAWr90yAXDQDaD
Yos637JhHiRf89RNBat4vgl6LWqiB8Ne4Q+a5dr1QPehzIxIut0PE7ulWIzyDqwVEMhExCCr0weo
LkRFGAlNpPITHCEuX/IlyR4xhynGG+bksWVMGe9avAGEzObsYrb31eIP7aCBI4HDY5D6QfUCNab1
6J+t0R9g/f/jcTeEmi6vjwGe38WBxrb8lg3bloWlD4COqN7gAkNVS60wDyL+FUEk2NiKzYquo+I0
WDkfYO4qzkstR1DAVX8OLpgRvSjL5Th14OR92QXC5HBDRJWwDER3O/AoHcFfQ8MOCWZcZsIJev6s
zb1gW7wS4Up6DdmFiJNdXLgR+CsoIBz0uI832O4dEfeUGeM8T09lo/n2XstjeP/2kFb9ispAyf5W
qWfMi4ZXhZeOSKjyVY7Xz9F83RESR3cOWCE1/fuDbRczAI+0JbfOIDZQ1OTPE7UkwX91ALWXYUTR
JTAY46EJdCBgiEUIcQnr6yoo/U4se4MVGZnk6+SN38dyRjbC3Eff0Q0e3mA3LUNNx0wbqaAj0bBm
DwnXx1J6HyQCfVrd08dAqqELYMr/cPKNmOGSzcGpFtmFmTZsqSx+qZBSrwNjSIAFP15MYhXVb7KP
XdEL8U6J4ncAiHnpioh9MdRVBW4b0aek8LgnVktoSDXS+puLm9hDp3N+x6ouQZDdAJpwvHQu2uIa
VuhkXBdyk6XHJs/n07U2o1M5TjYQ0aoeG5HaIzcbJVExvGoYuhUHpoVqDywhgGKudRR3TeDeyBMX
eyP7o+uvQIK/r05JjBTzo6walG5Ul3JnK9tklZZHqoR+t7/AytBUeLfR9SGX0eWUqwtlqctWHwy7
Q9V1PnS8R5WqC8H8NUmTHbma4G49BXxIUqBd/aB54FrMz0oluvNw9FqASsyF21OzsWOBbdEDzv0i
4+P5AIgREUBH7k/24aX6VCuJhRogUvZyVseA24RmOL9ikPL8LGUOnTg9XbeJU6bNRs5fSNgmHepW
tZV3a92ZLkJBN7gnwPPl+VfyUHgvT+Dve8jJiCxz7H5LHz4UpgQ0NJmSkZtnJRAov4UerofsT+I2
k+K7JPYQzcd23Alb1BcERsOp4Qf4Pj7mqOWmBGJcxsPSrQnqkqxP8PqPNK80zQHWmoyaN04bhnvC
4AfZ8UtwhdkMuhp5v7CBWQu2gchTSjdV7l5sFKL1fK3DEpodY6PQnWGBXOgA/tePjIgTiDCx9MJF
jEvvCSJ9GIl0SoRqxJ4tTP+kiDB6KRj3iWaDehmp3sr1y8dM35OM8aebC2DNblyNQLaGTMWW3/WO
OkFgiowLxYlB62JuuNFw/lZWca8InK7TZk2H2wmFIBkOM2waTntd0ylwB2zbhjsWcZi1ps864ccg
f9zT+3Cdyo5F0nTpy2DxweE0SR2MMYtwXvbD5iQtBGtG0VTPiSqUSw62A+NmxF9RZ/x4I01gSU1Z
hdZRA3aa8S0wggFBr7ZGcoZRnC2TjJQfbqjQ9aZKvK2oLGa42Y9VMqZjv3YmbqlmUd+L6PzNOLlP
GXz4X0OdlEcD3ITXJ3GBO7XQmueP9i85BKdRFrL7ynn60r6ZjdcsPW6D7xPY6ZmanX4VkzRqsBO4
UgYrOHVCAob+KSU3q/+yQQ430uO1FCfdwK8x/ye6ssHlxRmGogsBs8XJJ+95CHlcRELb5g4EINuD
mHrgszvismg2CbzqRormPzXP+un8pkvyVWt0iVEIAin8XcjmQGzqHEJRIkCW68K6FT4NjfL0uI9B
2oqkc2Xm/0L3oHrnmHOb/iQdhCymkxrDw7NBiz10RGNvovInyn9i3T7OIizUQUYFqG6GUe9FAtWD
U1yXLdsb5m0WCNGFOk7fb/Inr0b8WzijvJ6KY/A8CxKqLUtnzlBU+KFK6uSh26lLDd2C2pvz4rhK
c5L7CEJ/LMxKufIYWRyy4D7sMcrQvz31nx27rV97JG0IQ4RmZzv73J/VcoM9oByVO1hCe1ClZR3Z
TBMPSsxDoXiGI2CoDiIY9yGQG8zd6LgFhij7IFBA5+k7Mf00VJfY4fJa99eGq6zNhdVP+L7YGR62
eNiICGuoL+1v5xtY+2sSZk48npYMflBK51d3mGHkFOYBBEYHMJH3nK7DNJSWuvo1Uo8bBYL0d++v
q8ceWIvNKRQVJ97N0INi1sG/ExZYZFa6LECYz+LW1Fj3mC2/RX2+efqPylpLzAe/MWvueq1gv8MP
l5KEIiYuNquyCr4GzVvN9MNLhlzp8F/+NxQ61l1nYXoBesvX2Hd/a+3HxLH11iIMojX4lZpLN5Xj
aaWESxNVik9mWncyXWWltKcUmGsIwiCeWdzJi5EZ6TqiJltLcFT5koqMBAUuJza9xCmcJ72zxWcA
RSwebSXG945HrWUq/9BXNvIRd/GuS+s6EfPLuJJJe6Cd6Gpi7dUCZjEX45oBHyaUqILgaYEoKQTL
f9KlZnVnnI7ZOTc4kh5v/fIeDhWlanbPLgMdB43fPmalp4Y6UKUum5kKitzmOzVkbNAxPqUvpCz2
IIAQTgY3SHHwdRjFMsHOfuUWCq9otwSYhRnDv1gpXRnw8UxXTiIwu6ElsMxQbPChiKcAHqLCDz5f
XVYKsHdPe7ksqekJNm6h/nCJKMO9XIVEmdrElYjvk3JI0MSNzkNWqIokJhJdU1EkefWVP++JFGYR
MKuDgtpJnfH+4JCSN7ducNRkG6zvbYZ8/Tfzwj4mj0ndM6S/9eZJJGXqNvTl1zV8RiVFSmxP64+z
WIwg02Oo6qJ95RkhYx/8nW/iJqm2brNpS7alJeVGqW+q/XQVOyIe5m6K9uGeWIlDEmprxZDalLX8
nI6u15dKKIwDqbepJtW5D5fvsQKoA8l7JzxeffDQhztOVfRIEKC8Lt8jIp0Og5/XzdK1p5RGk0Ke
iqA+PlpOTd6NZlapwhxI00j85eMHEdWW/rRCgH9Iiq72BAxq7K/6pBEIELjXTdQGVZmqYs1GmIEe
YB1JQ04DuzpOXH7y21ok087R78J3KsB6MFh4ajiBrUkAGx+clcZCoaif0lu/GRlYrG67f3l1ywzP
nPbUpv00+ezIq1aEpZ7b4zSc+ZSv5NXNCGzWeOCeTkdEhL1zuPV3elLCzbBY3ALttgWSkCkEev5D
bhq9yIT/9CF0/IB6L8WklTG1LNnOJiQAbA9nYY6zw98S7yz4ADiuSlZquL9S913toh9ia5/LXt+l
xCfzrswE9WeWHkI80npZEVGe2xegZvLxPPpi7eNlCw6K0IUZLD1M5i4fExvVy+HJgZUowxqSEoxM
eJc/hD2C9APYLaqwEXEGwjw4Eq5TPuRSuvw7rCnLfCEo9Yv1qus38eS4u+bzFmWDxthf1jqiORpv
QuG1GU0s2Tlh5qXwKpKXsxN3qR7yJ42ns5+frdXu3D9/balCJ/tibXVHz7igvCyjJlHMlAhVBDAX
d+pycN9PU8a7WkQZUp1V1qBf9fpOtUxTiiIZAsOIV4aMG8SxLo3uj4D0RrxekcIrr9Cce9gTg8nj
zyCP6D75BppyndsDFdmge8wYNK/KaYSfNEjZ5X0YX3hkMl/Ejtreq95D8yt0VcnU24sFO9EbwPma
auT+oydLVVzgoD9YIkfMUrN7Yr0NI+SzsmAsN8o8no3BIlm1my0MiyM7mij0ztAM7ltKQROp6/0V
cA99NM/HKwfNlI+xKKKugyqAUrpv+jo5AGcDFEHaxmIStqA1CPsYB5C/gWmX7qTIiPzmJ4ds7XNF
2aXAwKh9k+w1gXsW+bE8UVRISRQaZvOwUwd3k5y8KsYudC5xj8PErAj+s6c9Jrh/rgNMVriXzI6R
+I3fhqHzZRZETv5H1irC/aI/GTsi6qcDuMKZ4BO2v8cv69yY9b+ZJWY/GmuW8SAL0/Fi1MKC+FlH
SXXD4r5WhdAHe/66CdKMe3xsiJ0zBqiPW6tHLfKdw9Vf5zB38xd8b5yGMTgZuutSwwhIUbKuVUEB
Zw0Uv+Hh69PSPwtrbNjgrYCgCxZcMP9D3mqQIy3l/tY1wjZ81lmUiY9WbrQyB4rArVMbcIrvMukU
lSOnv+rQ5l2v48FD7nY121zw18sByX5FOxo4als4lThraVMnBAT5qtSSl6/WJLaqQFsQhpIUy746
O/RhyBTYiVLy/IdOpUwX8unV+5JEu4FjQZyGu3/4FeaOjsb/bX3i6MoJoAyFxQ9CGB91nwHrDtPO
daF9L1AhLss1O42tYJkluQVP0xXCSarEq7uwiNqP+qMroU6zDvqW4H03d6+0tff9g+HZJlVw4S9w
MMapZ9CJIohxjjKLqZY2X9znedDujDGg5jchY9lHcNdw+FRml8s9CZBrJKdIRUUkwzJq1RSuiqQ6
0I7lCW8dGpblTqwytc9u7BYlndTtjmSU6sLjMJMmHfvOvCwzugv17I2b80HXvy5gAFKo+R+TAee+
As78+7VqTxbePas/3k1KEy2L2o2Od1ofnqkCXr6FyAw7EIWmSHrv+1I0S/k+1Svebx/57DsCb9o9
0+7ytidXTKxb0rfpgPdAfWnLmktvtImDJj1ShUWnbXL6mbW5jTmvGmsjZGqjxs0z8wMevCUQIi6Z
0oG/FIzMYXEoay3m6JXzC1HF5A7HEcs2L9BqF8mGJjhAE6KJU/nd85kGKWbElkPwMJIdTYKv9BNp
qzb9LoRWeAQZOXwEzJJB50iXJGkdhXK73QSRGoeEv1Cc1+oIXbRRMj1wKnLAvnyV4+n9fQIfsHXz
i9osDlON8K0t9dJ1BvhdTMGMep5qBu7v+hFyNzRzvp5rEBhgC5i4+1gbYxzF1JofMerH/8Ws9CWQ
Q7WFcxVmmtYgDtyfziuPT29nIDhCDp5lnN0zzEoHvOl4DwHn+2Zw2h6DQTq0gwLwm2u8QJEm7QR0
JI7CME2wQrm1E3NqqKdMVlvU+9Ts3saalAJcnEnbeeIo5VYmUYoPnS0qOO1+MiA4aaUCrirTMUr2
1VEtUhxuxEYei2QEQJCtKV6ym+pCMOeuG7eRQtwyJf+BVxa4wcDwZSS7T4XpBjYwV2HIuB3yP4Y8
F1cVA0bOJ+Hoth2+aI/BCSMHhuK7uIEmbXJL6mQfjYNeG/2jr/AkQYsID0WqHZGHxK839fYpAPoE
nzSB8N6kWmYvmMla6XSlX+aI8ROxvawfYiNlAkXoFQ4qcY3Z5LfBfdnqLAzqvhR/nfwUnURMK6W/
Lz51ulVgybOhi0Zj1YtqcsGWDayooyyHHrRUFXJChpnd7cG2KRRqPRfEnslbOAigNWvTFNzTKXH+
PSW1uu9NWcbqN00AL6J+S3h7xHE5+Ytj5mItAxLQX4ou5722migIm4BLkl3Z+tboRmUyEVhAowEi
jGtOah4EyFxozzC8hVNHUb4XRyQVkol9yd0rluqgPoW1nEFVBJpIF2ifRIUMGlJQYxIY7pkzFdcZ
5kjTRmrZ9ZdxNj4UhEmVRUS+1k/ASjKqLSfaj+F7HtrEOYxBR+pHbXcco/RUaA6NYnSpLAtjb6/R
UQVmDRvuELzZb1OmxiDH/NxrpFzUAUEEsgrOU88UG0XwIXjInyGtVydXJoMCi0tKJila6DCskzBQ
Yx+OlJufJMgsez+24nr5sHVgR1cc6mN0UTTGuvY+QUoJwahS6veUiKme45phN1BUq+itlzRMj/NV
KLrDyn7CieL3398GdForNGhWyRs+RAwY50zRg1hbW+KiqnWeBLh8cunZRZeKkoAfDPLiyw3LOjzY
5rPnTA7TFa7dQ39Z4xPz3OFjRiKIIa2qcwX/pYbWGkg+y28CiMw9BmBOfqCp1S/5/ol1sxLya8xU
BEwXmGSNBaOF2fcCqTDq0NddZrO+JFY8wZjATqgalzDduqQUr3pstXo1fEzMlF97yH655TfMkYxR
ujAkgLvhc92iPkMvnVfrJimpFBenogTJYmG8VhOnJUoC6m9xtHxxvq/Vxk4fRn3IElWDSEa4MMqG
S7XwDIC0p6mdLnkMPxJBYWgI9J/XkEG7ZXmnop0v8XYgNsPbsoPsOTXUUeYu3cKMJ/cQFUALReON
SLpOivdBSJOgn1633e5CnHEanmizMY4jIF9eX6T0v45roui3YwXLxXBC7RDW4LSaxb7mCv4ZvLcj
rbkxMspOQSSG3l6f4QpO9u8olYHQLrRzF0FqAl9QXDXUOBBwjEuWRy9KjfyCeuDOIor59rMU9wTw
bsR0tG3jDqshS46QBYw7bB8wTrReW7iwHzbeTsEp36J+inaeJYJ9hq7IiySRBdKiOwUzJyBpmTCY
f6cLO3rpIh7bkgawOeLPHs3IEn+mCY9ltLDzi8YI4PuEHeIa2VQphzh3RnsUzNN1Ry2z3zfbdtpF
oMVNOx5NmdXnxLbamwKvvPxVC/xjRG26oCpi5YWRK8R5CdKXsNLQiekzuHSCqUex/b4WSRlQ2qRB
HgWXk9Ew+6XyAKtqXbkfyy0g9bATolXL+i/3OZ5F5OI2qW4P6I5W0j/V5vs+VdV/prNPcNGKBGyE
awscOQXIixNG8FnJKBlyycgBC/hlcmu+g9qATAeJ6Vj5ZGtZ60HHvI8hQftM30yEykbwc/R2XMIU
t5uoAoonY7kLXmdpdfgJ28J3m7w54EAdCMqV7xyKITfxgSgrBM4GN1CR/fBtdbWXoIm78PPYZ2ot
ObHDjhnpzMexH/Gk/8mJ1zZI4xxQf3UBUusX5HRneNRDNGlotY2X9FQgDxH+QzTg7jaCXLbItJz9
YFAWPxIShhrafkYjhA4Z27ceit39l+HVna6Mz2xzNZaA8YEJK12FYrp4s0PKtm3fGmsEAx9dLcjK
KTVZC5PUVaiGRMTp56fswO0FSIGSDAwn+WMLG+OOJj/r06kM3NpAQ4hSQ0qiNIJfPgq3YDJpAbTo
3A+c0twkL4Ix/D31KhehjMcRXV2iPTjP3QvW3Y/p8IRJ0QFlb6UIou/Ai2gVqmkTjkJLDxNKPH1L
SFQwhQhhTH0h0JD7IimL+cCRFFu34KV1O5e8VZdt841iLg3aT/SU/8l0iAs6FnF4gcoVBhfCHzPP
hXiGDn3ReCGOsNy6PZeQCWTnqQ3EqOA7ciRJlMhjn1Jos3mWn1a5NY27uHuzsyO2bO8fY9lAFkuV
wodPGHk6xEkMzhDULb3464CQzHKqhEMm3qnWgiZGfCdsBzDRS5ahKy2p17SBbrTd4Jy+YiACUCMR
JRH282B9GcX5BY1T2DBYigU6eGAgcP96Ol3W1ykosEVVFy/JAe9g6oj79Z2A446E0k0C+ZuNXJHD
UVp4cHYJ3NoFzgXZnrOF3gIsjEDk0TYRU6+5iji1BzoZDV+SuVRxgNI8nWCTy6x80VX5kwsPyMPj
5YAhSejrAxfkv6Oxx54jDBo89qM1r9z7DdNXVeaRJxje47R4Id6Y91TQ4xujy87mHrGI/zGhysz/
Am7nkYC0/SxA5RmAHvujtprwHyEvsB2y4QJCaW8e0VeaFz5+elxjqSFTGQ2gmszaduy6wu0voZEr
altMeqOGfK/wJ4FBVsDJcZQeU79Dsy1VAGdBf9m6fzdfXXrTBDR/Hfzd8/+nbIqZ8J6oQLi/TCYP
U47mDTGnRkJIWG2g3nLqbvhGx0vJqtIFD7z6Bk0hMJBEIS2TNMNh+xMBdvQmAftxGfOT36xFZq/i
lqoDJ5IRVhCveOSCiMZa3lS/9I5Lrd6BaeUmgHffgS2LBNw6anHo7v63D6vNnK3agvg0Izo6hl09
TLrKsDvk3fRg/HaL3+NCvxtsurL2ItBh7R2ykIp9xmSVM6a38st1Nd62Goq1SzVj42FQyEYJM7Gm
I2j3m/LSguCqLBKsvjhpcqddxZDHz7FjRNhw61lQmo8c0EayatnKuxSm1V235/bUQLYdP/nfD9Re
nwjhVisYL8sbu/9i3f9xzZP1FA5ZbAkD/TnTC/9OkGJCabWXyhiFMAMltUT7yfkpHqflW/aM98le
73+UylULQcSpaTVeIaWHfxcuTf92iq+4mGbsu0qMD0WvWDmdm6P7+iRYfmMj1WslBFoDbQ3daDES
CzAYAE7oPisbiGZrjxFaOz+h0bu3OhIXqZpLkfQjEnTXOfQn4nKR+P4mYb9YF+fOuOYb0s+1JjSe
WotErSm0FlQ18fVx/9xljqvU9JYtPPCed6XyfGTG7gSWlJor2NlFuJpT7Jl5GJ89glmTwCCYPLWL
Opz4VJ/eUDg7CptXl55z9XYGC39Ql0O48PxChw8PM9zYcRlUJ9WI2aMhdYHCVMvZkAmTdw2w2El/
LMgAWGbw6YHk3XUuuYGiDQl/aV7gfiKCGlD67l439xI8f5cHolilJY+Zek0SUutcZf05angXuf0p
o6Y/e92YbDCo1h1mUtJZLFkg1VNrcyGUvwJNaRJILPXXILogROeTIa6//gBzrbmfBnJc3GoJ9v+4
hFhSsXwetzSaV/sjBsKYYQp+fiQ7CqSLMlZfXEncBHOup7k//Tb5hIHKAvsRjDgPWNnuGX5sercw
2QRQtiUKcqJGXVKA/tqZ9ZuDyYeDvrPAl+CkcCgvcIbUb1mkeyeYWyeyhiKCHq202VQEPxF5xEL3
/rEkmi2NNb/pKp2dH06oFpTXrr0abtlIMjggbNRMBrG+BGmVHxGzEvnN9nrJjo1nOKmuSRubnoAb
eaDCcaCY2zy8LSymahr8Dd2UyTPY/x/+ZYfLjmHGOFm9OE61/VPleguPROruY6nlvLYsDuCF0Gdz
6q/QozYOa7ol1/RGVLCxFYT9LQUL9n4FXV6DtcnQvYKQbogqUGDcONYJEbwCoEambfi1DlQnGcPq
uhWeuT0SJVzD5YkDBIioPfVWH/k3JK32i13Gu9fgIgymG0buToFeU7+vA3pvyhJ2QEDB1WZPd3tO
fgsAfSKOtx/cRHkiHRwkgjmB7RDxu397TGaiTB93RMgQUXsH4WBHiU930wjqUI0JuGg3xVcP0Jj1
cZ46JgBdLajV2gT15SW4YHI3yLm83Llb4SJRvflBppjL3lPtcEDzcXZ3ZLVZCok061Ai/Gglcakh
Sqh72xWUB6r7ckkOFKSpkZBo7xoXD5Y3Q/yfd/FiiCdcUAAO2PYNSLTHPQBqr+BpdK+Ib58gmVSI
66x2xjeuM8H+9EXloMy5vQoIOeBdL/4vky/xjMM4N5ZEZSxmHc3MEDIeCck8c4nq2Yhh/RX4lDrE
jVvgvfJmYiagWnEs0TiuUuHfSzkAE8Q58fYA1UL9TnRfD26+C/jGKRhcN9ow5P3Z0F0BO0xwqca+
/zC3hiN369CLHRZuadbHSrQ6cB0G1u3luJ+pPu+v3ieb7tJhR0giwMsNIVPNas/DuDo7v6qr1ns2
6QqH3NxmZOvca1w3yV5YqIiDmK9nKPQNtjx/bsWtcyCkGL/plU7efCbu3KYoyIhKYKx/AqPoSCst
aSjuCUzF1tqTfu6DMmHsuEU6VcUFrpVd0dV5pT0TS1ZJWJ8Cy3kojleHq/+BdEjhxUA4F+v+/6DJ
/H/5pL4R8vb/hQkixLmaVXJa7S4vZ7RNHdp3L6B6wno0OY+lcsS3bK0jI0e6aZYgaCsBTUX1bAUn
4bLTp82Irl+GA8T2oHluTbtawR4Q+LE/0Eww+dKhZfEax17ERZhC8pM9OsUCFS9YQOAsyu6M6moU
oc/KfxY0A135zCLA/q94gnIl4EoS1LpHplGRTxQJMKNj4D6UGRYS3dc/5D1RMy/M8EPGCh9qI3hH
164Dw3tiUBddg2+D1pDj+qnqKrL8dKkrenZyJUP9z9TX9ZAd7XgKxVyaT0yIF8IRh7pCKvCM0duW
8DqbO+LywZ5L8KQCo8IzAbQZAqylQRpSjA0h2o8NcfLCt7WMneqxPYgGl0bIZhudmGyZ+1uYgzkO
LfEFuEBM00rW3MF5N1GkeXI5L8iXVOqUh9+edY1rwA11W8XUH/amy6WpMuoxmK4JlWCYFGzrOUSi
ayPXf4paXoD1HtM/7rlTUAK7jR+VPoc11YtW5Pr4IiE+gBK9rTl9VflzsuU88Uzt0qp87RKB8Q21
gooRyPGkd+2poCCqKF6oaT0Y/UBMZxQK7DVaE4lF55zJDFB9oy8vp5xSOGw+vHEVzbbsN31G8cWv
vVi50F7dfTC7nipaCtAnx01jIpcVF7RjLYUoA3CHUgfijdXrUz7jQPsYBKRF/v9ZFe7ZOX/QRgLN
xI+xmEOvhitheWrOfgZKbdxAiXFAC+is86dg7q+xQg8IcNsotOd3kD02ATd1/1AWWpZDTxrwzp7z
CivYCVR6UU7eCdQ/BY5USQMHSfTqcOgkiUXd8fhzUaT08+eKINQRsY+KpZiz2i3s11bfYOFoyorK
Q16083dwi89VSHTW8Qwp+9ogSq8bTanGNwVVu6L0D48cilYY+STKvLE7o0kMAAZP29K++I9ho25w
56Eh/t0n42fUn2g2UyAp4YFlQhEWRL2ZXp6+Jbcx2P7B//d5CeFmYulGn3A+YoKxtXJQPkv0QgiU
jKX4aHfusVW/d/KNzLbGF7ObuU4KM6v2bHtiIBb5JwnrviU6Bw7WDFrabGnmS1k3aS6XhyxJgIHB
+3pe3qwHfGgaPTMgpgeG+TUaYNQZ7fcxhovRW5RyFAWJmW2SDkeQwjZcuSwClSRtEGybFAdChftY
m0BBnC4NrLENddU8hSGFUiJtFEM7X2i9UWHdueGdLK0D0w/BTaIEQRPRr4iYs0H5f6/P3HdtLyfu
PXSgWj2eMIqt8db8i6QglbXFPWq3LWTjY69894gB++3BDRqtuaLhjSLWVNVWMaQ7tTlW/Ls94MOB
OUe6KTp2NnoRRglTRpHa4dR4Q5Rm/6i1OYrFXnszTjWNy1xjc2OZRifxOFboG2LMxkyNJgU4CrPK
Nsbbntyw69WP5GmK4XbXDHgdu1t2S/zAah6vyYNc0+WZAeiHAKZk5Fx7KqtTu4XdPdy9MNnzAVdV
fOzuGtX10hbySxrySetSJom/O1sPImnKRd8W4F6GzwfFv4lY0oMU1FhW9gLMu9efKvLkeizXJ+mE
fF76mk5Ler54SzsG6i76HXxbqtVUcmF7pmDE2Teasni/v31aPUle0+WvUfjbWcRmCHs2U3dweBds
R2UIS3YjbiadE8H3R78Yb0fG7OLV6pFbcMbxDCrlS4ZtcElkCdpmjhXmlBJkLo+VPeCFuTtECXFp
iR6te7RerslmtjH35GzdvsxUk6qkB6Uvclp5/C9DBtfAK7WsjfuOWoMDZ5T3Mf5C0Vj/oVQ3FJFh
ZerMYMBEuGVrOnKIHVfF4WHJTfTSDu9uT+LzXCh3Xh64EtiPpWHYFsqHmFLuzBjadZBdIKjaXngU
C4kgy+nECdVb6xqDQ+Khm1hToLhitJOGnaILl0aemNtWcnvP31bAKtpUhryHuoQ0pQvfyxZfvfKM
fan+DQX27b35TLkvTqkNx3zRYwH0G2GwbaDx3Jp+Ba+F2v8gLCIxG8JqL8gPrYtZqXj5xWIOuLjB
bnReL9JUJSJtmEkyXI/SJAZCwe3BrCgu4TXQTuYSrMdSOib3Kqny6YGHJZqOiovcr0LFEdkQ1hrI
HYzCtOSl0yldfC52RWf1u9g2R0zvp31Iv/cJ12chn3t0EeGZI5uc2e5D/VoU3hMmqLzqIITryzSh
yYFRjToaRtafFR3tcmMIPdkcsYowTDQjSm9f5fXfGGf4uV0ZqgdIOGzH8Gyv6WlNk6NhIpbn7gSu
3trUf3rVi49w2ulX3dEMlCRg+ITZ93yhDtnotYfJ1XJ4LMhekKY9+RTI0b60YG+Zl+2qq5E4zcIo
AQ+Qyv2KVGQ8MP6XDUeej0opyDuaBvCZihzXCoCr9vzr9Ke6Sak29KIcPaEuBUdJrMfkOq8xSAQi
LVv02sT03I9VTgVZVw4CA7c08KtePLiumMdbt1BxH8sSscRPfRpIDPjygZXrugW8IJkQ405cgY3y
EVeYnaSe7Rn2d2KIHOgbGZuh6Fe1E4zikBu/w60ubmYAFhsJW9DTd/l9rUlTaDMPm0/SSR9uUtRB
VUpOM46H7AlcfjE2pNoxOSBkKIU+/8L4M1wzDTYD9NwI62HWsQLaOaa9Fpznnj64OYMdC/57aMnk
qLY/uV69tiss9edquG9EOREJIbPBoJWJ1tDqgOdE67cxyaEdQGPetI0oM/UAtfY3Y3ES3fBD+Gvh
I0r+vr8c1TCz6rpl+4CFWIe+W/lMlhmPh+BvPm3wBLn7X1tkF6/dtVYR2uSYtGotKuWBaGuWz/i8
8zkiG3olj/97QjN9Fldh8wS6yPWjBo287G9w4bXh5qKVVm+Bfa2pD8AvBPdOM2P3vX1ZoGXY1id3
rELqClrkfRyCjA5zquV+ZdmDp7F1mod+4xNaIPXstWRONn2v63LVh+xh/zFUa0p+rtKWO+/a8WYW
hxWVcZWAd1PMq21TxynoBps2GliwgRwLmGbuJF9PWXX9CK7UNWskIn9fUCa0DcviNDgC5WlHiGHO
WPFY5Kr2ovy4vO+hQxWMd5qI5/Bl4LfbYtolEidac8tED0xJHm5VB42/z46iY8SC9O8k9/BO+Oj5
47EhKQVNJITSh44Ea23DyeuqJ86d7fmVSE2FhIzYJT/T/wMvddBhFUFJJVIwEaKvudz8J39iJ7H+
QDKHFFjDvZxUpdeZbsFrB7dDPkMqgvKUO0Bxwe7khwXnHFg/jqugTGO292bQYDyDVbvDbS9u4ltt
2kxmWtlMmM3xjKfj46mnIdeNCKyF7rlrddMG5B7M30fMg63HPquQ/R7oRMVZTcLKeQLwIsNDxACo
ci1t5MBbE5b3cbicX5bv/4T8ELwLalMq7u5J4rCrhMWCC1vrOT8www1KOXQ/LWPHTeR47GlM25lU
vanvf6mpsLV2EoG8pf5vzLG4fKInx5AZc6aVrWjjTSIh8UQBI75pCbYYOfNGFYv5EkKeOZ6zzEpL
xgWfgSdVIG6tJVFuRzzGP6k8w5+f9RZBteh6bw0srmNziJ+U2wuu+He5/1bytR6lfWPSD1QmWUKG
l+CJT31wRnsOIMkEog/ULaL6XWzLrfxZ4D0dl/mmwmAojDY2TWBlaKNYVd2kjy0JFm6YqWo7Qd4z
53MbxXsvG6i9Y+7q1HaCabVTs5KPOzC841x+e+rlYrfNmUfN1iLbEXKmTBsdGGiYNaHZSd+XWJhf
F/tFYI99cZMe3eB5Qgho3b+6e/nNNe/5tNoXeLrhX+OJhxE3/3R5vvWhnpcdzlDRj1lo+lGn+jgw
8lYMjr6zqJ9E47vC5jrH2OBaOxwIIewiXRJCQLffkREYa9MJLCCyRAACHSyGrbnrKirZeiCruuQU
bO7U/pnD+8oKI5V0EJoSukLzsTACcElH2c3tGzcsb9tU86JBHM+lqGdQ+vRG0S9P2YDMhAFyYV0H
hm2vn1R7qODWgpQZYYAO8Sq3UQwjLY/yjd0mTFzVF834LKOxCUH7ofScIBLZo6fs6iBNIZ0RduSx
s6cuS9yuErX5AJlWuhbp+lZEpI/XBWuVt4ThcPp5hl1UkOffHsSKxCH/kvp+PH1ThUYyCIo04uiM
1Fgy0vQP0AIPDVgvDYnWxtbONV3z/xx53I+JzOO1wF1Qs9DBP+P96Uk+0Euc0BV9MvJpYQsX67sR
2jZM1gGx5a33ZPDBmwpWPA20pfXNuW2MyEVYCDxxdBUqgwZnHLAO5ig4Sui6Ltcsosp4n7XiRSqU
5L6TmFtxCJ10vFqWiRO3BoTGfO7BF9LD3lTZO0VUPME/DbnlmpSJZtpizo5Lc8pP0xJ7WRPE9+iE
CoTIEoIrEqgrKs0rHjC9sxfI0iKc88liVGcOcP6a/M09l5mv+XsrT2/RzLKjVJFVn4Kyad3HJhGW
qNOh0mmb4b+8kS4Y4Fh3QECnhpE+FgjabJdWXOHVQqXB66InmZ1iqieTmH+Q8Uqts+Pxzq1ju1od
creER99Vi0+D+2G0ECEzJNQuXTrCVA4s5ME7aeDtXN9mc4wMBTbw/6IT1PtyZKO+g/9u0wxeQpSP
ryf4pq2/O9NmU9ma5qab88tlvTsWtyxBjlrvxsMLTlva/ZTdxLMeMhkyGmHMdqbX92Asgyrqloe2
hnWYggv7cblf1XjUav5DOpHK1OQi+3O87/2B2oprmM2XJrQh8idSpcCOSEfQMAJ5Hku7bEdHQmpi
FgUV4K1BUOv0mgMm8vSRHl+6n7fpDW/XYE/Fyh70Ua/H0YzkkLDantu3PzGijPvdDES2krYFym6O
BS5lYlYugQ7yHU3O7XyM4dbbR9ORscUUNC0aZ0MEh2XHAIZr7XhXgHcyWIgocuubS7QbQ23qnccM
UNLdMZz1ox7g3zQBxkPc1WMWodajemh90HaDurN1CwAznYJA62KLnMDhvLXwV1wslRPUCNQQfysI
jDK/zk5n1Z7j+4FYS7rOoJVhg00VUinPS/mAw+QfMf3LJlaRYFXTIjgVlDLleJdsjHN3b5HXG/1h
amZQ1+5ktkEYcmZJ7ZNc0bPCiycauy+awaQXluPz9/HiUARfCiRsptHfb1oZcii4a53frz+m3Z05
6pxMQefBwPOyfO2GNXWk7Ze9JYEqTLbwQ+Ikbu1qxaqyjjY2xNJLmrQAxtxetgMEafo5hrn9wBuf
6K5G5W7SD9BRnR5NTfy4+CiscN91d88QEONwzD3PMoM2ZMHvzQCiL7y4wDswyVwN8CVMG/FY+2HH
6AE2V1OOWobWN4ivxS/0TwuLFFGOQ7H0cXAhawjBnwGTfbKKaKG29HyZ0v4SXhv0EsMFy3fpoRDK
wuvZsg6KTALXBi1cRaxXg55DFEnpjMkcHtrBpk7wDJ/WJdU54fhFTsmKmg9k5KznlYB0zKI31h1Q
MSdQafJRTHVlZiAxJ8miQn/dFVWwxc0bjbdibv6QNWvHbb1FDjHjN/By/9gL8HWBelkjyJ7XfQBL
kKXoYwEedD7RREN6VyHOSCP45RVlCdf7hlPjXwlDfgBPc8VP547IHCzIFnI8cG7LlBsUMbMMJJ7s
7h52jzmCyBjH2ZnvLUqwwqXbbI4S6G1oylFBumpXEHCrZQElrkYlgAEK6Tij3xqrdTUmPjMvEPYe
/pzvEX1K9bIF3D73yrd7zfsi+Oeg0WSlFIhRRLev5XdFSTQCkzSH6YuWRkxzZC135IzLSHrt4gtM
YFXR63Cn0Shwlz2WUlNICvhZiLrFuX30B6UO73iw++A/SBoMeXgH8HvpQs2PpvaGtaUfHachsviy
fKc0clFDn+qWSQnSNKL2EDurtUHiqaEBdwXb1zpDtXNe9SfWpRK0Dn/dCXgYSNIiLjdkwNuQF4kV
yrjPzOg8teluqd2dPta055wvHBV4Qc70LldDwaxMmDGjBJG/eHMmIj5TLaLyRkkZBUdLGSGlkumz
pFzXDdiLK4P0tz6cDJprV9jLyhx1Ep4vGEyYfrsB7eS8N2vjCyat2pzspsToA6HxHV3KImxYMPX3
dblrhZC/KPo7lU2zq79quEUwVDC2XCCKZUwiLwbvBDAc65AAlmxw1gC0bGiFNOCqiFXqS9OkVV4C
AAg6hWF0ZjcvviJhdAEdapVSop6o2/ITVM0+AlYgrDTsglRyWuQWQ3a1e4FzSNS74QuZB14dkkE9
pjcyh1yMzPoA3tUg3dmrNPUf8bYZy60JYnyiQK0UHrpPQozajpN58tUutQdJ8m1E84DJgv/oVLlH
LKigLD8asDU4weealR7cfrUGXIkpbvhenPJ9Lr+DYEYU+lvLNEN9SH1+S1FCBEbxPRApHcHb6eWS
ovJ1mrmBNghCMb28QCIOdus4pjoHcazePGjDZAqo1+m0tzIW8pBr9aJkE70GV4mfYqnXNF0Ihlf1
I0XQeW9uYtpcilRoJlUUcm671MFC7DoshNXUBZ/HQLvY+C3tBbJHS6A2kgOMVmzAzsDeLBbiev2N
ez5/SaBi4cyuWBuCrbbC9SmbsMX724dnYlKVDmqhMh4ssC0JqJgRaeKsrRFlM5rsszMXaEDDQVeK
kcvsCOQuvO1dyl13m2tuGTDMa3utMEvTw9zSi6O+WEhLIyWmXmK42ZPzgG+WWVlnUkOPt0NMx8kU
Gkw0sDhNoET8BcGZpFA0wPUlSAMxCS/PAhCVnfacs6BnOClMH4+hfSABJZvjbnwcNs2Fo3vOzc8P
MmDAbgN6V+/r+wI+RuoRBfII5Fp1Py9xH5OzZKEyA4PJqI5qGUxKQ6B8C+3THUokB6bWGTygHlIE
QAgN4cjDSz4qfL8YhA1NTDjkrwIUbKXcUMLsvGKxM0kzKwlqDiAdSu44x2Akumq+B3T+5M/M1hOc
7hRE/RH/w35kR/9N5ssbV1AUt/jF/OkuTvotYys4Oc3mm/goAtPvSOKugj4Yhy4FAvNxYhSfLnqX
wJsWFr1z0omL306lZTKlB7mx2sYQs14KzYtP03OxJgvixTGr/1ZDRMGHlaMi0bqx+2/mjvCloVsM
hw+YXf1/D7ZpS/uMdwQOWUlbE/SIjjJiCy5t1vAKT5S/bjTbbv0es4hmJNDFeNUZx3rR/E8c5xIA
wjnjiLIKbrqEkUEdcgrNX5bCflmyavPloEpsFy2e71M4l9PyEbBVDEf0PhHh6VnofMtBnKZOgxiE
L4viG1ynyMdkhLeJzwGG1B7HzWMz58GqPqwye4JMoW5Zrlic/4/k8KamugmBpuK2w/9QnSItLxUp
tbllkMDh+q0pe4+3OPwQeIrIxfLkHUOk7wCVMmJBPHH52Fl80XYElhriMRMQL2ql9pcLMjS2MFyK
LKOmmF1YBmT2FylpFL2CHD/zoys2LmHkKlf28kAuwKKGM/N218CEkfcDRetNNATF8gSYtFndeKKQ
0xEJDIbyAxrj0VLMAHedkUXhFT5DSW3ud6hGa0Z5ckx8CmbM4ra9MPK/Aft697QrG+qV4ptGJmnx
HlE+RWva8gxyfuKQgvrbIdaUfuJMg/Yu4AbxGpnzU3MgqrzE8ENUm64rH1PJWTYUaNzZG8WQi1yF
tMmONfxf4Xbo+o4No8hFLSBm03s3rLH5zc9T+WNKchIZ55tAvAukxIoV3d/bR2pHRj+I5Mvn1DKr
8YHIvUVV4wkwTVvBGJI9jroUv0ObdfrmH/smM5Jc/g7vQa8e4KyW0ZWslp/PwwwNCNJGnbUMtvbU
hselWi/BV2UQ08z1/49GrBTJ+6BI38Qy3ceERQCVqXGlUMGAUK666+TDdUtifNw3tnkIWgP2Euhi
M2lmWBm3CpCvQDsORw9nFW53ccObkrNX0rPEcyLcckL0ImRcZ60YiQ+jez7uSg2ioA2VmOKMGb30
Zxyllq8BD5fYmm1S0TEb1AbDYkRzfjXVdLjZsJkpk3RWZ8TRXIf2MtFzXs2o4leyYf990bJg9yYU
nB4ol6aAvBCSXBKjqehcVFTA2l0duLjOYHnFtzb7sxjALAXE9liETChTFFMXgCMDfRj8C4nJfMH7
+QO8pSJ4atNHjOYek9YF9Qi8Sd9frVbC+cN6+vAw4+8cSDouH+kE2pIvJJ5V5rYUbpGJn5DKv2Z2
uGWTymftDNe+ZKo3N5hBwYyR/MAg4W5gKpew1bA+lw9cYu7uLo12dcUtrxclK2y2cOTFJpfAnTjs
FLZKuPaXebzhd2BTWAxV7dv+kdnJV9q2Ugpe8F6+sIR+uP9WfSSIr0gyDtsXxNX8IVyRzYp/zN/I
3PXbh9pxidOIRUbAKKB587iwbAHT+nJqqF+fc/NYSHyjX67GQ72Mc73V/XzWdQcyV1Hvt2y7ZTLK
HisjlTH+Dx/2o6cTLDmepoIugAHdOQ4UEgb3ODFXE60ME3+4zpWwu3tg8DOu61zI+nzEG3kYmRUF
eeY/QLVcvCc2DtFTsLbGdvsl8hE7u7a2ceConQhLiu/NfTYPO73cAkVaykwm+CE7cacvE+F6ti/w
Y22foqFSGyd/NJTtyvPZjYg2MiJIOmW9tl1SYokw0bVSYf5F1uw8+CuqyGxH0hrXSJ49M54OyjhP
2w0zcnEnfMfSOqfL5sDggJ1y5R+nTwUhSuHAGfSoWyGrl5O7KG7YqVp69HnOXbnwgbGLqY7A9HuQ
4J3hvyXAIQYkex3DH2bd1ZB47UE6gUMR7aPt+UDrjOsldH1wPJpvlSwLzpmWxw1H1buXnZxQQi0D
S44BFaHBhqsnIMIJdM6/EWRm1fEIh5Dhleb9H7AZtlclu3206c9HC/Rr7WYUSLz8yyQfJLwhY7WT
CWnJEnmsgQE/DTTnsAkADw3fD86nvbu203MRmBAy+vnd3C04Z6Cyc2lRTYAhzBQNt/sVwqEapyXj
+k6rPp4FMnRmDLTexUf6ysEYv/71LhumnRe4iAhmicOg/nvMxcvDnTjzmSFsmDnK6MRY8VE7VK9A
sRCRlqhkGM06IpLYdlaUYEhvOjryw1F3Z9EMwUPGoEzFrJIgB/TJfbM8hMUdCDZ4W7w5XteeE05D
UoOdsXiSuMWrk0+VmtwihIp3+LTZxSRHZKCHxsmFbg+MQ+IHPMLbjELTHBNEa3hN0J2NAOKnbBiE
IXcgSgfJHtgnM/a1IbObUJAADOBzpQHxHOOu8NTRTkhzeW08zsBN1Tuij01folqHKv92AAAsNh9o
sOxA1wdeZUm4VRweNyC3oUS7vW/LG3WdL7RlKQIK4aD5H08wfM75sa8/AFlAfPy0lzBq9uMJz6YL
jCB/pARpPIMq/TO6bHAE//vSmwuG0kOKOeYuUVax+JsQHpOfjWzBRQZOuWAFDFEDRiKUClNGiCsQ
gVsYprLLRTWBl6v06HDDRbu4guwl9p/Fsj58vMpaOBVK0wGxDFsjuMaBiA9/Gj8YaLdRmUWrU1AN
PFV0EWz7R8IHN/bkdTPCvAmIhAseMaPyxf7pURrkxuIJtShQjbQFYdv/wcmKbQd1oqTxE9HS5cpZ
Nz8qv8K3yXmz63c816PakF3vSBbzSFsNNsCjVlVB0xr5bS0tbwk2VY1zOhBT8DATE29pD/PI0JCS
EQI8/kVVGGEYWtCVmN10UiDloPF+nRrBse/M9nq/0B25RYL0L9T1eGCtW8GOJcW/WzgvKSiZJpNV
Hz3bv1LF2PUDAiJ/2YfK3Y7II4OvDUw7dUgQOkZvjVR+C3cGF3PUhLHtsKLU9GHT0/3EiEZ79cwc
De292HmWH4zt1LMXCxpXt9jFF/PMwhwbZOIZt+yNu9soOR0US7JiTKAHGDZoDF4PBTgg9Cbbb8uy
GNMJPuW4rSSqsmC+SVih2ytvROTObktIi+4+rsAiQh+G/HnZRQYnSG3yuEWarXqPctkwAqJzhXYu
5mv2mYHE1luRhfokNIMvpYKRrH7Foo1SdBQN6QOKKfvWRtbFmU4N5f713gruGew5JNNoIGjzgTyN
NpmlJysdLx7nGdObKkrdvOsks8xXPjLJsyDxhBiUqpK1fu05hEC0E/FGqlHxienBcuF9As/XnbBq
qTJFDeuYLaNH+Ljp9+QXfhmuKTAdOIE63g22YdfLcbL4XIPYZhSGAtDboUPwBZaiyfXdRxH3TVD7
hxhupFk30G/NhGCwa8d9PrQWnislkV4339bRnG4JpCzHk4ji/l+IBRMfwsng3mhp3O8gZekxS9Xj
Z9B96q39Qr/JGAiBlVlVBKJj4z7ZtdKoFr+I+Mq68D2FhWRDBo0kYk2LN1T2clrV2vARU6pJkn/4
YctlXJzYcdz3BiHyA7PBdBTgbANYBsux0FJlwxlVS3lMJGQqMdJBzMNOmeCyWMvWvfg75vn9SM/A
fP7SKsPdmiDDODsvysdG6SevVLMp8EMQmVL+wnmttZ/OcIlT/+ds5Ggii6DPR6b/vvn0ftABGwRr
/dvYppkTHxNt1BQuVs8fDVyczMQY41dauyNSa+o0zOdtYrfK1CFCFZCxV80aRDGqTfzq7Hf6/Tas
eiR8koRVcefe3Hd2dTYtLEJowcVM431Xgxi19YEs1XsceWEh6KZY/IDDdxErP1TmMpwrb28VXqcd
OdFaFcNw+K9MmsTYdZi/izV50wz9hvjFmuacjPTiH5quUrSbtvoMQkO4lU8ggBu/E2daF8uRSgnl
5LTBWwJqwbg/zuV7bb0eQKkm0VjCuOtubMyqV577Ka9vh31gwRiaZgpgjtzFWKIXp4mOf2IZxBHG
SmnYCRa49Y3Dpta/6FoVH/lX8EQuPPyZ1vPk/c8t52vtFiNUDlecNTqr/WXJ6Uq6qFTg/WhKlOpf
GTVXeqNq63mZtBNPuQH7KaHEGT5u8fpykUE9JkiHvfyhvAN9cchIVR3vvjAVd8JdJnYjiVN1BcCK
K348TP/PJMEkGgAi30K+FB18KAav8VhOTRwQ9pEWYGxU78XThm6jBqx5slYx+EntZWTI5Uq0hCGm
c8PlGRtXFHLFzz1OKEcSI3Duo4qzahpLbEiYO/SF3o09ZMg+3UstBT6c6mpzGemLGomebO5dY68a
8108VXDpsh29ghv5xcMgps4flCQGLAH/n0/cE7QHw59DER4ZyhwXIZy+h0kixG8WabR3Vr2RPYBa
PlNimgWGij1w8VsUzVvge96CgR8Ksdai4ZknzccfOYPArIsf2PPSIPElyKmEL2QUywN4+fDnjfvu
z1ltfDIz/2ZR2r8TGLXUpZ/CFqzLJDGUFPFWEQ/5Scp8RsWbN6sitM1uumWEg3cON+86D9IaD8Im
zY7exLwKFX0EmKYH3HVU/RaXIgUU1CXDU8v3YXrr6fG24DWWOkY4lGdb+bDOAOLVt4Ze9jyypChU
KKXeQTHchnn/FzNF5PSU9qVs9XGi6KAdYJpUuxdfhUQGfeOIGSLpOPXvGig7ydkzcjym71qboFss
DF3q9oSmPcBuymAZKfnnFmnVlt9ZI+xvZOEoehIDIilaNcKPUqvjJsRwKKV7kZ536+rQfm4hZa8h
GK2WMMRfaztiAEXaWE3HzX0KAPXR7agWc/UH5N27zhqD9Lwk/l76g1xC8TjV/d9wAktG3b5Rn/ji
/CNsGs6+zk/wkClEq5Ap2cmhYuj8tPgMk0eDCQoYYH1Weobe69b4cZVoOpPES+0R14tYeHqLDzR1
plrTN4cz+cC90kRR212TjulSunRFZ+bhMVeYJwc2WuZs5/MD3zc+V/24IcYV2AAngNhZEFwGtPU/
FXGSrooTcfO2WS+YyB/SzsPkePCaTDMoeQ3wOKNOGrVqdeOCBiNEqUm7zQt7HJNzLQA00jO8XUoX
eWH+PnVPK56hH98r6u+7IK1kGyioR/Tsn/DxKMJoldJHk787AfImhmD2AsI2zgJPFDcsHAMuFnaH
cqv1pKaZGdP8RNxbnIlttfiF8uQPL8n5xXa5/6EWXPXHaYlDOSn91J7gIaTeTEb/t7qrsZaK+myy
Y/LJgd7BLrnuVGHVQW79eA0AOvoQ7uCE7E0fb2ekFy+qzFB1l2MLGpzHA5rzrsBuGtKoakLcyo2U
LwDiwTBS7s5nEIDqrw4lkf9RL3OfSZfVf38Z/b74Q3PVUUv6zHSVQaSVFPR3IER/S7W0gWNkvzMy
svo7Dh8dOwLBwEtVyJYQY326Al2j38JQ/HcdOVshDuwVIWNeiSdFYst48RCaBfaBYPSpK2TG0hZg
g1GR2dV0zkFsOVwuDarYmp9GZIeyc7BkREphN7gS4+vlroRENMlcovAjSQD3OO5laPvREXnCOccI
lWgJOIJLDlDZcR83TL+iqIMFqBJJM5rRUspeM9mNC8SoK8raHZb88XlxzaXfpqC78zAojuEhLZwd
HU8Qzx021LRSUZPzkvEba6zc2ihZOmmc2LWV1Crzy3yDt/MMyqnBZj/HUuCysW5syPKxIzdlv8YS
IOa3997+PdRYqfGaMRCKJ9wifeJqY28dAbJXsVPQPvQowl+cqb97rAvWycoIrDw/5quNdzVfRB8p
WGsRw2D2DBJYKBsNGWscPyO14kpKuJTlW0uXXnBYOBvBuDrCNuT/xr4H3Os1RDm+xuPLj6CNkGLV
dPsYK1WaTS9gObWU4nOFDbWu8/mBcFLXV9HxCIFqWTgZV6qTQT5KAGio0flM1MTMlDLUHjqwo6rV
/mKJkkecAFKDUfqnRjQVVLCXwBu+X7vay5RQK36o/ldXEiDjTkLmt5FFgk8xI5musreVYI39ydMc
1286nlrkiRkEr78Li0Y0TP4/HrfORCCI695akH33kbXYARy+RuI+r43OeFeqYvRjPVquYyj1BK1q
D2wRMAvEB/lKBtQ7F3o7dDcWLX3A2LBh7X7jYTxK7wVc0zS2D/L58reIgJ6O1b8NWPaoAtQnKt92
YpQqdnGxXRg0AqvUJHINj/jh19qgk85DBfSzhuzNg7y7LXSsiSHxifyI6o/zogLFjcUMISPneotn
DN9bM/MjySR8D4xXP7cIfGNQaVjqzst4dl9ZwVCGLDRg1wldJxXRLZ9A4UBSPM00oBdMs2PCcZl7
gO/x2TJMHv6hkfSQaIU9fqaQRSu7rEFowX5A5VL4wVQJ6fyp+Zuzx7Vgn9cx27yyAd7muw5xzCVc
MMS5MczDCAqqb13gfD2WriFEEceQmHAj2A+8s7XSqg0YIlYCQJKYocc8r+ECWb2m35m+apv6DHLg
gDkRDsGIsLH8/Uk6kWlbwbDMm82MJCtF0gxzFcd7tv9FfJrxg/2RdgdtYlnxMHldW6ZTKsGJoKF8
dTEqB0G1x62xnPmX13TWcVt7m55pbU0gXBvxitk1EaD7iwaJKAwn7HoG4KfLnN0Vr7y7W2YThlMT
S2issa0aU1ZGBk7pNneWBp0FZKbPRZaVF7qqX7Lykum8TiQXA4V6OJAk6gezcyQJJweni9ji5lfm
hchVkkLdbk8LlRC21Lcf6W/+RpO6+KastwS+GM2V9tqZr5iQE0Q+VGacVmcz0JYVTAeMfbsLptp2
DcmWdHpkHNDdo2Fzjpr7d0pnAJfD5GTjgsDAwYgJNL8uUT+3bZTJiq3f7bVmkOUPxIsJgY7h6iY5
I9Bi7QhAiqaZeAsFa6ICvDRCGrDLsNJOgs3sZ1m8VKACiheoD856Iy5kA+d5r/Ycr2bM3uWtbM14
1iWzx2WVvB+8LVuSbPMPolSd3phREHZpwfN7Ol3Gg3A7B3bhv7jWMrbrEy6AEwgzTdKIIMtctOUw
g0nbMcwh0734puihHIMItWBgvlzlu9GCWKoTZf63CE6C8yNqV/TNMI+xvtAA/5NQTHGn8zc05kNi
49sJ7e/Oje58RsXOErX70juFK6cbaWp+jgmEck5XDLgnJbEQiHFcECstc+N8biyOtydwLz2sMPfo
Ef3XqtJPBPsQ1vMuU8kZCwHdUogMfR8fbhMj5ByTYVl25UavxrseX6SC10MvrojSqfEt1CkRw4Sb
a55vc7DAuGIOBYJ31J+WOgzV5jjtOofkeiBVFIHcjTGOTtsFW84OkQXWhIeF3OqnS946aAgM1OyA
2McHZqHW4DuWgraSYyUqMCcwerhglc2YGpSddNnLJ+er3LXsCyLY0SIOK1E0NdwYuO4YZu1IAjfw
hy9f3EY5eTiwixcNSjgzbUYc4nZVlf57mFEiN66ddKP8jgKOVsyfaHTDc76dLU5aNg+7hRxi2/Cg
qb8LGptyiOQnTU0sLDCxTB07cZ3G4vrsTak8xgMzJaglgLbM4h/W5WgfVrnuxi6kEd6cXHJMlkjv
f5A/FICLDUgX7wIyJpgjnEtFpfYwa+gSXl5cqQ2L0KhMk6EgMkbc7b2LFqhF1JWzMO4UroAvI8R3
mxsTxi7Ngq7zBs1pbmHxWrtlCHKSej9ZcbauWSX7OK5MK0GIfxRSJFfRqD2TgIGhUSQigRzwMHkL
DVTD1F6p//3CIZyRvQSuhPubtVHquOPMTBnGhXfM2P9I71NbN2cE9ST9JmkE1nMCybCB7/WrcyRP
MyrE50NFpaPcZYDOP7y6ealfTBT3AcqpmdVJ36pWsBLiX94CG8inCQC+IR8J0NMq+ZB0Lp2/OKZS
wJwLG2E/uzXXIJGl/cmdReFflc4dOMU20ZAsm76eCLhqSF+lnHPolztOlofUqF3tU7zNc2UYOJIq
TeF3dIbgjBT31csdHPMy8YZzR018iGq1IbXPecyJ/Vj03xid1XkXYSEye2kgVwcga9oIlgfe13eY
0cIzHSRwe0wJobOQTop/A25SYBd1TqVPBY8Xff9r2HlyA+D72/EViLEaqKcefwaUGH1khEpneUPt
jGDFthkPFVyej4JXzQT4O0dm2x465UCybVuAkr1rwCKpWjD1iOpx6PF+Mt4vJ/oDMME9dWE48Wbe
xY5IcUc2pYzfGtzwlJHOaRjuicEj7BBA9M9wCsp2N3AjFSMdQpASMxRtUHaCtrvq+DQz8AzBvYoc
MOXGqsD8mkjE9tlZCIYCa6/ClMS5j3t4ARfLDB8rkudrAR5yKCppbISIJf6sguaiVH2udkZbrawl
0ixptoaqmMZ3Dd0ILO8lLJ2IyXEa53bfesU7qd2XOcKPwfnnb3t81jkQ1EmJSw7k9qJBJRgUbRMZ
1P5Jq+ERumrnPLGI6fTo8WuL1/RtfTD8qd5ryPVzALOXuaJNTT0JeFUXrnbmJ9ylr+Xmm5B9UH/u
erUoSt3Ki/bDfBXrzZzspdPbGtpnOzgxB5v8DWOM6pKo8HjUW7PnZmmbG7+2LNlknD8mxwxuDAEu
kGiWaw8RJ3IpdXOBGUo5AOPXm2NZO3M1zqrXnzOIk8gSCdncORtqsYEMUZHiNRlF2+zUnVeXTCn0
tTIBcte8rIi+UDLY2r9zMbDcE214oLt18vmLbEe49Kv+gkUg8b7aq+oFLc4g2DHICFzmVy2wA96z
8OB/uZHD2Zy9bQ9a+pQKZVAw1Z1Y18USV9vl/L+xMnlBwJuqc1FR77igNsSs82uLYy7A21xIUdLM
aSliGHairCbC3/yLKU2JB0t9gq1ctL+51TkHIk0wkDxSzOGzYloMkYNZ8oaWDSnpPjhyLHCA6e9j
XwGw9A5xsUAMejRqb8Frk7H5iVNjpDoxFdxb/TJT0XDyOmHsm69WUVJD/Lntcx81S3Hbuk/sJctW
e2W9M8Zl/2wcG647kLUJbshmtZ1cAGEubu8DbknEyq/cwtKx7yrXrjIpZcOmIIrYp2iDSjrg3gCQ
+b3fUmpFw+/5mNhjKNo3FBE99qa9s9Nbxzc2Pv/n/rvI4aUprVqvRVQtW1TH98xpVrAu+m62hibF
KUjULk/HKOlxKpzS4sDgJF6nXKbo2iHklGSHukTTILOIklZtElvbi6A2Cgh7oRegdVYPm1lGaI8K
WRiGYzM+u/uxWGxk2I6mUF/eFxPZ2u2QtXddy1KN2GUG1wt0UrN5cdnaJ83dbd/dP7ap6dwVgF/y
kKm5KpnWk2fcG/NiHF31MhpBorcri1zDRrdUPBO8QpEpHRowWRr/4BFYI1qQ/7KbbiYdNqEPJfQu
5r1+xj4dkomG2pqckMI2WuHs525iEVaE051JDeBEeVRn8F7dpuaK7Y4Yjwx2MwYVc2+B1a3ABoDL
gCXQmgkFrd2+1f/G2MM9dYXFwPSJqtQ2sZxdHWZpCCG/nZ2BLqYQFQq6QIhI2SUtJFEUazxrK9vq
ce9EqDUTC9/qWqZme8E4g1mRUhKKKWAS0CGRCY3oJe4SPjy2Npy/IJsqODYkiekLTu4HE37YAgGV
Eld1vtvGBmc5+WMs2EXsp4NTNsSNM9S1ML2VBHIcqJ+IR3031vt+gvbt5dxFSTBlCIbphwMMAazd
BggxW8xQMMza7ABK6EYe0SF2ouHqiZxOx6PcK8Th++a03x95pXvQNRAz2gm2mw7fsciDZ1nz61+j
SMXRUxsa9VolttQjaoutehj5zaSzujsNJsYcXoRH5uIPeBzBzmwEWjqq3fgIC3YqTzpAS/hzRbD7
whD6hqCW3Bz+HcMGdnDm+uebyw0wdAfIucL9zWVeQJc+1lQZrJO+2sobIG02BNiA1bf7vRpawEWe
EBkB6maZ+ObbXfGRFDtUUqnZdHi261V6+2mwMLcZAGQ1gcHTQvZnQKA4YEpR2KzsUy4fMwrpw9r0
jEq8aOcEXsSFNwvyciIU5RsJ9L5CdwLYeca8hbdDl3UTgG1oWpGvdxEUKiQHYDPTNQxQV9PLznWW
gq8O7IxcV3nKg/lOSxkOAwVEFxzLZzzFxRGMbfYl8vVW/WpzkaNSD+L4w5lNKlo+DZxYFqn+pH9+
E8vzAt30UNqnxwL7wz1BQIUHk00gXbDOQVYrIbIkHd+LImvHZfXoGNCCMJbkeOKdiiojJNpzA6kD
f1skYENDo27LgsLLNahgGmdMuZCOKqpKoymhLOeqcg+0I+IazIf7JFn/BBA5zwtUV9cidTSLdXJl
iw06CZrVlk3cmCHVT5xZjbGXlAozcJYzmMLwUEadeinvOmvdnrq96t/gq60fe/cG8VZQr4sMoVys
RlSgieSc2vRmEUw2qu7Vs/ZVIjGX36tbEusSo31LCfDCNtMN59NlRaJxYcn4x8u7g1V6BJTd5J/i
Vgf0f0Q+GHuoWKpYQ6y9Gz8pV7SaZYAiVkKvmRRhTyPxD85l5nNwmdGzSpz0UBanydLDpGB9VJps
siAeGwyXeDblb+CylcIyX2kZ8dY2qCzoozpkTHePy/GKstmfUTNiCo6wj/HkPJ3T+9oISOdkMy0Z
0OBdFag42mv4rRAPbz2+fHJFaYMjVt+X+aM6xOQ7IhtckqArPGwA+udWtN41JsxJ8Z1L1LXfzmOt
IWdwH2z1xaYgyo1If2BzoQycBLsZs8mPQJI1vwSvC9CicGJCDfbXxTDvx14lsR+nbZyoA4HEAsto
ndaxc36Atw/NREQJ5Wi/H6PIaUJXKy3XszWN7jL7OiViVfxgUQkAOqrMr3EzyjHxsWu79t7Fg2fE
OKpBRBZaDr+1LTOgckMBqjbvm/ZWZKJjw/C9NNOjI/fcG9TUmbwGWrsop/hzvwBTUxBxKoMe+nmP
CvZh0T68OB1jRSA78xb75DOZTd+l/KzRPABLR8aL8mKUICRtLoA6qkqyP84y03fMMZjZ4Nw1z+8q
X7BjGtlDrnRfzZ8UT37Y7P3d4bGz2/jCjG6tUB7Ot+QEyQaYE9CPSmEZNVXyCkyyV2X9iYxqaJLB
T9+vbaKGH8h9nXxKclvypC65wBXU3tPW9EUEURAVr59TSzqBlZPu4b9RotyUPD3WNK7LgUt15SmL
iPs9HLLtiZ1d2DOMmYm33IgWkA0hcPusFGdhCt9Qgow5B18nzM+SZgWC1CuNUSpsqHJn7wJ65ySl
7zOKFSBmkHNrAORKQR+hSKYC+zJ8FCrvEpFI4/qBuT1rlGpofnYBZ3n1DIs107rtx2UCYDhHfgQK
tWPtOFGrrYUllF8XZA3L1ziqLaM8uBbHlp/3IiaUmSnMavt54cVRa4JGYvN1Y78UFAIpDF0Lrghq
yPXsz5IprhZnJNjILTu+TOqFD3qEbQwVrOm8OYIfPDDIdBauc9YGCH6OIhV+plkzsg6pF1oV4sxz
yloLr0R/WToozhdoyZuAfmR+J82RpZ2XX1NoR/KzzeGKJi3MiZt1+f6HEbBoZxzcg7vyDiXkMkUL
nixY6dkwvbK05xJKbhTs7MvhVWPu2ZrfHQUgpSz9w8TESGRWetaG8b8krpwsCGkUG3KPhCerIaiz
o/cMHSC5dYFC33S2w9mD4S6m82RzGdo7tln4vXqvqWxh5rWsy1CwPXvEMj2KwnZhL4XTtCLQW0SX
/i5UoXByhAtVLUqJcL6hXGPbH3xuau3CNbhEdyv9A9Z8JMcx0VJkCvK42JkBs1o3CGWcXF+YIwWM
YFdL/Y6qc6vIxwC/LZZ83ASeB2VCApTsiDZg9hUfDr5rfz+eBxT5vPA1CU6enWNYFrgUvIug86SQ
FxnIyUPlzN+A+Ht0w4ailaEmGBCHrbi/ddA6Lqp6vSjuebqcvzydANzHvi7LLIJKgXujHR61/ZVU
eD1TJB2CftBJu/w2r4aE5ixRg7ZOJ9rYivB5aSXlxjviYDRGBJ0dJKqzdTSDMz/jhPI3g05Bs6fl
m9mDAnlqbuZ1FL5gZnt9hLZLnAHcfUFf78KuHT7E8WYkmPjWA5/Ob6gvB4YmLUfN00pOzwTk3eHv
rB6gBz6drcbQxMf7rKQsUKYeTaV0x2oFHz/GA+KAwqZzzxKFk3xUwINQeln6j13SmMCpgjotJU1p
oy2Hwa9lousEWYCkUYqkTQnPIxM6AdpojsMfJJ9fF/gbkxj1Nfe5siscbuv0KlYN1hmNMcFa0vuI
5MbV+YwUzJW4PvfwUEbk1N7dtPCZJLZqL4gr3C9agk+eNx36KEo9Jqv8Y+RjhktLvMq9tKEjrTBr
nWrXs+lAm3Yhm8BuId8hFSfgKUeF8Ua8LULP4uH5PfWk2NTaaCTeoM9gH3qloBcSICmZ4EsTED3U
Qoc/UJUM0h6xNJWXbtmFuyG8UjBy/8RmSw6nCQl3j/3jSWZrLUofSdBi0yzUUXDrFAR2DWryey1h
pOrfYI8uFgxZVqezBth8C35IxHSakz9mfPTrVl7Xddia4ctbZ+rrTpQg2up34ervSamWGyoKCmqZ
Bvm/SH4W9dVzKlflaIdaVLdTSN268RtA2hUvWFtfTswlANAuGlzzfiki7ZKo+LJ9XlqFAWAyMQ8L
8yGkBmTf7J+MvSzbumNXis/r7Gdbo9Bv3lLUa4zrZNYIFnhn3RDow2p6710KWWOhiHueKzBF+2UO
+gxYDFsHL+tG1KDNXkSS/Tv3Sipgt0QMNLJQsryhQe1DyIHbvyYxU0etXi0LcuoRJG4+9P2kMQFU
9UZZko4YNLSw0RqK5rPbDJC9Zi8niZN8NNI2/yn+5NaOAKlTbRbNJ6JVS48qsAWzlWzyqHIJAQXh
+dtVnV5WtJADyZhr1fwIm23z6PNHABGMJXxGGc8gT1+jWMqyFhewp+pLPS2TI+GYcw2DUoL6gYOG
nW5ugGMe6pYAzKoSFGUhew7ngUMZzpRkDe6qETWLVHOihhmLcNdJIagn5f3aThNYfTP37ebPgLer
WJ5ey1plGwbFjzWZyC0w9eUh/aMYPHqayWsLdVq14Pa6vruTjDfiivkXc7Z55wANeqW7PqEMp+OR
9EfN8lmSEjBSgt19q6iW8UruU4VjzX/dq4uzS/y9B2bmKWLDF+rl96t+R8o63GWTFHuYwrvtTdiH
XVpDPWZmyHI6tLr5bHzQF3AEoVd74bPLnn+EAAqjkx++yzd1oNIvvDbmUQdzVtSuPOD6nD+0UuG7
kzOhulDohBfsG0At7by8r4Bc3m/+KKYFGa3ekH1trIozGJBr+8G0IUrvNF2Ky+2vXmkmvhypC+yT
PH3TCVDYhphZiiat6tykQJkYUyVPwczYtt6OB2QPHz9pVw8f9je2waxdq60ti98QheNYEMMsJkPi
vMjvh0QEElsUyAlEkmZvuutHHvJxRZX0g1mtcMxMOFEAQXFuRpqik0WpP523TmDuvYwd9wcMYSnB
1IAyBake+TV8qxaMBGkJ8Dnxc4NPYV0A2x/fUrw7adx3xCLpkAkSCcHzA+yojOL4huU23SsPSyLM
fKxyzhtqq4Wkica+bVnDjB/6C9xIjmhlGcBCqz7vHwWCvSBCbzLQfhZNZJut6+6PI4DVModaSQiy
9GggQPdUQ0oGwvwSKoxM4F9j70d942KRWD6sMeLMhq25SKWE8KIJJ9mhXuUb9rTB3wlJpA1ZO+IB
jx+uVUeK82qVioo0NfU2afiL7nBKVHd+r2Dtm5WbghLgMMxXvDX/rzD6IyuM70BCDy6DVxHmbFN8
naUCVNoJ+BMxQ0aVjDpR0AjKYU/QFgQIAE2Y6RkyDFsxdNAF+fRRHVlLNRkMoxIVOTVty9Ni6hrf
mNu36wnOKAxi+scZa5G/bXcS9MHe0WseDZvyOSuBbYkE2lYIFUf20vav5Tn2ZYMghKaNywFxTV4p
dFSh/9m+DNugYMq5vje4S+DBzi71hjUEzpRAY780wD6KiaA33Q4aqwu42VKv5yzaJfdlewvQLlFs
EDxwlat0aZ2tyl8oCIbl/rMPQhZH4YHJwmXevxa82RvQkJ35O29gU2jpXnioaRXQXG9rqSdDjeph
tXi9Mwf/HIKSwMebniGzLe4aLX2q1iiWL95wfsSTCbHLPOeuN8sMmt8DmFk5kdQTz99AQ0CnXIL6
ExWf4pDwfFKY9i0UqaHTWpWGu0KLgXzsA3vpH4Rs5nha0t11bga8q69KGyLonRES2Hx80b5eCfDF
D9iQP5ghVbNg53I95SI/2hWNcNCZa9sC8JFK8agps6vAzEWEMvWoWj+xDltAYzI29kQxiQRvRLTd
CKTwAxsfWGySScjjws2xdzCJKlnkAXxclL8crKr5qB9zECNEQKla8ugpvksGiembAlEPmPK8gbuI
0DqePKXsrBmM3iDd84Po6FLZ2lYYOvuca5KpLwSTJlTekBTiO143y4VSLDXyAaJ1pUptgYsWSRqR
hYg4EPNgieVCRMbIi6Q1bo+/IDTQuBuMUDJ2wGNvqi3vDex/KkphQYXPxWu79Vo2+Rppv5fOhUKL
qotGENxH8mzyLMJx7vmETAdn0v3RhhbhSmUmLgK7804EP4qFYfgB7jRPaVk1UmUOR7xP6fGmO2ln
JU8prr8Vn+4enfbRU3+/DTph+27Cf88lVHGkhQow+5+G1KXvXTDdPOI1VdXiDAF3kt5hchZglrbJ
iT1LbOwY6kjPIo8MHeKTfvMQ1UZeOsbs6V3NM8NBU5xK+rWh9yoxQ5+PUVK84O66KhZfuN62cERp
VR162F4D0Bbk3gA3l6Iuti+MrW8wyJZaFrEDaHIlk9WgY8LYuQy0NutHrhPPTfCS6stHMCb5Kdtg
xsRmIeHqEhLK0CmS5a+WCs88PTykxJDZ2LWUEuROGBr20yX3FKDZju5oZ0sBfU1DyP58JyuEx7DT
/Ej3TLVwd2d8G0DGe8nO0s5o6ad5c3mot3gTcxBpUpPiKwJ+dwqdg+pYmbBI+h2xmqs8zn8fK2FF
8cn8QZ/47ayzIWR2QHBh1PISmoGhmp06np5n5uhUwOVjlf18DN2EBr2ggz2kLrnGM/5TJQ2viQHQ
hhqVbrY43lv8jYybkqa3IKsnyYG/eRIqoDmYa4o1QtsPwQrYcz0YObxoUjeDPgS+K2eUT+HvA7ZR
9zrpLfT7WdJ+nSfc0uuKPFvAsDawwav3YCw6bzu5F2FlqfktVE8FDsHtWmm8CGS/cQaXXaSSUSkR
gFN4oxsqNhIaNPqDObQaefX5OdsOvSRbdm/7n05m3R7TTq3nCFbAi3mi0IChWfouRcXi0uoHZT0R
igMTqz8mLAZibDDwHJkMnJzXl8op8AwoeQwGgEMCjuKMobuOPq/FbAfrkDvMMkv30O/9JauZJ2gd
LfD+OqC6jxvs3QOwznUu9jm70s3n4GUIsHHOzEqgu0gla9RDnsjRQgiQ+u8EjiMn36+KEonqyrKG
SsB6M1nC8i55sb+jd5eoyppjK49DUpnR2bg9pl8LyR7yjAZNFI0KOz5Rza4GZZ79dMPSezRUAZvR
FMuwXnMp7JNKgVLwQnsymQ4rAiHujHXoHUBRo/5CRgomtr/4WdHxOPwKNw7Ql51iQC3dJaQGRBrT
TGnBD8JaNi8ImfaJkg6JgpsdOjgs/0k/I9GBAx6RQN/HglDU28jT6tGYrISTccrSA2YUrJApgFnv
+pAO8/KzFR90STPQsr/AJiUjgtzHxFsmKYkBYCkAXGA6MmRMIvwLKE2vft3c9CtYPw0Hr11hsjJj
UIOlMcS/SK3l4Ii1FX2Qq8p7Y2V14+Hp6YvCbaHp8WKGjU++mJzbw7KR6Im4IE1oTOSMb6FHWUzr
yVYfV9Yn3t7f1yyK1q0+s/oCTs/EniOANKH3XKhxkVX6bFZcPBcE1f5HqPUMxzqRl35YLx/6n209
12ZBhOew/fdb+p1HFkSDfdz9y5Y02z2lRnBz0FKqp+srcwhEqfCwI4GU2OHuNwOHh24zvZMC0XHN
Tsy1WHnOs3+XsAarLa0rT0dh+KBb+DtoMkWurLl7dWQ9o6mFwN2cdKKOOY0itEVFWZdtqO7k4pSn
41M1IjC1M7uLK+HhoTQGnUNRlBpUN+gPQn9W1dGpDV+ufRfeDLuP58ytbaX8JqfoT5qJQf3pQOtV
2Bcf2shvNT12V5o8g3QMWH7fzM/tawaOGaIdan2oXXmKEm/DnD9rV0JT4P7G3jUvUQJbJ3AkS2sj
eNz1Vx1kpaVBdvf67X1KbcJ8sT2ppsfANbYbtilNFramfk2PrHraRuZVXfbbkN/se9Q9P/mLwUju
F0v0MX3/5XipDN4OdL+l9DDKc6x1OfL4pcCuliXBI4JFpbSmv0bw7/qtGhHbXwGkFlSbA4EV2euS
zNSU3RnsDc2SCWgknKRMRn7Or5B0NCK05S5VSQZBIdwcZe2sL+62XizMgtc+VZQwv30bxxjr6Wh8
l3Gll8LxMKbafq2i+plFkvGfTqqOx6xUbhYL5pN4doV0HjzLC8GjdtIBVbjVzjy9pfvYJdMambtI
hhuHC6VrS71/EQ0lCsBc7+FcnQgcL9Tgcp4zB1VYCTawnZgRBggmPSAj6ZeWnac0yJ/b2yyquMyC
WEE/Np3rvrRfKDGaNOUQaJBRAPjD5tR31PHAFq9JzR4scCZuS2YWg4HBdKmYUt79wFnHVw4OSE46
SFiHfgfVqlCjWuLc5uciUD9blIAPfCzEYavPrG+XTGEkXTcrwDxwNp7Cqjed3jyl57JVU1bllhA4
UCRbJpq9j9vg6rdU98j4fuRs17+hj/6CUC9soC8XqLAkwVEzJYpj2M0ilRsm4we4WwPIhjVYSMmu
aksqhq6OhOS9ojsjkwx+CPaWLXxnsGDPs2RFJyz+cmmgpyxm2nIRzMOx1aa+slgIzqyDQsQwY+LB
JLkWF8ECnaVY2vGCuIgNx/oKmdf4fSr0BYCFkIdlGaaDvE2mnqd2eI48fCC636Lb099dASWEWqvp
bOQy1//XWw3PeOuiF0t6KsttyGuaDDi/yhEEZ9ZFKlKrAyJALz0/dfE6naUw2Q1SWnsVDHayVmK9
5StlcQJ2YIP0XaHrJCw83+yCE2+gRqI5HJ7W91o3FLae2mtDAQHpodD0YNxPrY9MA+JPvcGntyZI
ZEF2U5czXI+6ba6svR/gbsdsMjOuT8ONMb5cWIBJDr78KGnxZBCGpqwtlrPiFKLPolQC5CTwhfqx
QYrXEqhdJMx8ynjcKGTKEOLvwC9A9d0Os0HIVhs0NEbYrQ1B5f1UoX0GPpuj8ImM84HiuWHKeCWU
sjDVVqkFwtI4+RIb4chKlozxH4xIqGfg3GXH/0cTH6xN1/zCkGxthsewMweWbRe0GXguOa6oZu8l
ZKwC9BjMaKjOPcrwpxVF7YbsowA0NB9uzJVBB/Xs2EtnshW2QtAf/z9zX3KYVGWRCpp6TNCJMOqU
XJEWGZ4dnTjFrpTd84e2ZOC8CYAU3Rz6SJXEnA+zMEvOxcj3gjz44SSUwtfWWO2ECZ9v6YdU0RkO
ikdEoeZrUuoZfUG7FsbfRoDhl9OE7D/jwk3LsM/jUrTdToxn3zsHIcMy6zXnjJtn7cD3FTY4yPYu
r5kPXJsaDE5dTqfoZmqgCYF63tEX4PW+i8Ik4nneKduVmfKe9fvfeXSC4tIGyQeAkvdPuPzQ2rHL
XgE/AbWuGjMpS7CU/LU682y0vKRcJLWKxZY3QMTOQKgasGiFI7pOja/x2Pim7lOKCEBl117TK99C
minQ/gl9X4SWbnZpeWNY7z1gIMv6FOK5sY8nlD8Z/kU+w65MhD0vAa9GM/Eeg1H3BDYIzYrfBuDw
jtnGuMOPiZCr088JK5Vz9Aw0D7BKOGC3ln8fp81U0mfSe0vnGSeR+YRNmZtoV0QS8GhUIMdrZ872
U+riqUjmCEA0jpTqsM6frivog6JhyfxWbDTlhdsNa07OrSyZw2OI8SGTdg84qM2XQOrmWiJ6FXX8
GpM9OR5Sl22l99hQuCBcE4rfEz8ddL3xUjEyeqCbpAGyLWEbg+8rxhQxsVQaPY6KYbngfxfI0Q+k
gt6gic+RH6nf2DWkzmIkwjl/SWTTlw3yTRVHuOM24O6iP+9TIC2DP8ikuqnrbvI4L5QM//7hkG4B
sv/nB+YseAIByIVPf7SBy8Gr+9hhfUMiImgaEQHnJEpgUhiuIlVyqggQsE1OgJz9joMidcoz3Qr3
ZMxYf6dPkXSoTRCbMd9dw6XKx+Mq5HvFboqg9VJK3+7SRLSQ/O7/E8BP9gVSdZFjgTqMeON/Cm17
W/mN8nmaL2PE+rrUJL/jjKrXZUAtxddXuivd36vnCx5eI+R6brzzntubuOp8p1b0z/fCS8KY2MNq
xFW8YPypuAwyQGGfZ/FGgXkm8GslYNZ60OLjfkJK0caHTpIkkWLRlbRFi1XiFe86dQfMY05p6g+A
0ppAmzN8jj3TLqN68lixU1TBQA5W0Oal1e9GvpKYB5Yb+6k47CR0A4hVW1v5XChDiQ++bkP3oKqa
dK6/09XwRlgcs0RYl+6BPfpymsMu/xoklR+UvgQUb/6garF6/R9Fei7oI7vbCZ2MW9D/ZOLcFZl5
U3Z99hEyix6X9T3TgHvFoQMMxGbNoyCKgwf1xeTJ63c+PVWIaRh1BVP8AfiOjU5xMYNMJc3/CgW3
cb6m7SNutGTwsboStdiGZ7arTvXdeuahotszUKwvDrAIQcpQDkSjE8QwQlbIiksip9MyCyhgu4w+
KhYBf7GqmtWkeD7dh6lTupONzqsmxGd+7d+caISVQzTkRcJWAkj+SpebHJsCQd7KU35pvIGuZHhY
o6AOlo5peZim3Q1ih6PvU0AoN0qOc+gI9XscYcmGJ4LWwfA4W/f2yb3MqFG2Lu4cLx8MctAkv14Z
ps8F3LILAlPzTKXVz7Gvc62nejqnirHpQG1Vz99pF7OkT5Jx0cdeLtQdYwECudnD+GmOq5qij/+o
7z10i9r1WG+WT3UcwdK7qkRW0Oy+V9akbaCVisr1xCCaRSvcT6QFWcSpocnrstl43cCozynwUhBS
yErElv/bywL4jZ0tEJbCuSDfhjl3ExIAvArPYyBY4AJdmXnYk1NUzSdv9K3n23HOGCAxRPrFr8WL
SBBYyIPDcG3z19wjgvTGIfFxsIFaqMggTC/yTNWPBjuJsYEyVelKje+Fvlf6m5k7yAZMAnfASDVQ
SJ2TzYuVzfOWLyD7iXJ8vvB25jC0mWQWixAKNxztdCv+qgWf9bXHAU81hQ6OS5/rx+wmEnckeYQ1
17F3xEpzOiuxQ/La7cGnU4Tl9Mgs+C+aLj977dELmPvTW/0OvndOR/VgQ5jo93xazyF4YJ20bjxo
bxg/td7Nvds88oZSegHAFC5KhCFkRLzhXguYeCJEvpjx8Vf8kKBXx3nRJNcCW84iL2t7mfr6oI5h
j7b5oWYlEQu8kAe6laZhJV5Pl6Dn0MXbjaVKunTJ7QKhMuYFtQu44jELl2BU0IJwOGRrdXpmEiK5
35VxT9fpTbvN9y1IGnrqjcrRYUULjAPyg93JgX66gMZdRX1XGeaZvdKgGpL0KjbgV4D2+S8DqVjs
KT/X/Ni4TKzVh7CfhdE9KYJvtjLoAen/W8DXn28J+GihIi41U2rjUVmonQ2w02iHm0uqu7352m7w
JTEpLpR/TkyshMT6vecf341KZSUnNk7Kgyc0SCDzRGxkmkRdzix+Y26z0m4Y09kqj4xIxqfcmE0m
CUmanPFtT17ciZnwgJbWINREfIAnZhUBOKm0Fv+Tmf6+oKDAbdtLLuUVvv0Mlma2u5uyrXkbF5Vr
vzPCLm0Z4rP3qZKCDG+pRfGOWmSgGEYh0a+15F43t01GZB9tZcfzC0uUNE+wBrtd1/h6MD4saTz1
Vnqko+dMYx1jt73ZAf42UQw2gAkZe/CDO5e2YM5YGaKrtEw//x/8Bpc+OHH8DEFsLVxaiw+Gvmxy
eFtv+aEv0oqzAzfWgsWcTxhuWIY05d8qNFhtEgWKmjg4ijyHxU2qJUzJRjvg4Zha+tv28FMkFaf7
TCMJd1rf8YvIZvK3yFfuxdcEtgnSBaP5JDiqJTi3SbomZeentX9j4up4CUTovQm/aQ4G+vNOKnw3
puNxKRHkaYXe9lkVDzTCozvnwz9cRVi8+sUBiuBMeqAw2Oz7QoeAcvR3TU8NtfseW073efcGlFt4
m131kaQgK1eAeJpyyq/vPFUe+yzaV2HIDbN+/M17VhcAh2dU3gWcgvcSjkovTUVr4hsw6x1hzzi2
38MxHvrZl4naCrhZpVDe1VoiK62aTUg0eaq4WKs5Wq27sXtI0JS1NWFSzpTXiw3gl9tRcu4fCoQG
ec/GIedDYv+wTkLZCagI3lvQWO17d6YkekZrrq+2v9ErzS4n2Wx/Y6TGxNJai7AnfpUgJKLK7lxR
59vFwXtRrK2rbPYldu31PA4GuD+RZhA1+hoV6adxdSh158BEYx5oJbRGSKmtep9kRaQFsBE/nqfZ
jhPQ1DCXWNWbxQvZCBKG74ZcqNTNjOGOtxKf/L/Wtrn/QJtVvGL2Ypyr3pu1eDmcdWJo6uwaCnnS
dAJZLXEa4cGykQL+TERdTYSfRW/fY0jqLe2AbWCm2PJIWzky32Mzb4D6Sa4ztEVzxNTRL8nuoYIm
uMo5Qh2fYPgzgLp7RVjdqVb1uxrzXK8fYitDnvdDoGi+XiIsGR/RkIpfdKwhGjjn08Zgyyip5/r4
HWmsPVD86Lq2MGho8yKcUTJrF2JV0lJhfU9QnaIhwN+z6Cykp+EPv5/VKPtnmaaloUk2fQD9RaDk
qZWCN2aoAYiN7r4q8ViJPUWQMK7QcnxS2MFs0wK1eRaTJYA8Rh9AbwFWfsE7fXZT3Zfe7Pcm+PA8
v+KDLLn8uqqo6gyez+6AUov7iJMMvs3wsSCFS2BLyw73PbBSBWu+4kKe2266UiZsFPsgV4W8/SJz
EYpoLNotH/snw9oSrGeADSGMJrteVcTBMVHX6NLQuWTTKoAk+Yy3wOL9wS1p2AEcUGD6aIjVwDTf
YiSMrVA0l1X6mDPsrs7RNJnA/VukCgGgKvRULZsa0zrpyVN1lmbWcNNKsePHGuXi/2K1okcI0xT9
bCVXcKLJVre2bQIQVjGV6kq9S2i+qi3vDEwvwPIcOCgyuGF+G2kwT+bROJdOzP8KsgRjRnXXAPfK
xIaqMjLyCuuHiuZOSU220LJS3ieBBB6wNTH8Wcgg0fAg7aCOGGd5XMSIAWMtssxuQlYMaMHf/r/Z
ue/teELGl6Z/JjUCxFLdGy6HR9xkalg0hd8S2qTc9LYJInpdKE1+6d7gng2KReijXDAvQj1/4Umj
UyzN2eJ3GIzIGEpBzKoGoWxCYk5+MyL0TTj9a+cPucBs8uVegqtG2B+hYTvbOBz4grp1t4MY9WP2
78EztccGq2NLKaILzWQ+3upl1p8LhbUOhWJoKuyYTD+T54KUEEqMsJt3AnNqW1+uKt5oud3sGSPZ
+22ZyiCgMdOelLOGM4Iwn3BC3sRsjZTmpXbxbCx/yYOmfyQ9X2nDcwRihPWYSHKQQnepiCx+XyZS
0yhFdsftbLbxNnUAF+NFkqFIYU7F1SKlHA21TJAzIPvPMw0Yj5B6cJLBtaZ3zMBuWVS91fGOxnBd
orNLNJD5rC1AN2TAf+/+zCQpSMop070W1xP4xHxsG1/KwJJqIgSwa6mRKurptQHXwVDkQsHENk23
LXEFDm+pYVItwrOsNwqd2C/Qa3VCrxeWvLmyYw/HmnT9Z8gjaBgeT+z2OVtwzzMArQSIqg55ZEmt
X+Dy/pfUcyKcGYI1WU6rP96b9YBnsgu8ePHdfnsxdeTVWnKAP5jctdzGYNAPZ5n29XRHpsnNRfqR
ukkv6WS2abPBXgP255BcRcHflI0HCBFcMOtYgwYIKGUx/ImCKIF8L03m6RNO9LOUuoLYaXP9O6aD
5GJrFdCP72Z8Yiv25hoKosmMM898QTvfvyURrz9jDbAD2p2Reh+Kr9rWASNMNTMJJnxVgTAOzyTr
1ilkJuv+2huTNPh5hZ24kOkXx7F3MWZYgwINi4bPTm+gukmT7IwM7l+thDx5ZVgny7DU1iTOzl5W
//OnOlXaAwBND3XLgRXnLfoEqXrDHikRx8THoR8Cvz/++d3RkoTkhdcxl+2FlBx9y2e5vvzeplX8
m1I5nOkKW3r2vtmKmmyMTaRSXVb1Y/IiGY52NP+u8jmPWPlnaCl9f2Ug3Gx82R3P6JGSvPyGMci0
CbvSH29p0WQD2ecqyNjbxSWkY9CTJnjwMFeWhG1ObbaUu3zHQ0kbKT7Ugfh4nbcTgvoA50IWjpTL
KsmuiPQSjjh2Keql3GLU2G3Sz4LgDyryHTq02qkMElDWhZ8UQW2R/tQ0wkN2z3u2aQytEh5jV3Xm
GriT4IioEubyvLhU3bZJe9+CT0qKIuQ6h0uzA0RySJCGz+rs7O2zFQjkNSuZNrdfkMxWL1qFeDRa
SNcivmrYD0uMqTFSpO82LnpkxdYmWkMlhrOFnM+eJC2hgIQgbqyHYcMygzwh4/vnh7FxmOqebeow
W4ova6fnAJfUKwV5xocMF5EXHAgIRLL0/7k2v/ZAuepl5Vv7qMgvMt39DqJBk2QyMoeR77KvUk1I
rJWoEucPn6lzLuXXAnVoPEQ/DvEPN1czWCVZSfJz+d6iDUeEudmNfpa5VZBxcuhszVyIcTIqtFSu
4yyV7FBApOid5fjr+vTEuRZi9aOhkxyIWaIEB6xBp4UPi0Lz3ZxkTNY3lyGy0GHtfC06PiX9dOa9
o80gW2LUHkHW/E2aqxkmBveXRKOFo+L5zK6FPp3Sil+pz0tfVeAGnCabW9YKmTpBjduG9Qhp2U5j
M6qJbITaVQTeYgwHqt539Lp88PZ0t49b1kBj09pJ3lQlckI+QvQHsvn6xc7RsjZGvw3k2i5hbo0w
T4BGvcVBa9tL0zh6yawEZZvT1ZoiztV5aeQxsGHX+Z9JDKPCx0i6fG7yPzhpHx1vc/E7xF0yWU/Z
QMeLNzyEjMJBc3qrTALjddlmgqSwVSx5aP3bayLb3Qyec8pzaOAf8AiFIANqmQyzqMra0V1cIqFT
rvSGvlnE9pzCXTXbgiVHX+S7yGEfqDdXeUD5bO5ZJSH6Gy1NiheWbnqTwjoWTuXYv9mjM49sU3w7
T2Or8ASFTP+22tPZoLmnhixE6nvXliDa4jFA/wjl4fdkinRym3BwSWN1e55l1Zp9M0r8KxENRnPi
cBNTJ5UOW/v2sVKj5RnebxeKjgzyBa1Td6ALGiAW9jbl0zw+oe0a7q+LboBoGLm1zVyVSqgbhzM1
zjd3DrN47Ddx5WYbpchms1U8ZKze1JfPW6iWuuYFPXbIcJbPV5ibaH7Jl+7FL57tysFOhZgwAIRw
uWoOMdsvJt+KDJlk9s69nZ/WV4yffYWzBUX/Rhnt4IIVEyY+Cijscm/LIg46TIrSpchgLKgeVQkg
MvgdPaLj+LWNuq4bdS2qdx2EGKhdM9Rr6GXnYAC7Mp7BHORKvrtTz4dxrfIoDDLkjiUHxLECazTu
N91MZlFH2Ki2mlsoGkDoNdHf5ISYGtaomYRMk3ny70Y9S95OagUucMkZ7IsMtSeIAeYSc5TGBrvi
hpNEBfhnYh0Oc5y6O0p0lO7zECU0hE0aPZHB/lXs6efU0pmJuWHpvZRbYIMv3rXeP9EzN9goFcEP
lNBDBzV7wLHg4rC7ewFZvF8eNfM8F2Q8/HIlQwNkotapDps+WyRd4bqDv+C/2HkKBpe6DD0+OyJ3
socoyhV0WOfWRt5rDwBGuRXvtxHjtM0pGCa9rK17W6w+RF+Vm/Od8uziIc2VDbcJD+6hgcDOvnXf
5mEC5H2pIinxV0UjxG5xDtEKQ8nKZYKiEx+RoUsCjPCS7SjAjWEA3LBeg6bbajuDUZzCzWsHBmHF
XkYfK67XNzgakfmFwhWH84hAyC+hDNbtfPEWeV7i847zGR4zfYkRXYEXn3ZyRrmoPo7zKiqf1K8k
PsqUbCQmycqbHvkIKMHdRSg7kPRMlQmXQrp8bliCXrKSxJljgCO83ryZ95bD79HmsdLFLX0218UR
EEC0H/zswaZkTS+s0S8pw8PF18I131bxGDqTX776dId8GX4iqUwUNg4+RubY933mWoT+W7fhRwNH
xZ+8XRKVP0cG+qbuR5gjVgiYOtAQ/+sXoZ8WswpduH8NiyVN3CN8UrGkd/TtBCoh9skfiFcWGPZu
AhLBx2x8bwHjJ863IgE/eCygOQAv1krwmzfqnZd++yFMWyvoyQ6o7JQ2LDjr5fwTDT+mVBFTBh98
PiRZsRhOFrjiRpDGCwJTwLeW27iPfO/Ru+xz5YllzpfVw9Z+QVdVgAi+/l60GGX9ZyC0hyL6wc1l
PeLROGgNcLEVhoKUAsqPWI48UsAR6iY0kASGJ+C2oTJQ4OTt3vIuVYn4zBybauBceMwhrRPjv5XJ
uulO6Gcae7BEXakzYtFapRJgKoas1kdWjOpSr4ZlzPY3B5XFiHqGXkxrseNsjQXx3BF+ofGUOYmr
1tlfk1IGFTKq+KKcVBj2LhZ9t0PaoQZSUvOnOf7V70mmczYHuTB/Q4G28+6aVk7sf+nRhnaUHsiY
1yRQjG0yE3tv6lymKCtRBGfEGIKcFOj8KWslyIF92zc8VFnz3lRMvDjzeILJB9Mkpf9tamit8d6C
EtxdbndunxDsInkWGzt+76A/iNcKdnrS0ZC0wx3PXjCd82n9r94JBSm63iLkJP1I+ZlEYdVsg0+1
xHXi/puwuc/ilwRcxG/nB8zz/O935YOD3D25wvO2Y3AztCJDSQ4b8T1fpmDMRQCtRUWRScaJjkPT
43AAPD2kw7/IaSDqrsUBip4IwtbNLi6LQ7IxHJiNjPyt01OidX0qF3WNk4Aoh4dkf/5tzerrv2pd
XfLEauJsOvFlqgIu0N5x+FLby1dSgULNWwMjUAx8s01/osMwUHGUiCetUygXGJ2pPzVcwPPMnv4E
qhlYq0uhm2BH03ofKqyy50zM2HFUlB3iic9h2Cue39m2A3+1Xnlg//zetl/O1uvtzyA6DCgFYrsq
QNVsZ7LgwWvizLj0+m0FVwg8VzmvLla6M+39tIU+fukXt4GhXJLqKGK8ON0rwTgpIMEIT38ekDYd
ocafHqAxuNNhItl7h1rSAgM2xrJ/lDeSNH235pbaPmZVawcXRsUIZ+Ig+c4gYpGXJ/0h7olyVJ4e
+tFXXzO2aEzRHhhTCUvBP4NFrwvvWgRR2eA7imz+fukSvmHtuch3tETFDQVURAy6gNyHJN5cGj9N
RuFFzwDTjzL/BAbUghPDn6ZNDkrYoMsHhyM5dm0IG86NW8GpvzJ501wPfzNtuTs4tYwqhYJ2I7O2
28EXEma+kRxO1/42RIWLdAa0+jxMQODZELVUsgRsFrvnJBqq67yiQDevLSe3akTPGs+1ea7/Ovb1
Szly4yocSTMXQpj1xPgghHfYYBSPhbO8UZPynFJkbdAddSwYNL02O0TcSqD293VjfI6e6u2sjPT5
6CpV8lG81cYbb4nrvEa3McUkNMP0o4TPzTcHwjc03aA8C+/Y+W5+Ow6A0tI+nQOP6TYqs2Xnqynz
wjUbFAOOOpMOzM7ojqNl5CmzCzcSHQ/b8omMYpfaiRmwlR+RN7lRwTzvI/iQzk+V/EwlXwEw7EHG
2wFWuyfqC14XjRxPrK74wRIvkeM9ReDjPXwVmiKHIWPnXs9Fvm7q73JO5nTrEkLl1FwuWhKhVkhx
XLpcrFj7FoH1urvY+9ZQlaKnplVozfHmPK/Tmt3HO5wZ9kS4WsH0Epf914/uwQdwIzkcLmKIFWN4
GxQ2zC0fw27W9iklN1XK37WdI3KT49YdH0pKyl8Ix3xV87U9hgioFRoqVzbthiQXO8TNVwvzNZk5
0v/o4sY4q4JqmqHTkKicr8XMBi1gLQUW6c03w7iSQqSmWRArm0t54hC6Ywff910u1L0S4j8anSOr
uENzIJjz5rdamRLG1vCGaMvcNw0HKkBI4xhEESRWQAy8oJMPsX2IPfx7wdzyudVfNwx6201mAezN
58sQzVDIipk48Mi9xTVJePRWmNK294q6BflzETDXdhCU6QUxj3aTanzgB7F8jIEgJcaGdmHno+BR
sYaVVF7FXa2UmaRcHJC5yIJI1FvUAgBM6f5KBCxvUv5us/QZXKEoopI3ylNeN2MsYh9ZTJWdCxfL
oJwj+2YR89XoSukPn0yE6mbpItvpmunYW7rADW8zFlkWA1OftES6c+if2RwKGTis30YsVGFUK+rM
rji2QdpLpPVy9VKZ9mJ6PeovCJsHGOztr0uCyzAEuBhWj7nvWL9Kb22SyZYTyy/KzmHp3kIhz18n
4JyW0j4sjTYvrU6+4NkcdheVFOGnSRqC+8nXXg2aZIoRlnLZbj8VH8MKVBzZAcet02pvHYD68ONC
ZcibtuD647DSC/XO7qxrfN1l7AQb7nKQMNTUwXqY2rr+oTgOz5Piu6sps+sqRU3RIDeWNSfd1JoQ
YT6IV9foUu0JapXxf80h6FtZAchD7PuYRxzuA7Bi6t9SvJ8WU45GDRy+6rxg+bVaopTenSi76rZ4
E9kWZqm67ZKrGtYR6wFubkOn6hdo6Vv5NtMrjevFySibelqBwfTNYXmtDWlzn0wFKVM1mfCDMYzI
Mj/gUAGPV2SLcT2VS6siyhT5NAtu5Itdv/mI46PbJoFTekDCgw4WLqJGaQdoVb4oZvMAnxg+zm3f
WujVjBcy7SDpajXwrc/PoCzAO1BB148pQdmph5/dlshLzYZ1UL8TlNJagWSxiuu4Ytqv6UJPlGHF
McPwyaPTIG+DM0Herz3vTDKlZUPeVw4mag4a5md8caIPgtdI7oqtQqAVwTu+8c6iOL+ZjcUixWs9
gdgLCGWYz3iljeb3CNEdXiTtuqx53KnDn3Nx1vVUST4vg0mOnwhA+OjfevdsxBVrwjO5hS2lLssW
fipoe91wjg9+y/HoCFGkAdBB+v6FhiRGs9S3kwebCjtCyLYh2o4qmMO/9PrZikbdzFpBKCMxO4jw
Qo1Wq7kD78Ix5ymPkiZnrgP3Odvr4CzZ5ii45EVRuDwIN5HLL73Z0JPe5Q5YrRicEQ1165bn4kkn
RszkeZ5ogknWEx1qhkZpdB4/IU/6OR6UiSvfAg9uPMCoaI3Ifjn2GcMgRzDGsTRzia553H7zNvpD
BlV56IWiQw4cqx9vNnF7pXWqzSHW2AkPPP8lRzIcptP1+Or+zJY0x6ED+TwvdKWGPHZDxd0vdaEw
7GSGI9zA4Tv0/a6pKnU9qbdBgSYgXcsQyQJI4EvyyVSl1T9yuHqCJRNTCP5GmvKmiJQAtvSbvC8l
1NO0Th1lUnVtIOjtrvFRD+ik9i8PhxtsITKNuB3rkGOcHlKs+DRinQ/HJtHL5CaTPzugQ0xFBQXA
1B3EzR3wu+IHNcoMqJM1CkI4AtydhouNehRnW0kxMdRL1h6gthSSad7onYEQUpgXuFJ4FqcvaaGj
8xcODHAEuNIj3EbXDQfBgLfs6dKQFzix4wQ/Y8IafRaKs0Eo4WNrt60R5lsCGPvccSvZji5q4O2X
w7cjntaCsWSzdh0f57vuVVWwUR2piYyeEAgrr6V97cYQNESXUlDEV8KOeLrRg2UTKFnP2Tl4yFYP
nT71t/UtzrwEsurHe1cs3wF5dFjN7rFQUwFFzGOv2OAJP3KUIfmLVzbvp/rIV665EzAQ3vc/2pY/
Zd82hG3R/t4KDKnzcbVmR/levkb+i8MNwLq+eZqqDCRX8YaD/t5rgStN7/YKqgfvVy8505xl9Yw8
mcgIb9sXyhwFMuOCy0jH2Oxfc7sHWr7BzqFlNZ1tqeHPxlGsE/BHLZ+o1H3oo2OfWb++RE/uLt01
h6/5oAcC4fSDYbtIHr3B0oXJRawoMQESbIIHAIprxUpYtDmS+ZZAW7UMBVmOXo0RhUXm/GE3FYzC
H1jrPxVgfchgpXpC0wF9HZQiF33TBLVxS11yWP8/cVaI1nx//EK5FLC21rHZFUy8Rp2LxSiDOyJY
SRu8lh6ueV02Bw2WGxbtS6kwMk3sWgABTYg5rC0vXtDpC1gl4Pwmax9LRNgcyl+o85lukQu3D9aD
1HYJGzC8G7G40TGj/pjFCHjg863XaEbR7r9p05CZfJ/YHMuvPTnabm7T9NsgjkT9TcbSsj2es1+W
SwzkZel29QtxqSocLmVXXztmzNl+KJZjL/5qLPWljsuPYpN9bld0KafFp1GN5+t3+8qKfViw49wj
0pzdQzbe58dZqDs/auBaLCZMU5kh3Rsr7pMmb3XpGFi1TqrzxmBb2Jxy1qTmLDesuoP0IMWaVgW0
8Edte4J/IfcQSOogcQBNkNvSxHdTTzo0mmd25+mGfE7JgdNik8Z5dQX6LQUjhRYCr/KqXDNN2iyH
rn3/17Wbb3NCKKj/job/9W4URu6uUI32EV3T7EbxtIZWxEkoTueBe07wA1gdgnwbm7fvmzHCkilW
WpeMoHcWduRl/dT28dcY7/v04zaZkZIBcO3PUL3VczaYNGkr01F8KhNcfbqvaBX4JTu9fiA7E+MQ
nvIK/Dt45ZPbStrRE/fd2QhNZ3//PNKCMg3fe5RoC0TU+cIpxJ5bjPbYsak2jPkggcg1q427aAtR
hFHfX7pQOa/dX9RF0VW5+G0M269ulwU7liBkGwYqkmOpSu4Xmz/2C/FdgHpqMKV8LTohKKyq0XKC
RL4s9QwZIAdq+i9wEZlpcm0kGuwx7Y71p1EpKAODZyTEaEpzQTGohoKk3TzoIKa2UpCIQzzCsJZb
prTOv4OZGHQJTybQzrqNTBBmZBiJ2tHJZdgqXctujb/u3yGI4yFnHZ6wQYqPkLH80gCkDVudrTFR
ENbcN9fxP9My6YPF3Lf//nOVpsEMANVKDfhI1HLs3EjtP3t6kZYjPs/0MAoJi6g5BpBgeGZCktba
aGtmuENhyGcRMctMJ1ohq+MkJxBve34FrnfKMwZI4YbfT2wu8+rAFxB3gfgjHAJDsY92R0v5jAV2
1QCRUz1y139gPCyEGrDHkj1+oLO+xGUJ0IdtO8tqSzQDIaUTVI8vyWUvphO+jJzyvrPGs1fbo5gG
yqfdu4oJ9iIJCNsOTab7LTEaWQ97ogYjlCp7N45RPOWUmJlF3UMyTg3JderyIO3JEFV8WSxPUTCM
G1B2QU3RAHWWCol2530RhTV49FvvI+1CqgncNfWJlq4Baa3ku6J/mIs5xQ53yW+/HIorJndUFA6b
mHR/aDicsZSjj9AAUM+vqzjF4ScfAYWtrqkDjKDQZ60S5n8VfVCvbbFbn6HTWQBMEiv2yJ8f9bic
4wQGSOaQdbrLBwtu8J71aJ70fcWtir411uM7Fa5XlahmBuCUOewVy+tzaT/HW+CR5Gn3edoBKMx5
W9c/XVKIFhtY/xDdQRk9AC+VfgER9xx6edRC+NIAeydC0VCNNZozKilVfv1PaLMukYU0XHETYBhn
lO6YoFs1Y0s1CHHAgJ7r6cbAhABl7la+KHMx7bi8Njh+x58mA5/HqbW3zXVDIel8yWs+k6Ntq20Z
Rb8W3KiWn3O1K/uLLPleYfa6NI2iLScZmD3Hh2dSrEanvJlDFY5WvUnzwj0G2fblyefiWyjQjQvF
mjrr6WKCqoCspOg2qzkvflX550SLZCKmHe4P6HtVxrJMhggafQvzcL3RWpIlb4EPTsMal4VkCNEh
boTc909tLC0mE9jVSa2sz0fbeytIhs83lS0uFFE4CjHGgLtri9BoiO64TO3XrfJrOeqbYnRetzZE
kDAt4xStq9hwXT8jhKYYTXRNPAZ8EjL65OYf6lr2qX01eB7jzxm3NPSyr4Yho9/ubFJPssejMkqp
4zo7pedIX8W6gdwxqg9YkU3IzEc4nMF92oxuNxbtsvan/zbp285ah7uy2PZfO8BOBCLAC6MFO8bl
sA6T1YmiytXK9U/xOORp7dBfYY1oDW9e2lgpXMP8n9/WbNhN5LJlkYScFrnqou42AEEsuFw/ixaH
lJXf8fOb+A55wh0J6ZhpYge8P9WkzWz+4a6XQBrJGhdwwSCJRw2RL6rHeH/VJw3gtCFM2nrnpgXd
0PUV0tnKEvi81CG4chgNQA3cCiryO5MfYMNOKrZUImhDFGdG6ev1Hx3Xy71kwsWULAJqVMSsnOIS
9uU1AJPryb4/rXVQBpbj5m5YsO9d72vzxWK56CyFZYxjsdxaQiqB9kyeNhAtzAaQT1T9Xx40m2ad
Ez1/sFfKztnSJfjDmAuLZ84V8oFZ/GAg2UGkBbGzUimQsOJYu74Bk4oQYDrBAS28UqFH3nQfWqPk
s39GTSKWegtU8Q5hpgIqKie/DDcfpG/xTeefGwV8v8AbnzCyEo+6pIENeM3eoRud6DlLP9EpevkI
0eeRpfKLNJCsf0mgh0sVCst6XcHHJx8ilT5F4PDfw7HPOoUEF9oZlGvS5kz82yrdNHyfceQYW3ZU
rtrfoXvxdcZ5TiFhnUb4JKwzm/JA8J4t0UzERs5894v9fvC5nF20aCS0lvLyb/eA1IVrmUisf1Xv
P7eJdBvgsrQqk1GllJYztt/r3rlUa5VacnUVccw/SyGOhwyj0BHB4mvKRmJ4hfFoH32IyFEPKUNv
r6mRGPBdsi2XX+sU6XnpamwMUX5raPBuX3JdFkEo/zliFJcdzqJzN7e4E6bsM+oy4msfTCJISVvj
2ffnyrLdCiKdP9oLtU2uG4SME5kGIkirrbdHMVln/l301h8QwbhJQIxhzhco86YUVmgPwxQix6Pm
7AWIzhSlYnmadTfF0y+DFrhhRI2+zvfakYFE/Q1vkKb/eDBZAJO+zUvfPufn3h6ogB8+guMB7Mfq
p/pIetcaov8Ooit11RlnaJbHAdTbF4pUnXW3wyQKw9A9qWycFg010t+xxjb83y8cWoks9dLNxeFx
eyt0qjcg4DgswG3A3PgdOTFDryRCY1d7nWsWEgo6Qj60ufpZgwK5QZwGOt1sklrKwNl7qOop5GIh
2MlEvaLKnJvmNMWSoOUZbTGf5BdmuWLLprdlhe4oFULWSMEf7m2SwIfqIdibtaC8hqG5CY191ygd
86/64TD+sHF4GJzaETEgx+Nq0WEBGRqoTrriCs25hxn0m8+n+9sD4ayqbOmY1PTTA4vmAvnxieWH
vSXKcHPlCELN14jXpcNb2bFh1DBvLIDBf45qWYIq37SfEYXO99kVClyJJCD7jKWhYpWErSv/X+bQ
pRyNND9tvzH43W5IoaDqt7GUY7IsL5nKw4HfRmVXi62MXMtnrLkbp8BPC2mAHju7lPVinI6kO+7j
lXnDchAkoc4HeAFUtfgOPVFwSEboB5Jqrd0lT0ezjVR+1hu66hoNbsC5yY0y719mwmyncwpHV0pp
FFXjtByRqYPey3tJJvhp/QVjxZhLSJMPnjgiGk+sl1WZlD6uKKaxi4tNIVDisCGAaygBUnsGp5eI
I3pLjdyrZSBO5S3QxR9tMPBFtxAYpOne9bJ2kq2chaLjYmjHCnDqaPNGMWJNyRJus4OgMymCVUkU
rmyWAH9UqPmSMCOU+Q6WdQSVznFHedrPDon+pWkzwpnJQzoHMAC2SJJfDDzdDQsT02R0aPNoFvOB
Lt0jYQo7K/uXjEH1ml6nBzQPEYswnx12/MXruZHnusGKlH0k3hE/X/cbr+SYaVOQAeG/i/T97Kd9
bXu3tvgk9m9fHcG5AljhFaPS+QEE2CgZVOP8Yjt/d+WVjKVY162CKndS5jPFrTK0z9a4bu81hfVS
nxAK+zOOgwbyhSryeZNE/0Jr0FZywNeDg9ixMXsrF/omcyw6lgHC/CDIOCCjoXp6INsDY/dcvSUl
B+My3n1T3rfQ4/FqRwrcvKQrlvXrpFXiBNqzeQYdiYjqVnlR5uBsMLUnK5TQ2Z4nrGw5KBiXKHGq
bXH6sTDVy3usc0fPYyupgCRBnGLbfVK5CFlyEJO/qABUCazGYw3K90As80bb/lFENy1i0UVYM6Fn
dqEM8P1RMGhyFauKTEH24+t+fsFtQA6tWxeRBFPhjEbvZRGX7E1ghWOGadSPEOWjKgXaSJEQgU1F
df4KUaT9Z6MBZ6s12NUZCM+dCvuNvXtbMY1Ovb/ay0oIWZznD5jJOW6xPTjy0TxsgEv5of2X6JVe
SPHOGsBthm5QPC/CxZWFRPMA5ALSv3gAN85aWTEfXdkB7k1HMLWhF+8rzduISp7E1yFf28/8z/Es
NIndqaRP5lmrsyNKZefsnXWXqZLWJLsJvH6F6hYIXqAHSTF0RG9lGjdw7T1TivIGM1lyKbnVIf1j
y8eS90bdP5dIt6dSYbTCMpT9hIphNY69AxQCP8aBAQVsE7pp5XoXhDQpWzbjwaykCLiFke1msQwG
AmxUtzmkpA/TMrB0I/eqTeSTmkj6/HXbp7AR4KbnBll0Scc2Aj4ljcI7WnGqqjwNJaJP6jA5z8WK
5FuCsxy7oxtWMQXw3+71kOY+nNVBJiS2IGbZ9Wt1Zj8NA/UTNCm/mlo0+YbZPXJ5zWGGvsR71t+H
FPeC25LtfZc2bkM+YelO1WOHIIlmoRkQn3SAklogBhXMX1rU13L7c6rZT6iay492lIIvt+DevOBO
zCBZOl3IzV3JUZUGv+0ldhZbB4nA6Bkzchn0Sasdra9yU6uQEDuuqhN2rvGN3dnLdHVMRWPsDSdC
CP15w4LStHyMQawLBoa8xHYJfZMsd8D0XkQWv2VOxaBx1geUbmd67xBNh1vp8+rg1Tbdzf5grveS
sAowxIjGWgFFtTJGnHX7x+/PBaDs06q6LrE2ic2h4HsPXY+WpG6qePoYRxcCrOVEVcF5Xrc4S7td
+RPr96pPdNS+cuQ0ZwalHl8BNqoHG4aKJgbjHq67219m/Bmi9Hx8qrqaxKO8j7NpTVHy9vpQHMT6
2NRG9BgpcTnfN5PmJpxBPxobxxUzHpfa3rS+BMWECcikADlVcGO9cV/r1H4NUDeAKqBlJcEi9mjs
nt6v0h2qzYWLWtkgIr2bM7NWEoYpd6btDT+O2PKblTA4cOiUIJmcxMQBPj1vhAtHhFGAUlHAMaIe
TuTHu8E8I3e35Avf98h1NcdRJnYPwFeYIQkYMjzBtjaBQKR80CPdiuK/f+CEgySIj68MOGYT+IaR
h8XWYWyMCIAg6a4NaJin8mafSles8fyUedSzNtd0GdGGsYjkhZooLr4C2U52mGJfbyzGaa2HUCxL
MJAGaG682qi3QQrmxLBiP7R1pWIPZDtSDfgbQiSRhogZbyCWgw8GAQ1obmTeqhEFzLZU+S2jMBu9
msskUeDEeEGoQ+kGY0SJEZhcBgiofmcHAzjIkqpTbug2lLFmzA1sKaqxAIuTA4M3PL2u43nNPSih
/KyLh/fVZX5Xv/xiYtlB7ZvPLeOo1rH/nYliQBh+RXcrE+MQCp/J0VL5kci7tpblplIgMRjxGHEl
HE/TmiZn0zUzY6LwWR5aqddY3i8QP/qSB3Wlk9RAQukzN+QqoIyxwZtR63WtjORlaYlG2JrCuXyP
Z5usdiUtRs8Rdgy7Ltlsk13KrAn3xZbfGGmxMT8wZNAPWQRsbifb3gxF9CADFaTb8AmhMkYz8AFg
j+BqAbQutVJifmSCXmyYSlMGk9kvSOL0VaJotiD0E/GxyQXiEd768Fyf90B5RDBeBXqJmIwiykEA
fk3N/OYdc3siDXfVWJwU7yJmH1RzpjJaY1rrIpM7KgC1aYt6ef3xul2/tRXvk2by0rlAb+SFalzN
XlukFc0qXiQP3twraZwT7R7iTtLIELJGXJTxhxGU2A+q+k+fO0f7EEM4lmkH9qoYlpzeXDducqBc
PO5dCh0qmS8AksdczZZmCHJm4r0UoTpejfoDWSLvY9lGbKUerOEEjUj6QR2UL5CKKlh+3i9fjP5t
bQ1epXBiL3VC9COUUPuJ/eoQLSF0t/wCRwCWXlIX+nMJ9hpU04a+HuKcMLAByZGJ/LfI2/QDPplF
XJR3Sz924gDhdmno5mpDh5K1Bi6se4CvW7ydELnm8EGY/Flds2D5wSv1yQ6x6FEeXWrYFKDo61jQ
Vg0H0Xwcc4KM9OOxWdEiW2aqM5VKLbya56aNzviDQgZVHFeheEo4CPZV3jdIM8w4I2w4GEKbDBi/
w2CF4HmeFseQ9IulaW5xd+8IekcS+MoometON2heyezO2uL9PQWFrudzytYTOXPhLS+jGw8VeR0N
qcwLm0O67iVzNVMvg6+4THu+NBlcLOH4JNQoWt0P0zF4PNO/AQ/7Ktiq0+24npO/UOsbGA1YgiCJ
v7Gv+ZXYvtDlbnAZT/i/G0R9xh8QG5oaNMWPRnAVkeocV3bvurqwhKa9FAWLZMtpVQf4eCELsY9M
y05+5y8euUHp2zzwCfnPZknwdBubP9lhIMkHWdBTGiaGb3E3+5QkMMiPjTeBqIve/yEd/L3UEMJK
9iFPikzK4YtICUmGT7HZE3DjkBz15lto68jnlx+Q7UPtYU/MDPrnN1ySicisWUMBcaNsmpNVdzsn
VOSSHzv09c7EtcQr7rSkqbxBA8xRuqTZp3Ae1lqtIXnNq7MCdsLPG/GJszKtUY6zYysXlRID5ftA
XM2U35R5RXLbhowcwXLywpzoulocmlZ8X1F4uPveGVr0kEYmM6rsdETW2oAjNT3uKoBwjDVS8sa1
bPYrDzmvMAkRJAM/eNq63hI+qyu5ekNHY1MoIKaTG380BaZS9NGh0iEqCad+0C+UqakbUBugsjj3
xKtLFc+MluZVIXs7F2b+MuYTOKJccU+2ihnl92o0YMguheygX6ifHPw7qJ54lYXbD1ACB0MpL9kN
VbbMgej2Fcl0xD8Xk4yJaSDZbO6M8Wm91psHDaagG/rbOryHjy1ecQpVVqahJWIj6UBXrRe2BpvN
gT9sMtn22vN7A0/23/RhiKyYk9syS0jWCQlF3iltuICWAeQzEYMR16R4bcw3PYKi1bjSdX2pk24K
5n5FqE3k1Bhr4mCHbLgIeTuv/YlX77LGYbpVx/LyL7fzjgduBanwwizGOC4aeNiT31GdMAsKToNK
Tg6VvXYfjSuPxVsdBukxkPwtWsu3lxzCTwIAX1xdw4hzZitVsNU2tKNyiWkLlw6QFrx6XofRKih6
LC8MPpcGaxjjdzcAY0rE38V2JbUL7QGOrcdi0uYwN/4KYOCCqiCSlcYnP8krFV48v+hGfETascx7
WxPGGOA2es2urp5rKfee7jg//TXPY0Ado/QOyy3X+UMB8X1LOKU6MLbdUO1iFn2tjX9VhizkVK4h
H1Xf1MNwVlM9zrsvjydhZFPd6ypQo34zajbVMZfdd8aVx5B0ZMgkDf0UZ6bd43qyV7FQLPqtEnxj
lQkk8SMIltZ6PZV1wcNmhxFUueRc/XUXfoqrJeUtAUnTwxPPyzRph54NWvfNsXCvftfvcwKdZTNh
oPlPfElcXLn9TGB+IQIN3TPitNnYzzxhUvlBvzVGmg5uhKOv8rpf/c/K5kdh0uE95wSb69nIdH5Q
wKc/abUJU18LatiAmigIivCR/PYk2QigHFcsm/m2jdx4sfB/tkXadigUw8DScBVUQIzwcTfr1skS
WTLKmDHrM9IxQcdO0cbV29UoJxW0/IrENYbDSFmEEjByMVfGex2UbhuDqITLYgrQb/E3+MdTGTJU
F/tkDrB87bTn9u9hMh+Sl56AiEfwTKNrwkrCBPc2P4O10zXG77gWS62g/Xke7/93ZmyCxP9DpWs6
XrneVfYxuMudt46igLrd12hFhomHZ8tcXKt6Q5ESR5H5YP99wnn5lWAbuQHrYWufERLHNdvNh/Q+
y9LSLKH04yc7FiDMXsaHb3BiQHkEi6AknUFJGyF6ZLVtOx3xiokeL+AeiEfmyp40O4GdYgGgf5vZ
pI+yRQtbYjEKOBkX2kVkJzCxAfbhjOpigr+O6Tp9oWmtFlSeZf/uJA7K9wUwmwhD5aF7N/V6zn5m
XC/orkxDnPAwrLcpDO9iT9155m7seTzJn46FBxO7wx9jI6omNG1x48flw6H8lyvcmb8e9HRUS+kF
ckAhDGgInq4I0+jnQJt+IAjQwlVkDX1bI9CIv8AUreLqkmV7WRM0jYaIPZiCKqK/F/mIaL/4iAoA
gsny9IPQ0ZND/FcmA+2K60GdbZHj6TyTg06qWwoju8uRrjYyEB6Y2bQZoDBVkAkcTyjj5ER/Aayg
+sxDB+iv/svoxb78c7/rkjGrG9U0QlzIy8DyFRzXFJTZARucdkhiN8P3bCkRY7bn0pVs1b6mJDXk
Zy8Zq4bRh5D5+ehM/sDyBEJ90s5uwYX6Icb8R4hk5XaKKcjaKNHt2z2Z/beW0GejDhwj5pKh2TMT
az0f+QrZMEWjGdtytJ6xK7PuIL7yy+wFaPCFF3sRvp8xqtXkBCXeDZevN3UB3eqAwXX+5SswkopN
Zv2AeUr2EUrUOqTbUkk0/YaeuJySi7vmhYGSmLxHcZATePB/Qtly0f7S6XCuLUf4qpQdPmJqMlkN
bE44zH98Iv0PEvMZ1yz+SORhYUacj09FRTuosT/u0aDpQwu9H8VVAyss7rOBYY0xj67ihL3Mh/vI
ojSKEYwhrLu4uWOnjxV35OkOHCMOj6VYFTNrh7Knvg/Lv/PYSVT7yCNUCCV+7fO54QmyFYqG4pFS
FSH9vT0ZpH6F/rnKwLWHkOHFn383kbmXgQ690ahFfLPMcx0zOJR+Hz3I6JCZsQ7bLV57c0gGvGei
NHY46M1c6B/g8FqKCCMPJoW3VvzDOElWJj7xRU6No/1qauBWVoJwQLCVy9B9Ipwpa3HmCGA9Cji5
7hlo+hioNfTZFsWSDthQ8CqVyBmLJbIpg/pE8OXxvzBS8VqbOLVV9XM93YXeTkrq7woVKCIvPT6g
cbxELAuhXfI7rQXyxF3M3mWgDPD+Iz9GRhZUW8WoeEh7cI4U+kExMjI8y2M1i6miKwtPcw94ZztO
JEJHRWrmmRhmACowAkBQM2CiqBemajKNEO7F3tZmHyMMzMgRmFKEOxiLF2uAMn9xpssMM1CNsIVY
jxUjM7gw33iKBzZl2IsKnQIeXeCPV160Hk1KIjwQjhqrwumciPSb6pRMwhMgt3cgd/pxzzLo14Yt
3U53C8vmIwCuLh1v/KbSSbGnumUNCZeR5gf+DIfdrPT2tShYKjTzfrVIkI727MWt1oW2UyikemLE
+ucj/3DAGBS/+jp7NqNTZwMY6F4DwCYmv2ViewFgMGYJlWuvEGFPDvLJzlVLDciO5MtVFb6zwkO2
RBrGQKZwfu4GmIL4bp91eg+uur/N713J78m+R6n5AFl2V3ebqZNBDXI/5mblQB7tTry6pIZvYz+t
DGBzrWkxz0plzPAJx8MGCJIjlRHP3FAocp6EIVVsxOLNsI1ybMKj1x61FLJMPYGXtJa3eWxzEO0S
rVCpUuRSAKtZjFIowVSOlz68l0pDs7MZwET8EwvfYnOUCMDinybYNlu6wyWmhFwV9ycwe893xLpn
IsPoHeot/eiU3hNqw+pfm1wxqtaqrSDoHdB6XXkV2sWvQSpRpi+dO4yLJ1lYRWHSph9cQv5QJr25
TGpO93f2vswUxya+sLqv65GPq8O7j6ilEqnsvqp03W8bxubN4cfRZc9oF8CvNSS2mMyZkYU3w3wf
VFsBNeTODPE9vt4ZCC5j+YKZ76k0OgCFWYNMYV+LawZDL1BE6eOjA8m7+45ti57jhiVELyY0irD6
t8mdnnkninRCzQa+d0fcsd+b441sh5RqBUUUt1YTl2ho0spOA6hyUaqrrh+lXq8CMbRcB2VeGe/Y
FVO5XBxaE9GdZiGnhEP7ClLd+bwEZTY1BeNH7eG76QBenwfy7In+Ym5FiwUGKNrJwtCIKVZaPIFe
KdeYDVUUZtFiXLt1TEQsWwKcCVHQiaHt0dqWdZJJZzz+Yp/dZQFcVMhTxOR5eXzE+TV/x+4IhQj7
3EJtVCwCEXaIEf/UitpMOMklgx5AFyIM8xuUyx5g11RF/zjnU7aMgdAkLbQTg9E9aXrlMopGdq26
8t1DXzk8r1iNHliyvE2QfI5pmMY0bNgWEGLtARJtquFrDX/hF1dTM7VRGzH45F4nJaf9gqjSzXMp
OxfFYId6W0qh3xjcl6tfPzrCjehpH5JN2fH3XRDHqJuwdFxRe9yrsb3vcWFLJG+Sh/J2Jrx6jt8R
/iLvyxFVlwcL9K/FPXrFcOslHwDhT5Y8Reij8pGBI9CYgPwCiMpnstxre+5kDpn/ne73pCwRsl/B
SR4oaSWwX2YD8HGtsSvPwXGJIoESYic6cpoKTisNz23z2tDli7qAk6YlxDDcxc5OkrLvTjjCRKjI
0mRh0LejDw7ihtOSp23bG3GlZuABnpoTmEAifKG+rAFSSuFa5th2gx9U6SD42y4T6ZfgDuFxkdBA
aDZKBI5InMBXADzcEkqvggHwPrpxeUmnaGx9UE6buoSrAAYAOYTMJ1jv7RepxG8+tJOZ0fnr1Jmh
atzEv4VhacWKoa7frDj+3em5bV/KPPA6kkSXRyt6ksOM1nLbgXxv0je+CKC7Kp2TTdgibBfnlr8Y
32D+0Q9dEhz9cSWTP1JOHJxj3LfNXXGoxfGxwcrXRqxqk8jdotgx+m8hPUdQmOeOXm1acQpAVKds
PM94KblC0tSOIfLbIUIrOgOfUglDysZriL6I9Cwrxe4/qolY0dUCEAcfvxpfmDEuTz3ho2gC7yPG
gyVKXuHuTu6MA3eQmLewi8S2xAMdGmKiUV7CswrJWiUgUwxq9nq8qU8DUiPS/daYHUlhpioTie7S
vnx85Mk1YIaQUFTnOZDgv07p8TYgZtrFvt0obkzrVOcoQLuDQTPBgxNuz7+TFJy5iVvonvQ6aEEs
fmTgT9LweSXxqGhUUYHnAfUnQ68xsQur21DGhLoqrAxspH+cg35oUKM8tge4g0sgfVKr9oPnVzCd
E20fHX1PhJIGbCIfrh6byExTBlgHLocy7JALvePf/YehEuuU8y5K42p0yp27DUWZWhBUi7BDWzQL
csG71b5qtgzY3iaSl+BLGOliAJ3tCPu1Aq0lORy8o8SxiZc+97vO6QzbTJBq6AtuoT4tLrB3w7ew
/MW+GBaQohyEq0Wn/oWEA6HupAUsL42H6sE2ow3kwGv8KcpNerc4kuIE/pV0yIZOS/Xdi8RNnWVc
WsTVxG2xC/RwH+YL3h9gv7svvEHk9HEZ71iOZF2BfwpN5M5xJOsl9AZkuKLaIygYNgpCnZTz1qAm
/sT90egVRa3HdxbJe0FTtnkNvtyR85XowPPNX/k5Ez0K6OB471TsMgzRA3YQKj6WHSgVRyFcAF3s
c86PE5fLNGwQLu7S9SkM/XXgvvLys0nlA1vNKDLGcH5dqqXmVxPpvGVyeZkWmZc23E48tqhWxacN
ULe4acqS4cO2wgmDHIuhtoQa18qGrBdKOhlvkaPC40wBA+11oDgzzYYdMLNxDbIVSPzhaFQ05nXq
x7rvZXklaszAkY3t77FnEAcBMB3DdFo9Wg4+eamLwLZ0e6Cs05wtnQSnDALIq24PLmMzsSY5moav
VSXsqb1CgvVCiixNqTlVio2UXC1Al84GsKY1d+YZcBOHMBNwwvKlzeUA7rPtodRJIRiaK45/VWk7
Vj+O7N4pL+xEu88v+AdYUqjgFAeaDJQc5AM5NAHVZdaOi6vU2ZCGVIihp8I57K/L+CUrER75slyz
t0POT522XrMSXjvt2IohgKMUp8nSxPe6tpasySyEyaCvuzOGXJC6Twqlqfn+J+HteBHRc0QLdSfP
Gdwqm9ZbZU7Ip06cB0Ooa76a4f3yvkjFkJfCedyIVfA329FJdUnhxjs+zp5U9XTbvJ2b3c+wIH+J
maf1oW2BoOjLl+ag4uYHFe5WjcUXLmuqmysvR9Ka9smE9L3T96znPdzW/SObhVwyDcGn/GNBBL/R
1xNRKuoKzu6FescruRmye9H+5h6NOoPxoWWqZXc+e98D8e8nnqSwH/njB/q17x6/Pfbij4xqNwJD
S4P00RCV1dfFeOcJG3X0BFCFQlUQ+JjU2VwDy5HCIl5BIgeo5c7QjP4oh9ok2RILyopaQV1q5PHw
mJk0mxaKCRFldSpN/VuF6zy60coDdeMXFa9bkFxz+ZZNB9mAYLN/zeq6UiMP95FYmomOczVTAq5p
onkdeHy5n0qFM3fvIoIbkJ10uHlUNDXRrOmTfhGr0GFOk8XBSa52pwapKiB4rQ3ltmtcaLtGBnN/
+W2Knprq/Y2FPkiOXsy4yFPxjnR866lW7scLHBLebz8lZ9Hj+3jN3gF+Uslauf4liKQV+kLh0Wdl
2SLr86p0IDv5ZbRA21dTNQMQ2IODmKAtHbWNjOcirQ8RUpIu0um4UpXZtYX7/VhVA0LgRq3BcSpk
4ffNpg3ICT1urZIHxKb3eg07YQMXvPNQZYPdt3W1k5H7DLp/1LdtXwanXsFnuFmQxNdbMfOfqhjr
OBPo9M4Vr6u9dTdg2+l0cRsrqDwIZ9Jd4AqWdFAR+3jADn9aKi/x4Ov+G6Zb+8DDguWWK8e7i+Sk
zQIL50mOzNyFCk5a+DDwuDJZ9pEvThE4mDAj2puJ3W4aLeQ7G3eFYaDbqqqzUpeqcPVbQ2aaYVuK
TKp2PNSXiwwAtHxeTTwHDdBD7/BqDcYCmqr20iZvPwlJ8+ZplwlhdtyPII2oCE2xHbO1t1wr9IP4
QS/Gt27cxxAjwO9aNkvE36kIm0qnUmeeNLJlO7btLwuyA4xnl9yBNjFfxnz6ChDEkHaJIO8idBYq
56LjYDdkZtM53ffo1aHe1NKsU3KgZqpAbyN9rddqZPnJWt5AKu840JPRjU4uS+9+ft3x4ak2D+s7
stIm/ITfMWjI9DhM6owPnVZZv5r13bQD7ZeNJMI/LRK0dHgJNY70L8OLIJ1EuorMmKuxSiW9sl1g
Wpv4vvp1VabAl0uuoBUIkKZORqmf19zkQDtbHmqq5iVjrwAB3a/ipmz/Ifdc4iZNszu9FS8kC0mu
ejHdhwtQtRePXQz6CukdZLyVE5hLFBd/l4ixi9cps4whJg5qn8nfIHNY1BK6YImsqe1wrjGJADSc
hR64sZ46otu7DohVv4ncMGmpukL3cLXqMMfcTlobxcPBIfcAziP7YIgEEt3kpB8XyFgtQYO+yEM1
uEwIQ/VcL+XTzoZ6rr1DMbN6qKguNGkBeO8FMbFSecE69gu0slPfxtKnmz3A9Iphgef9Y44St3SY
xIL3kQexLykgVAT75C5ePpPFi2iAW4+dMfQX/tvsVnZIrEDpIBdmIsuSvGWzuvgdPuTM5XKQ80Vb
oJG7P07OlgFoFBpgWgOTeTg8XLKOQ9taXT2D29aZlQikCYtt0Q57umcrE6DDeAiltsMh/n4GxGuZ
UFQMNCodpisQxyTq/EJ/OntOUouDGl8iXmnBYua25h/o1cIqcVxKcaGDcp91Przt/P2lcOX+Wlgm
QMtvZj/PXkYbBWvuXPJHtEvQ4kmGkGEeKaxV95FO1JOvfeo8tTN2aA9kgRhAy6iFe+DnGaxEc5k8
Brahl6cFmy8V/90rQycXlI0hfuhPzZSaW657uo71ja8jVgtledPuKnppt+Xxpy9qyXR2yYwsjM2l
zrBX8lnspZ3awu+F5GuDg8NVqBzwN5Lbf7a3+h0dW+x2yGk1l15HuWSeBm/MdOSSYk6ZzhSPAzKx
oEiACbeP3R4Ajw3MYSY7oP3fUkXsUKw91pYjL/QHRFmuqVvGqFEyjYmxMlTrVHwBIzKoGR9lZDFK
Q5jFL6JahMi8D+H/g/udfon0kZJ2UIN/QUVFEkWGVfRs8MH+IO5legwlddYtZD0tU61B4IEegHWq
h3repb2AQw4kVHEaJBZfoFqMINLLmMT4A/wtbcgOb857VqsGy5+eOFCzd/DeUaBer2aUJm9Tunsj
tSPVKyXeuoi5eSKFjSptrF2WipxoeWqGKSjlOx2J4EQ0JwuKCbUk/TMK653nzp6j8szdT27pqLni
GYVut+5HuX2EBDZ61x+/weVWgwO/zRI6P0Xtz5NRFZVX60V/qtRNxQkzHHwiJKpn9W19NQVli+Dp
3Sil/IXsllHN25O7h6ZxDCKExZ89stqarlWTY2sShym5WGrWTU+UFjREMRWYjMnkKCrwuiBBkQqA
8zA4u2EUZxgbm62Fd4CDedk0ijXGJQoC1aXI/j/YTaafFutU3mQ8UsCQYAPuLPGGM3kOAAtP3V6+
wPQKL+twSmFX/o+UWwJu0WPe0KI2AICWvU0yiOejgGZx1iuXRRKV1qgPH/btjKhsPX3xPo6Fq3dQ
gMKYzd6opcUWwvZyHj7eHQimSQFF02f+GQheKxJq6V3QKXapZ4ceUy5s7EiWa7eoND7G3zgBd2zu
GesmIKoE56YzPF/fU0GXgCa/9BG34MfrWDf3/cPMGryQqZcr90cm9NpGI7agXnLWR86A7+EpqnbR
hxCHBd67rBJ5Hdr+/9KqntUa8j0wacdteuD+BuTnMylbLtaQKCZHJ697zD4FZEgI37qsZvs4u0p0
36Csnu9E6uJnzBw+kIxBDczkeVPFVhwq4L2Zx0ZhmC7nMjWc4Sc3JeE9ozrOvUjj/+G5qZ/UZ2gJ
/hv+e1cdLxt3KouIMKsWSMBADlx8gLM1Q3ZReR0KD9nhrZYqDv0zypygkNxLNgb5nvalG0t+HkEB
aghtgUQ/QnVPrtyx+PHukWBp8PmKY6VtWghTbCRw5yYun7znj7KqfitUSAG6mfAh4vFjyNfQT4JA
oJLtwBF2Nu9M1h++3CsBgk04Z5Vr/6Z9Plvt5P55X8bAQTJbOAcOdKrpYZXXtmwz8rGI8mtz6Zgp
t7ALKuOBEAlwZvP2igFJbqxbVDEE6cNXH+Hv7hYcWcGdPxBnfSDpXqAKoB1iDr0p4yQ5cUMv35ri
LtdB0NQ0q4Mov3tO9jp6eUrUeCK7B0isAUFzzT3rZiJKpeCDnMno1Lxjz6b9CR3w8f4ogXAtIe8S
K2TGevSLTxRMGc7sbUKeh+6953zGTPsybPctLw1rCDSOgufu7TaVpk1Ze0yqB7G8iYBZ7suecywn
cY356ZstWNiOxshUKv1LQloF0EZkBhJXuyxgCup7E9nsvLoiJFKD4XNOrvFi0oXHNYRO6anBYXWw
shxiTKt1yPq3vUf1uN6T6VnBVvAZEjgEVWDiYbMm73XevIYIMhpC9UnYMsaFi3bnRRv/24b8IWI4
vhFKS3wHG2iHaScDcwrxTMfPFeXLu6z18n7d1pAignGCXC/5GjdjBsqUbSg12prwaND8GL8l4pRj
VmzZNCRwHA7iOO3gAfOvcrbHaFQJ90uiZEbg20hzRmxa8ida/YIlkAFcHmQXz/YuPum8s+6nSseS
wNT4przvkkB099LFbfMm94q1dS04nd52AoFxy85QLj+dEqkZSsWQyXR88IR4e66YnlThprVnGHnE
DKwC2NuAGdSloStBIf8xaA+bSJy/Sre7No//vGQfO7eBR5Sh/YEPggNbgndg2Hypy/viewIDsvRI
KtUFi5K6LuxkdfGvDtDmORL0AKRek8pJFfkyc6ZcCw22jdB8AgHj+8e181KKOsGPmoX/RdjebDEs
B0ERE9x1rkH5m0ene2koNIwA+4oJmmeuDCQGXsCqOFn2qsDkSi/rQr6TnVi1PvLc0Iz1ZzYT/V7C
YxrmdFEQfMVIuPs/nsNIou8iEo5TFqQka/aWwqdEVChzr2AfiBCQuJa71bVAXGL9ynG1I1I39kub
432SeY6vfn8dUDm7QuYujmNv56aGb/l6UuEZh+SIianRz3zTRMNpIVsVmhpcM8o2+E+lIpnyQxwh
cciYGv4JTRf9QjbZHKl4uqrUrBLb8T4KOLUFY5F9iVKFkJVzmRvv8fpSKwpvJoLbVMdd/noTUvEE
nJAEU9jFrOfzpsWj0ev7XmfyNxUKgiyZTlzLESqbGoJe5oLO9vuwEcvglH2LPVwDjUqiJ8rw9Bjc
iRMeTq94iwRfJpFA7d7v71uHymZth53D/BapTQrH/F/ieb5ysEL8ohicLiDz1Pq01XlB7HLnE+If
9KeEb640j9omcuDKt9izqfBSFM3vZ35JtFBCxjG0wdBHsqUcx+TFAJEIx7gYikLJOibqhjhwshtW
mLeBPF4X8yVBZ+ISZv3lNcqx6eHKG7DPPKOO0z/vo/jzeP5P6B9ZCFbehIZ82hfe9HKWXiVrSMgv
wUbciVuxARviD9ftmEP/m7PxhbXsaFHhrowsjNwdEi+hrUVZlgqmLevJDOqJUjnApW9GXmqdOClc
QIV2WOftWG6IKZTHivoPYFEe5ZdE9PZ+CleMXQRjWDL5PIVYi9HBE1Z6G+aI9xir0XBmSX8OSbf9
+91D6/U1/zbpmmyzF29BxujoP9AMZcZX3kJfLHTS/DtLt7bOIfRc2RiUqNWJeB9MbwwHd28xmr+L
63DUm0AuZYzzXCSKfWj7CJDfdML9yYcN8OiqaC7iZ0Yy0gDmO2Sgj4Fn0n/GjiOc1rh5ek6JLJjL
k2JeV1X+pbNI9QOxv9s2p4x4Yqsq8o38Z8S265ct3hYE5xPQWzVBBgTcG8kfttmCwdeStuOos0wd
OY2hGs7i0w7a2Z5XXP/7zXvuyHX8OhShvVZJYfed9IOX0j0Z8J+clzuQwmYgYLuqMAOdnoOZ0X5A
kZu8mQ6vGD2QK0JIAU/VRqJXbMl2/1uMQbR/fPwYXsDr0CYkergoUKL22QcvjieSat4yBCKE4O4F
A8dCEMCnNLTEe8H2pK8cMFj7CzjK5ECE1QUfdQKnQ3VD8MN9xsWz0YdUHQQrg5a8j9WxjTjkIEkw
XXmwB81mop3GZHFeE6kFTUtMf1E42qW80TvGJ7rql1tCbzGW5Fv4gC/ZjQ28Jar8/LVCyxElLc7C
EjTIBXVzIV2bhTXK3pgWomb9XJIfI81LjMEa/gxSIlzpS2auV8oRpT6p8MTpaffk4Rxj4K9FjNus
COVkrnUz1jnSr2LjVwLxqJUEKz2WYETjCkppZS1qgok439YKL6dBKu0wtdlnrf+ndqSV+oC02prO
ZLiph7W6rLv3LVUP0ixpob9hO+Mxh3TQyynCCYmtPSbQzFgl4QHMHrdpCi8Ie+NWO+/Dgm2kKJrX
Ms9gjUZTRm79dhOx7a7rmsIT5Q7j8/QzyBaLWLe5BrRUmq4g2CBS2N3Dzsy83AawkIVvbBDG/3oM
pofCpEcmXJ+vkG6Ek756Ig92SvBBw+C9ma7dBTMk1da7Hkso/FdggP0+e+z3z2uK/e2GSh+pjIhq
jDU58R5Z6YNpIq7S2PzuqYGpTDDHtY8vozCQdIauoPR2RdoCXDk9ZOWb7qiwpVGgxMnxirB/Doy5
gGgzIaznNOuQMsE4ncB5p6jAkWlXBXMVBymyyfZQqiw63W+pB8bUrIydkcJskcWp10SsQXRo5eT+
fY5BIWFEuVLmXfu9w0BqWRx9dS1IBrePsbKde+EQT4bK7JGoDRxSRB2Kig4hicn/qMhOjnknq56G
b7kC3P1JKhZMST5fhbr2b/Mj6YOIaCikanlZOzZWj44GZ2I9IoFXWyWYaoGvp1ZXDHbdq+Adfzf3
qyCSmt6oDlc5Ei10ZNm2JCfOcTf5Yrs7t8hGVNPTjTwxdsZrnnyFxGdgO2yPBAn6y9dGwqvcW0JR
QkateLYp2h2uGPeZS7Qp1oRWNEoji82Sh7HPiL+/XLvnJtGjkwUW1i1vljWRDhtQDG7MHijYoEPN
s5r46bYvhXgJwOA/pYfaWvUpYFTsfCgo1SR1HoVWIZTCsF5SZaN0LYY+xhhbR1ufsyi+tqHJaKot
e2utEhzT4OCrO/94hxVjpctxUkHRMm20Hz7qfbdPHuCTUC8SFDn4X/7rI8F8rBunWU8Shj0gd9K2
rxY7LwQKJfPaHvFdVYxMcYT9a6/Rpb+xGNdWSecBiG1hg+433NSRgFCpkf7yI8s4hC9bo4Moai2u
AbDJH+xV4A+UWRAjRrrKCtEzbnqFRqFwjVBYSv1NfqnmAS2doHCmpNtZdAZ9vYo8/dLTWqasL8W8
OzaBGhDxSYgot6/LBoEfRYMula5zc9w4sUbJqHpLKTFz5NWxERo3A/doEG+9MCs8Bk1nOn2FeyB0
VjdF5fYMPXEyipIDjSFrwBNWUV8IWqddxuLoJq/nSC4r6XtT+y9KgI1NJMOStuLiVJzqBd3oZnf4
g45BkmK0umIYC6ow3Lp9VTbYKyqqZZ7gWuCL4lft95VuUZc7eYuEX8hkAZMTthEBhSN4uHn4iey+
XN0hZHaD5jciD7AdBwJWyS3+WuveS9Vy8/YkICNvsZNXlUtkA80leCx8kldoXVzKJi5KyCuL5hkF
JYKlqSWyp5i9Eyx0/Ocd27SKLsV44jW/43QvMmpNFfh3rO3Xp1QDhKWK8l7SE+qohSSiwOOd9EZf
FuNLF0mSotLLli64f/Kv9SvPOrt04QldP3zhBV4HTYyIsuotzheHjkjuLYEz3/PHnsDj+ELLZMmh
URUt7wjgAR+32ZupS+bfmwwKVCi1nSnvQ/1RUhjYH4BA3EpeCuL26LyvSvknU3IshfEE5+c2QuD0
z+2whnklGHY/bZT14lVRuimAryoP8rTeohcCYmDYF5ytEphHXp6VHV+bzjuSY/vUsRGHAVqwUe6T
OdeE0lRi5WfWGahpUGGrkJ+pDgffqc8v9LRX05sjYJIKlYYe0Nccu+P3jYmJxy6pwNHtOl5hfxfZ
JampMM8EF1RU10fXgNgGiRRXqt0iCg5Ol8W75+0O2I4Dxb7IiQLBjFakS0ws3ARabxtQcYoPPhzB
6o1BD+e+SWwAOiwApTos/rwOJb97kqFoVdojprzuZGBUQRsslUO8xaxstel3NahHsRlmyMHyyuFz
bPgx57CdnFkksMe8P+qEvBBAHNQ9fuZmKYR75EvL+TyoNxQYiRpc6mdijXmDc4qq9dhivIChl0Ls
8C7WIQe5Xt3qS1k4ij1Ya//S33y6LmcbFBkc3KhiXoC8Ogy3m2zBsCC79n3TsQg2wsFW3R99lpkV
c9qzlIRNHxMzQRr4Bv3VlM8qUsfJ4oYvbWu+C2o4XOfWArocsUSkiqFDjmFCadNEaLApMLE6pw6i
zaCSe45eGao9UfK+tkgQEgiy7TfkZwlPvemSPj1RkB71Zp9xVJQkGRtEN5BDoa0Hk9NR3jzTZVkK
FrTT7azA20W4rnkbD8sb9upPAUwbX37EWtaR/vlUTk0SPGwNLOPVQFtHLyTCsiB27ly6jVGcfJna
1swIhKG1k3kk+mYJlI87R7CLNvcRT3gT1K0Czn55EAvdYX3Cv77Eb+JdPPtclcTjqeAXF/N7n5fQ
6Y0durzpVNDNe8bXE679Poplo+1kYof+dEcF2G6o5CPobLMu6P9AViPyJrkUvV7a+2Zr1d3FyEyH
KumcCIdDog+hcHzwT1GmlMBYTSUveMXEzfUF9dULNkc+JGdEEzbXYjcRr6WeV5nOBskJ9aWy3xpJ
Z5q/mG1GQPOUzfy1b3GAOK9qX9yaNMVvyA7u6Mt1j+v+YOg6u4tda2fd93daEMqeOBVO+nck6i/N
ozSdLpdqw4Ap3fbpTE6jPERey5npDJrL+Kued2eAmZJG1oRwaiq8ULAenEDOfjaYK7VSIOmwBolW
xo13mE3PQmoLim2ot4jGuuTzd2nJVGZ529jrDuHME0SrZzdLTaz2pL0DnLNENbQzjmhs2O2bUtDF
RnpIm8t5KA0mMWfmQtLqVEl1rsfi+aW5fv5bA7Yps8DKvHx8fwrpf+UNaWcprHIrtjM5RqFSikgP
v/gP9Wrh0r/jOOwLKD1RwElZdcKw7JU8EqUl7mmvN5p3/dC8fTAfPRdWQ174GRjvndZRNqrbLWng
ZoXes7OGWP2CWAZfmSA5L39v1ovRx3/xVO6DmQN717KA9U2fGD6kYANb/YtNvDRBc4u3jY83pBLs
xz68JKGZ5khK3gFgfU4mH+QT+2J+Ba45w4zSSzeNr6zH3dwJ/01SlTvCL81B59F7T8jELZedC2co
vsLipn5DBVccTXuu6HWCbPSI4pVRcde3bfJSCNYG6/JDjFr1y+EGdrG5dI5I2SDno0cLfk4HET5J
IlTxNv7I88ancJh6Rf7t1emkQ5Fzv8h0RGofpZ1qKnus8tq/ZpV0LpSNZuUfNiC+FCBdMUp9d64K
UgziBRyI4RDqQk0oiK2Y+C3pSDL5c/68YbYuvj1SnpS9nlwIV7ChjZlm/hLDQdMHiLp+Y0kiHfVA
DYIaSMUzlN2qqUVXPATDo2w2SEPa+ve44vVKgTK/hWsp6krH+il/0UqJM+2bU/TpFSkuK0JfF9s3
6m+wfUq7mGHT3wzlLOOd7YdRKxFulmgmKqOlDZrMPMEW3NiBQg2xwY4QWYevE0OTXeugPjaxE0Iq
sRtaRzD8F4KTKVrFBFzmqUIgU5d8n1Elf0TGZB7CiGANoXN94IsLwRAkBfdftNf+RNttpVeJxILk
63H92gR0xQAZCiT3JxnCOxUd59HlVsuuTdtCP7Zl8bwXKoppsvsZ9eam/wX0L+Lxr2y5n1egq5EF
um8zMKznHQDM6P7+gAiXY7ZGs2FfTgRX4IxfHZlXoTn8O6qvCzOnGhF73FyHtT8jKq8GVuKApmVi
7Wak6P+tKamF2BeJetZOq+IQLg98Wm9hxZGh+7Iw0K1uQoaVuyvhQQhIVYnqM0zWxIv4NPgEh8Ws
oWd8OtHdB8pk59A6HcTGPj4RVHVIFI+G1Pi8r762BokqDCE921da98W3EtMfGbo9bMn+29yFdESz
R5S4gG1AXl0MFhRclqUk/ityZBdxdwEUBPzv4kPw6hzBJtVcR+9pfXH5LHvYk+/hqZ53mPZT6+7A
AcLnNn3vsRplLD0MgAMYMysS4zmOedEOPY6/h7wxBrWhn8cDUFw0Cm3N+NjKCVqHeeAsmEj2pNvO
6ehdx07ovUkaiyRxR9g1xSNoLN6JmOe7nFtFc6zbfDKnPiSbvP/8JLRfgs7ZlzG5zjXKqO+mrS04
H1QPw6vfCYXhoQ87vRh63ppXbdwXw9gdZL3lWa754Ovg70n2nxi92I8CDDTeCCGO4xVy9cJ5ZXqW
OvXyO6ZrS+YQ35b9mIgEKhGkVPGwzSZyd8bcLq/NES4FW0ds9o1Z5k6D2auqK+l2wnqrSc1Qo9EG
oCPYfSWAp+Jp5W6/nWp8Pht/r6cmh5AEADpjjemDvBRxXOj5IGcMDx6Nswa5ip+RkPAkKvp6Rfl5
Fuw4H5D6bBwd4CeqrcqHddTSvlYPdeWkFWwdIpgBefxA7Q68zPevLNJZJSCiPBQnAdiPRKjOtM9X
vsVT638tKxaPJs4bkb93SKHGBnoTsKTxLSbyb71dHVTwOSb5jsuYfqNPPwnhSoFcUOBeHDdMRJKm
IqwGH08aW7D1gin3Pr87xqdCy6z54uFvx8+LbnJfNZ6iEnyfX64jCNypTSdOLOdGbD+tVj4sb5h3
2fj2P2Ltf9el549RMx6xn9WNcPY/DcmSdwI99BCouewKWHfVPShREohWWwQSLDEbcUZNOEp1o2Dz
RNCJaCAH9LyMhRVhh/DQ2LFDcQuLMNWVJ/TuT4XzgbAgikwwa5TL2xlfh5GXZw6/cvzZiTNgwLGh
6Sl99KQdI/HKOFVbfQNQ3n2f27iWWPDfDZUcQLyxlvEKvQQBYaX+jvZntidNzDAMiPwljkbCjAfl
+SRN6v4JtOhpLaz2jpz9gOSi5E/hGhFdIWcfRwXY2One4seJItdPbbFIiXEuI3LyeYbR+ueEbH7A
jFhFb8dXiQupO0BagOl3uWZ0DDSdRsigtRwrqxqYGMtQ5T1MUfNkwD4Nc0k7UzwWxmCMPYqiiZuQ
3uiratREkCVmAxO5ONcySUE+nBiLIo+F1W50lUrBm6sgP56z/lykpceXRiO8xhoEIsTLhlicoP0N
X13lR6pzlArFhdt3mbUk2TsMXWGx1wNEb/wNLVmRzQO6ave9lQANe76onFf6h91MLIorTpxPsaPt
7hUih5/PZPWzPJh6mhDy+wqmGfqVsypfa7iTAWLAn8aIx2jm1e7p09HcQjGvRQcOceMBc3zEt6Ad
YjF6thfqVqFQ8cjcGB9RHwVawcoHIrEjlIW2bUk3OhwHrVCzKK36iJZfTyUA9d2udzGfLZDMfnfM
GbIRW03SCD/wfg8NVSBisEKrUp0vfX737o1NkdMW+E+HYILy2T/Zcc061S9Cw+gDwNqEUdTd0ldd
YyK61KEP4hzoJbzeea8J+l7/vJYVSsES3SIheF3jo2LhOa/p3qYbaGzFQKh7yLDlO6bL6cTS2Ipy
+nG0KvWwKIea+0VWhMHV+Bo8GEJqjcQwcyGDPkTvoBs7cT5tuyhQdIettYT8SKN1KeQKra82wKfs
T/trI6kjzGeqU3W/uYJfu00ZG7vSSCSDqMcS6VgH7N/JEgSfu3aeXH0rvo9tl5S06qf32s0Qc/ph
4squ7M+kpSo+ugS3iGjsd2VacSoBPRSmGPhQnLhruH9G+FwhMJz5jzik9dfwQ2aUb7FBtgPJ64Tn
z4ZC9NeJWuXzN8Etp1BvzriH4Pt+FyWcWcV92dURoJ7rXvChbZkji/ffNlernz5gay3fX/a9wgMa
HOZPZhyEW3IUHJWjIxbyTCHbcKFzw7Kf1P08yKIKr+kYxwL2fLdqpEnqSNXaLOo5XXNzpG8j2O24
mB1/g+3TI3Ox/w+mqT57tzDfiZ1tCQQwJMS3KyD91Dj3PpLLmvftJgRPPajf7A0KfNnQaWtNoSSs
3nUjITX3wZunNoY2zVXysD19x2Zg+kT9BIIA60xxCIImAgCad3LTI8lCIJkwIhXca41OxSfqc2jP
c2xs7gnz5l8qwow8BTr/qtYA0SKtNx17jkdoVpaM2EM33J0P1EVj/gnLvfUyQm+cv9splxU1HWHg
E1hgoRiATvgkeas4N+VgDHBPkUMJYLAsd7JpMyWs+JgUpyJZ+BScYRElLiBjxIh39KHWPIXWomwF
uzJCutdq6K9xqzPYmJaCBZ0quhtfjUMQIeeHmEdfLgNEaUdmI/nHdp3MZSGyE5YYxOT/QQSXt4Pk
afqzXW9L3XLZchCKFFYsWfCSz2RO3rDnswRlgn39JdKLs1ibo+1wNnYb8UDw3egqtznMKV5HiuTD
fZAzbtdCjmYnNFgNJ+5wfuhYsZYASVheb2vd8IHMSiE2QcEQO4QQ0kBh4IOHzvZLqQxq6JMbk7qs
G9tltwOl85EtBT4QiCuRs8S08zwjE8cNUCL49ubpFwh0ALfYJM3vtkapiKt3UpUqPI3eBAKCI6mV
7ifJuHszJTtu2Y3VOuK61zIwxyK6M6TzimX6cd8eN620rnPydiaEpqK/6cvChc/Cw3N0m/w18qPP
/HeOiuDxUriGesbmYOtJxfpwNlXKjJcmHpb4v1IGyh+1zi0HIjyxEeOIMdQccf0PvI4SJmlkLO81
v6YheduB8XN3HVv7Hv0viWryzpZtQH7Iho5jqALTIGdNLwb1sBojx6fFZFwkNC1/trWaVrFq6938
ZUhAmPzZujl8qgwoALA+Zn9Jzhbj+ywnN+SdEE8Duad3KjhJpt4xFlTdhFCMwt4cyXUTlZR5/fM4
IW2GYesT2ff/Gz++Z65MPbIHM15r4yh5eVdIHQnz50yhLokbDtZB41K+vDiFoYnuBZnI/hTrbeXo
AEC3Ek87BYzbneIMkt5xj/Oh+Jr63cBjw7wRpuY1fw6n4ngOn68iqxgCCiiyWAt/TNqdTH7v4WG9
V1d+sgPcE+Z3n44zd8B5id8AcRSAXPqGDxDbQiAle5JrK6SEFawTt6bO1CiCz4V1DFcNHn5+T2+N
DobovTT3qUWx9o2a9HGyYcs+0Emt7jGTcxvxoxSpTCAqBmpA1Aa5a8O+pfBV8wcvw4xSCv5glwb/
Ew8+8d1ZLzzfs2At+JMf2+iflN0pKJf5ZG7sM9Na1UuYx+GVLAxbyHaM91+Q2P/p/4ZVoBPEpYO2
8fbvptIZWx3YI6cJnIfwjvjqgyIPlYsqnflpNiDAN3pKnqOVibSGZ5Guh9ofVt3O4BHlDTnw5sFA
IVlxcfoeNBdcG7xtpglpeviwQdcSfORmV8mjuhtfwyTSStnN1o6wp+znMmKE8VH5RUTRfkHVohu4
C19qauiyOBQZtJT8kJqnHWjDlTKI6GUiFg8GzEz4byfx5AHD08uT1ASyYyyeJ1MASEvV9PvFDg1N
sde0hNWww4pjNz1KJRT+XR7/uftAFwjr11TwROfyFNnn/HDVyYedzmlTPfNUy0rt7uojMqOwnvGh
i5o8oUT6I9jPEc8Ym2tzOD0q6UkIBMwGQwtcCrVQ49FL6WL0SzRoW8UtLn9+2czhPpjOjCuz3zGw
ZuljGX6//WSo31CFAGIz8vGvsv/E4bbpVp7IZJzRxYZ0xKag4tbKsNjSz9GEUSruIHtDOraHR0qb
omvpMqWwWdicfkafInj1f1gJIMCOeClIG5LMOb7LjE2IHPvMwRizrTJeHHu60607iSXU2a8guEjv
HFn4jIzcimO3QvveFykC8oGryO4uJ+SdWRzVZiQhK/SRnPNTwMr82y6bx0JwNpJ3CIJMHxzsnf3F
2a9IaT7cpP9Vq1sLDoMo0v/NozV3cq5h2EJs6i5LA8dXXGcmPK2BI2cPH3GfFKSMSKUa2jCFTiME
OA2McuiRhhbuHyt/MmwIYJjG9OVPjZt70t2XrvkvoHDjnPSvnUyaPyNwR8iPWoNtPPwigrOs6/KW
MPfjn/D72/mzJKqp4aYdsq9dUoqrt2wpljwqHU21rwDGg74rji/h//uqFet6qICPxRfafqupYl4L
v5vY3P/bSeSi1IXUBiolRI8kyyzJyIRV3Mk9B+moiIUTNTgKMlcoYjlrUVppZhrCIWcsgBDj6Mul
GFOSvfshSq3S1cOA7qgZmG5oK4mjzUn8hfsvBqKVHRy2/+A7oHOMVKENN3h12PlH7EClRh9ZjPpQ
NaU/4pIcOAgWT+9tFhAdzeUbONECbbqiKHBL0w5oiaKFsoZQIsR2z7cQHccr10vOla9IT6DOym/K
eUzUWlK+xLk3NWhl66jENXyE8VNS9aX2g2lh2x5k01IsOUu0dRJQSSfApvWmAEnbIoxI76mzzWLT
Scl3QTc/XOpiM+ClOgnlqPBACAjZB5WQILJkR7jWnubac4nloCxXyOnNDyBgI06GueWXJ7XmSmbZ
pp0vZ5CVgobcYAV+teo+FwqUl1SKTGjiHvWh3/Y8Rs11oMHd+8yx5garg+SLkzvXIyKyBs2gOKjD
TmxaEZxqz62yKzt/ENapZZUR8ZEBsYciawsw3d30Z9dd3RcVCsGhrewOYRf/4mpCJWB0BFjfeB30
hxo2KGbce+XfURiJsIO9N0BDq4kuJWiXMt3gB23qbki0rJPa2b794MQc/DNDia+O2meycB10qIen
4mQX6M458X5hYy46tnmklUGmZduAkaeBRnetvjPMo0nllzSt5ld5JBTj8UeIwoGycbr230Bvlbsq
+Bs9wJNFRnsSyC6YBabiO3497xfnw4xazZJyt5euInNa34ivTaSWGXhf+onoijL+1F4Gap77YY+9
i2K6J7KzaUzxiPtPoYvJaEU/9ezOjYb09SZUa3s0j/kY5bb91izUYu9Umoq1gryN9AA7ZrwdpNnc
sI/+O/fvwFqtDFaDvVtMW7nrOhzokEgI7Ke879Fk9VIzZS0WiRTtm1ggk+QyQ0IRPuKhYX3Lu7Qr
6Lbd6mvhGE5gkY75vpObA/zSeEnm/IAetW6dwWHzqtYhOl4xhebnwpx3Z/Qmg04PZV2+0zvUS4ZD
BGPOkT89n91R/1jKk1geBlSzQXBGZ8sPh8sREwdsys56jKNTEJh0hDROIlAzgdP0vIziQNVBNnxO
sSKEZDSzZx1F1WOJslrHydv51Qi3nqJkaRWgBQLKH4iuXL0PRtE/gl1K2E6FUeAU8G52WqPBsQpd
MIQ6Wi/5JxycI15tr8ULgqKHRPwbLBM3SjF55p0+B0Yh4aVMni/3I9T8ZY7RTyIB1Mgo+OXiwvlT
irDXREjeUsnG9MBuZhC7jDS9e72wHJxjqwKD7iqdcPaGuDgGY2JRrjXeC5dC5FbeoiWJgZOqrI0t
Rt6ZVg8DmbliO7CAQunWBI0CdJrKQEzhsoar1hlPrzIlC3lvWQRiDBPLqWHgmaZeFz1nhnQ64PRp
I+uxCqcDS1JihT0+Xh6/It9OKrnj4lUAeZkROKBb4T64xuRdz7t6aAv9sY89eeqJ5PoNBkc1itSW
PsBdQxaDvlFCwta86og2EpTLz6uuF3MPnUovZfHJACKkSKVoehEjNQxeowK9B9hq03VJU+PD18Kx
HjiO0ExB2KxUDpMHmtUtx4QwpMsWby9/TfN/dS8aeXtYfJb0/FVe4fnPEpsZJ2Vll2huZ4Xc2aXx
kiDDSTR8HtC6fozAvm6IxqpBePNUqWgGZ7918+5RR4GV3qAcoB/jdlVF24qAc6ehVtvL1VcNHY5C
4a1pkfjm0fKsRvog/kjgnRMAM3j8DJJHS3gZ/ZbMVGhetc+FGQsivVljW3aw81iQErnrpU7qvfU+
lozkEZUzrUaHYb+gEcAhNW793plxZ4n4/HA/DcQDLZ3w/sgeh7WGYsBqIk6JHyjXbfyMcPvbTTBU
Ci8O5fpedT1MfhlJJGIphEIhb9MS++QJGOw0KV0vFpmQcYj34wH0Mgd4TvHXbB+J+TSCtrrfPwu5
zOj7CZsB2NyrGtvprEsIxOSUXgwwwMIMXuCSgKRcBxN4l/ScIdYM3N5BzKsQCpLtnV+HwY6O+Ae5
C2N9AgP4ou4/aThNMNnn7zsrbp2TcUfeZfFSJuf/kBJUmyz85qENNvBYk9qbWvrSmXQPBm+bysg2
N1qTwvGTN/txFjYA/u33l4izAZM7SbdBlCtZGs96oN8jSa4pCcULkBQhcMzUr3cqFVJ1/g84UeAR
7zFXDReCc98On7iWPVor7yKhko8MFwf5ktp+Sx4Sr0oNhmG7ao3/Ph/ua0Us8FYYNrXY4Xy4jFSV
wI2gALWZN4uXo+MgQQjDdIn8DnYIZR0ELs9qyOcm2gGchdTDXDIieTG596ByKgD7ZoBF7Gj1bWrx
w0T8GtWQOdimxJRZjNOU49vesyneyrBPbGwrA43pd/iziNr04n0deQPeS1XmCabmxNJWg1mj1JaD
9TzF4WgQxbiSUOtgHk9Ca2lPmP0b6ClBhgDJSGUmvNLXP33oKkckXOSdqZzcxm9CRXzrcH/qbPcx
xya1RNBQxtbkuw0URjR48KTfP6jKEgb8DIUzlRl5hoVDr0ZUgwsUPNNHbRun4Ypg+2N2A/gdpRf8
vWCViFRyQxhqux6gwIOliz6/3TzqxtTb+3TG4Qi7ofzRshY4OwrhbwwdpzlLmXBISu3rYTKj/uxG
4C4vUCDM8dck8puAHLR0l1BYr2Ml98qZK3j0ze7HYwNn8N2LQpJ403OhrgzGF10r7wroNtSXI82u
qH2P+2jrdODNR3iBlP6R8DQuLJ3T678OvIIdL0pxP5G+nw5ZCbAm4DmZ3Yj5XBqQAVlKPkOoh/oq
OwVqA9hbF68Ruwji4M556aJsfgnX958mACvUJipcb15lvxSROYn9vSEB6T7FRr9yW30Ofj87NO3E
EzqxOOLPnD1jCQvavOciKgqaOo6M7bVMqEiiGaWJB1+5qPPMU0a6rOWuNzG9lzF9eRnvtew4SLkR
3z1C6/VqI1KEBndzogRKINysIWC2MK3DZ0dZk2SmzzQpEI9oN5bQ5rVloA6b0ChbAdhj2kjU2Hjy
+JzVn4uiPGypIWp6ngZ19ig++U9E7/jzKhR/qkJ2GyEADJX7rztRzfk5G8I7LolQ47ps5RfrS6RQ
MU19u/tm7JecJXcrv0HX/IICy7Iu0A3U6LBSwvt+TVP0/53fsHChvu7fruYVrjMOb08M2NHnhn1q
fVHRKDh5/SUmXAdNp2LiBviVDVKhMk/YGVlQ9IJYmn4rMZknrc3z+QO0YhD6tE/b6w8nF1umDrzO
YLAX1akEUTqJ8a6ank1/w5d/TS3sG4tlmQJMBOyR+8hy20SkyKCFaRDGVoZgiyadnOv0PDtmx57I
9113j4SCma9GfDO20ZjP567L1rJDtkNni3uXsmc6HgaI4f3HsmYJwehy5c2y/5FKQMM8eF3rBqDQ
kLIN2PbN3HPWiRHK/h4EOB/0eyL50bkNZx8NEYVmYyFubKmVpm+jWQLP4k/3xaUynlmqzVKpoaqY
0jqr1E746fqNt9lJt/sotM5eWgOpnZBCoKJ6tCO9ou8xM/AYmsQlTn5Pkb0phX5L7dRgaq83FRIe
GBMqolYXThhFZ3PLPdIqExcNyUvQpo4/n1xGvRmRUiqJ3ngSSIHH5yulYhjSzQzD+hOSlAndSq14
FigMLBgLbO+cAlj+LQ9OY4+y+MeWUc9CiLyq2to6nfyK/vYjKy8kFHeyx6rsRfWxNeQATQjlnP7h
OEQ+Rk0pZgNtsZBxFO4Uy6AaB08/df3nZK8jYhJDdIXp6du3geEMC3gPC7nDvX4RvYhq7QhHx4KD
OXdt6Z25BzAQ+wmh6CSSABkfP4nBN+lGkE5laOfrdzgBhLLxJRh2HWmX60MdSguSYV+XFldbyUKB
ZO+n6/4gHBsw09iTsbzFI4F7fbS+3uZlCRljd43AstV3QbQ9GRlcT0RqE10IBimH/TBYN2z22JMC
44pME7dUHsdLmOikn12abTZgGDnGjiTMzEWgW+QZMG3NPR8Sqp3tQtVIeFI3AyvdYNFdG7R5wgwN
IrWnlubiDrjX5y7hAhr2t722yfcFiGzLcRrAOHiSFN8iHEJnHv4tmtkmt352WV1pvvA2Sfyj8svJ
X94DrwK8D3MwCDGuyDQYAcpFqmnQ4Ru2D1rlDGjjLZVjUlHwFr5iE5oucnG+KhxT6MhhgdCSKAxP
b8a7KV7OgCtaOrEXOVjqaDpb35G2uH85J2Urx9q5RKFwz8RwmxDohcy1GuivStWCoPUZ88AG99UI
j0dgCQ3ls5AL4nu6znBuT5sE8XOunqFDVox2YDtwrR9RiUpIJwD4MYgZ+UA7q71Dy9h+jM7zHvBo
IRrbyFEb2lM+ByDcCD4tFhyRz2jbQlP9FdgKOhCRE76uZsuhiv3GOFXnvM/QN1uLz9soXXdnyRf9
vGmeAW2BPtyfhxJ/wdlheZnz1ub995bUfhoX9iNtuFeADYkpPWLXbblWHCHRSdtjzcSEppLef2Io
pWjPYBEls4kGD8JxP8lKplKCmBOeR1xb8HUXtWFGitiouQ139K+daDiLSXbAq8KSCuPGvsbbLGM2
rppHSWFh5ingFcbCFprudJxXECBe6dkzGVo0PqxX5KfLxIwk0i9RYfyEsNntq4T6U7EvxuhMtq5Y
fZAfXSz2VMyje0oXoVHdfp+qHoGx2FtRGfkD4k5PtzjEQse5w1aqMlDKAnLE9uxcpGOXoxofgYmE
dgNOBi8xCDLD1B8el0YkfaTwlugWsmTSw7PH9cqB2DwDAWOjL1vf+v5XFFXazhFUo+r5MJBxgQi1
WMHLX4mV/7oEuhZx0H0/y0IrqmxjDpdSNzjqYQjpaJcjFMQGgofSfgo+/7TmHFsLHAEeEer4o8aF
h9Sg9GzBeuiEoiUSt636LCI3qUeTPwWk3MSsSJ/ix1gFqffSB44mDu5v7a/A9QBDk57uriAC+rZo
ouqYsO3kQAwwmU45kFtKYk3UeTIK++q/IT4ZC/ugXnbVhmjMjmHipiGsBppegycYmmkBd1rSYl1u
sIarVBKAfxyQANXUrj6+YzaHsUmFV3pcDFj+fePwql1r2olSZ4cZCgkG70W5O5lsY9uNVnnc4t2Q
/7j/Gas7kYILEfvUXZXtJM3WajdBAy/qduCCLbWyB1YLaxExDZgMaEUKWSRWy78Y99iPCZUgJnTg
fXA1F+S4nA5cKAEFA0C8lSHH256G3sY16MRhyRUagRgnaXMmuMLqsW+eCvMCks0yb6JTstjQSbTE
C2Vh559ueTbkDqMf2G6I6W43wgsy49pCmoHQauOkjUTaH5HC1ZsicwxfNCpoEukcz9pz4xtIEU+l
ab1q60blr0rRJ9ZS0/Sknpm7TBZK4MbJWnLtm2uKvicysLldUebjDEN4ttdJGf7ZXA06gKSUjWuM
tUTQKIY5pC0IYkXk+hDdfNHBUXasZVh2OfK18NQSZwf8mwzDNokbAbTH67lbV7zi7eGFnL+XuHTV
GTj9oNfuqn6XD9e0GtxY0GDBEiXEFgxt5WsdlR6Cd5XDL1GEp6FwnO8Q46KXhaslCMjyp6eqnttX
v0o/Pv2j3DtGBObK/tmccAXJ3SzO87pEkhTkAscZTGERu7vZ0xNDfpeQbgAQQu0+zOYmFo9a6nUQ
rC5ChoT9z230Pn7y8Ke8UuhTR3+N3bs3qfdvcIZ9C032LCWTbNMEuuqsvfwcr+CNo24Kmxos6szZ
wo2+vS81PT/uBBe7pKPEMwEtJlbn6F3GgAQXmRdAFBcNuRqa1IfYEC7UALL4yuZqoJ9X4ASJFuS6
ux1tHEyvnViCpouOEQq1UAhmz4NoruB8V3Cx+Ou5Oi40dcYcHLCh4jTPOI45JKaK4CWDrCvPvn3u
32+W3Vyv9gm5BsQ12s2A+vK8vTig+ipHxvZ+w/FDdEHlQk/kM9Z/T2Bz7ka4T4ATFRZg4Bcwm9as
rHkBjsKJ9sd8pQ6sauzWXtgl8NQgvwdapz7Hw4xF4CRt+LnRzj2iq9CNgUfRb8rOwD9U25F5YUXV
h8aI88U0Z6lOtUS3IKtCa4bRAyzNEJgVUCxeHna2LH07QH8YRl1kk6QQWwygsCLTQSz/5mN1neBw
nhQ1emPrD7dqsPJsb0WWWA4Ay+/FGtF7F4lYqs1Nogx8J3Sok9sAZ6kA3q+gkgB+u0lyzjCQgDe0
LquSvx8/7y7HbKxMxqvf2rwjw66WWYRL9Uagv1TTgM5ZxT8Il/WcqX6cnKXzSQjRr0d6hAToTx0b
WtQhkB2y4us0HlEKtKXBiNQDCs7ieJgFlbukdkTIemZPVlzaPvLobjXpi0+XXrdLRis5VJN4US9d
7bNq7PcEbeqhTyLH7ma0w3g3YuEvgwcuE1kzwFMg3OfBCnFmzHBSahbsTocB6qGcUeCTZWOGOOBb
CszH1BgzKkHJgqmb2RQvofhvQc4q1Gzu6ByewKyBC11V3ItTXVCoJCsE8X7rTiPVY/J5TALS/idb
/UnbMtIoDQkJXQ3oKxjFRoQgC6HDzcEV02TZfEWW2lruJ/0Ubq6mwCCJ7GQhM6TdgQFX/c/S1jyq
4sxw74ejyJrczKMZFxq2FiXbrG5le1PwxCZiOkOVr0fcf3NqDpragIUEmjW1iQ9osMgxDkbzVPQ3
H4KQE/JwTFFT1nPNqGgrgurkh3q/VMv+W48p6gfh9rxV4oq8t46l2Xgg150fnmZbh78a6PmoLGZP
82eb34m58x4BRx7edWfEDTB2H106B20ORKOsdNCmRrOjA9UFAkPJv4Y6a0XgnX5rnZHPd7tKx5cT
o+BjChtH4YJoPvhvPd36fMYu6vubfjFgFbylkzLnZI6BiksoBU2Q1CMgNin+M2XTjlyv3P/tAYIJ
KDBYOi3WiWD1H3GQAv1hmyWTkztIIZ2ETX4Tnvu8P7Mn506tvRvMyNdM97J9Moc/mjYcTamc6CEk
2Kh/aKH23APg75ChLrWCR3Hzo9zGQV38ECzpdYlbbGOXFxhx/wiEAo8glSBuykRwbdj+Tihal2uQ
vco4sristqAApkL7PNm3nuzlUcMilkxP/sz0T28Iipvi8iIX3OXV+NNmci6YC/o0St01heu9WjdH
CVjBMydY8zjXe6KXwpA8NSZukPmONrZibOeCBHiRJuVGQsWHIKcTYV1uubGYPwHKNIHyfUK/2mD3
3BYKL+jG05oiSl4WCDc31ZJ/3gbOaM3jd2hS9YS8KDz8M3PPzUlyLRWxqjg7FxWHyscDkUS1UXjw
u2nRwtVJxNHJtDtGXR2suj/0UC4Z+iSHTiAxjC1slMDaWR1ukmPBHEJ92LESAAmmCclYJKv/4CIo
ZOQXAXLN0Yvn2uBAR3oAQvgCpTwYeMSdgc3Fui7SF705Nnx1lnT7SiNFV9NN4o2lFzGB3eohGbMg
AWyYvOL8YFlz7LoDklEi/UjFAHpUhntQWfj4sgaXjgWAZ9/sJ32/E+6F9BEJHux2bNK4E/7/DadR
Dv0jajtkj/8xE2G0fbpJ2Z1tV8f9sW9wJBpisWiiOMMXnLmXpsFNdMxKOEQ3g2m149qpt6Uxnouy
rC1JcqD4nUdhsUCTr+aPpcboyhE23rFuFzdHDiTGnmWRgRV4P+xPKk3/pwhC6GU3X+Ulhzos1A6/
BpV1YHGi+fLjl+j3ncVdF0IEoZ8RqzrODzkZB991dG22ZIU0lN+ax4GdWYshx+GTCE8fTQaJ9HVi
VVPJQzeiBRzVgk7wW2jnsJv18Dj/XharDJAsXP2HEr6d3YhETj9nYJhiunpVlj23RIgGKPQtM3Qv
PPbo7K+FXmEte9f5HcV4TTVOHX7gxQKLNTP/VhyOfUBMV7DV6RI4qr4rAS2Jn1NRLJ8n3oztxC3q
KuQMq3TV/TyXGI4JBjGxmQ/knuoLPA07GewG+mKvWr98VBAVz178x+j9nsNUKFnwRWD4UEvnp66p
8bLA1cjsQPtRn4pwIA3jSv7QhgwYd2bGjU+gyLlzRoKipAVSsaeF2uRTAyWHMy0jvCE83e+iAX24
1nYUGHDInwHHeGNyBQAltc0XqEKME5PxThAey6ctZHvzvNw6Z0GV1Wh9eYhjwdkvfsEktbkkpEqX
WsHCahJIyNAez92HWqjSmxDk6VkkQ+prhbccqMx6gqd7z+3NSo846Bn6C+5O8nZ+Mxdf86PMYn4X
V+zxSrjZOqMXm+KN+vBfWv9o4DL+sMG7OIVSJIQhJ58jep+BLz1W9V7L2Z2tO7DTfd3MU2RcDBGt
cdaNWYm0vz/gkRcljnbdl/ifXMibO4pQOHaQKGg1CIIIcUNI2v2kHyJ87U8BF0+DiC5vxLG8W+Hs
J/ammJKoYBlSCQiO/j6rrcBhdMvZaYiA+4pbqF43cNgoDa/vFO+7S8EsS+yPLwvdETT3JhvGOHIS
EwneFb2vp82yut1TqA8qWMPPA62hOYB0mfroavWE5ipPFVwkt19DDTZUfkaoPvT7JpvTQ1IPXsS5
5YcX4gnuY1gmn0lCVgoNCA62hveK3UTx5HIDhjNjsK2YUKnjHSMRss8XmlWV0inQ4zM6lj6+QyCw
ShxBZvQhbtWWUFaNJAUfsySmAV82LjRLHoCJZcMWlCi5ilyTlhe+TJIr3oMA+HN1VnRtXgcnMkU8
CgTU5ciXfMAuHKtq5RD24a8r2VWD+Ya2JXaLKPR7wx9Is5n08YaZLEBjYJxxaBgfe5rpOVQqoPFK
FgrFbO96Uoz6rx0aYriqUGDNr+/XbgG/QRTKKHg2Hj9JVc7Pyg54ZAojPR6mTVuUkqonjppnQGif
e33NMuAeWJX/b7O6IWMk9dWRlI73AGGkRsYE4r4oHIzAtVQNqJpJsGfSty17+xOvMYaFKsyGvtsW
W9GUOygtnCFPv/6UAJ1HbZ1p9jbPVWfuonAnkf9EDqr2iU30/mXveeK0BPFmrniZA5rYiicKDRj1
S31h3yuja9uQBe3YvNcP1Bz2HkQlD8tJobC6ZFn/TLycoT3ec3rIxe8DcyUXCAHS6cePo2PHQ3YH
fwt7vnEJ9OYJ6R/ca0gxgWNyQPpvh7jyYmqCmoNyDJZyXfdiWG4b23JTc0dv6YbSIb4kaEpBDERI
Q5Np+KgLNIMjdBB2DkdX0cMg6s0dlFV3cDXaUGLVvX0FwPlkiBR6iRMiFFh8ohRy61BR6IIaE3zM
r6FqS9kNqH/8TFE1Shmog8yOWFZwv/BujLLHXoGAkF+LIMqn5sZnfAYtzeCuueZ/tmn7O2XyBrVT
SpbRWuaZiiehKSCNtlb6IojG1Y8VbMpgfOAg5hTnRpSEOKL4oxQdqzrRyAyYZcAoeIp0pVOtaXsu
Ou953cg3f7h26XMT5DZ9TArbp4pfcLnfz4rnoMFG4hzPmenmB/SNFN79WbvcsS44iRtJXjJH1OUT
L91XJsdohgQa3SumWB5aqiEtJ0cDATMmmkva1qJ29guMblEjtq1Tl8SStdIFiWGmLV4b4AkI44nJ
8YGBV1TdeQe61Sp4i14Ox6vWjQQiNaRG3TtvmDnttqDQrEqql+In5YgY1hkOs5EcQcKeQ7jzM+ds
mHzCFvHGORrv6e3E9MBTDSDMouKYhRuHpDRIV9a+cMS0/BdgZh6JKWTeS3TVoO4LpkNDH7eOVJ2t
nPNFCK442e12ooaZKVgcUOidnyeWeYMPBMMTwRgw80EUl9ND8Yb1/R6TTytPhcTAwt5dWY2UNt2F
KQC1tmTCtr5rk7wY+wcabemXaYdiLc1bk5Vf/JRPatH/v2bwrUR0IFlM4+ikUDcVWpOrAp3BtVzs
KuTu6uZTqcrWnkLD4koT8lxRTDRicj1BcGSz1n3oPNLmq/VgkONs2KBHEfKnMyq9yerCX23jctLT
XVtDwmJHuWqRNt+yME8B4jFr9eNRuM8/rNWp+KjT6xkeJZ2T9wcFBASrzGsaK6qD6Xn7ox8cKIjd
YSjIyVgY6RKyEn0HSWU/+tfJQg0jvxHa3NWa60+3El22JVa9kBElwrPglkAmWdk4qxEFxscGf7ew
cWpFeHymswn/pBFcrVlfZBxzEPwzk5D7S1J0yDD2JT+Z7L/u+8MLobN8dVbLy0wz7H1yigpPkGRt
GWQCNAb0AgzWJiCCHr35s/XefQXLKxc8zqcQekqlv4s3eGeR/+5YlDJhdNRKhToT6Yc3EqpeD4i8
9inWwoz4MYJ49C6/SVVhSoNZ/pxX+Nm5mfdmFqwrk+l1BVgZ/NDaylnGBx2MGeKpH4OP04rqWed0
OrebEoLgUceapUpIKcbDEVLS2Ew/ftgDfiiRqMiIKtq3FQ0SXGXE28CxjGjV2R1FbHC0b4xDINzc
iD/Pz0V78pFoXdRot6hCzWAanwewwoxQ+q0JVlXUqwAmsOaCoWRJ3QDAvK0yjsvUyRJk8s1YdSsU
D4AfLLI/1KRFTvbcP6S961hjzqtra92ZjVn0wMZdVRN6lR11bIZaO3XujCEmYBYxF+tpSehvUoBG
pvM50tWKTwo8w2WdLnAiyyNtCe95r/9mIeA5FUDlomew6crBq8KIkg/rwpYVofVRMQ1TfvQromZ4
7pixaUzpWZvQZw3oLDoMGZ/nZRa2JKK4pisytqyxRUKTvKfhzk5UKvL6qJPGQEkr3vfTEGZewvXX
fO/OC9XUlAshfxYkGuaRbCCqgisT/0jjUzo8bqGbphWfSZeQUvVDqxDs2ApzszF6iWqNX2+Xzu29
hfh67p/2EnM7g8gDXJyYz8oAyXBOkN2ynmZzCzaQPF4APuQ2Vqugi2wA+yABrmUxoNtenJEuceJ5
3CAJaSsxZ7GmInTCvPSZfTCnqPkVMKMruFkP9a+nhiDqvxvbHn3H7FpdPrz/w7Fhx7ocMYaN8VV4
/LlXxr04O+srSIcB11SKQz1XQHQzOfKEg7xO7fsQHXBWUgBuNZc03XNB+7Lh0LeexVjPALwDDgJp
b6dSAb9btGnGqtYhCB6ejBdDntO041VD1EvDyPWkmuoDD1GaqP+qsV9EIQ+xfyoumxv3+B+bGoP4
NPzlEMNtwY9MNTNpuE36Pfy0RQVRvykH1BbK1CKRvUX2BpIkDg5w6NhMcYryGGDzSQIOR+gLOVLj
Wr+wJZcQ/M+eZgcvLFMbZJGPTLzIJixk3LtylPZUGT/Y6afzXtbCIruI1CBuudA7UWsy/wDIlMwp
LNAkxT3a2kVK4eAOLgVr0E92cYLs+yNAhw1FGHSKr6IyBmJ8oNdcO5nKB92YPSzLqSAey6KE/Qhv
j+EejyJzG4n5Nq2BhDmm8H71kV6lXn4lg+kaQYwIDJCzOZkt9+JXZZsFgycIcWOZhH2hYw98tY3p
z/xqJVU4k1MCOuQMt7L/wJFCo2s1glbCLs3MLGdKicqpBF4SK6FIwluJZ+QKKXZo08ulDqiZ0e6j
KvBexEgNZcanQXcYEUnfFAjqFE2EfxPJsANJ5F3eQk8oi02WYCC3db7Fj7SQWRG5meM7unnMxR0O
5SjGqZzNH7D7gbwplSJtB1Rct50z7FFY2d7UlSnxAyCR+h5ruLlbHJIM8QVYEh80/uZp/bMcyufh
0ZHQa03C90qqBe9PLMdDG/SbG5Iq09UgUdgrHbLNmrLD9o5iVx6l9ydmmu4BmT0h2oc2yhvxddDi
OkSwrL45QnBZZ0Kypgcc2bjPeixBt1bjqSqLKNp+P3XbnLjjn48SXqF6h1Nal/6smbi+5NUAkQPk
2Mn2El4p0xlWRfEpwKPOkrTOkVRB5x86aJFwW8wzncYc9pzAf1A2EAG07dcHZ7bi3HDInDyWptSk
ulin0nl393XQOtxKRSfUoIi0b1tTXYIHKm/AIavZbTWEkX3i9UmqL5T2GGmvZw43Nzi/Il0ZIPbw
1QOl68Lwyrf07da1kPgQgBqA0O1RpbBIt1SaIwHWfE50ZiQIhA6TuOLFvXfQSb/JwYxlk/bxS31y
HXKRJeATe/EjMXyQjnBC2ESOeziqFn5AWiUIVr5tp8d9WbKVbjBa59xOiQfmNIEsqoSr1Hb+xqe7
DgodqHwTopMAANofHVVNaDEYpq+thFxzWNRBtww9cJMPqqaBzzuUW6p2pAAU9ZCckEPcnIfivkat
KHAfnc8kID7bnf0C8ltp3XcAcwGtRGquv/pzWvDvQucOcg4nvuw9liqk07Fx9wOueswcFw3BJ8B5
kfZuhM8Bh7t8cMLdimIPw1QFtu2F1fd1ixfvul0KnNDqT9WCCnVmtCPl0jwCTo7mx/E+eygFIefT
xmc4CSsxBGLzMPHS1EveMi3stma0Lp5+gU5ZZCxkdLkjJhxZUU2Knuq2e5zlRP+hpxajbSWpxW+e
+bTz4QrFnVtxqi4hwIXx/rKMIBJnUy4HVZICslhLotVqA8r1lBB4I+cb43auCfwxp5aEn4Y+kyJ2
M2BZqth4V7mG/lxPs+OmKYgoa/Ad338ny6hL1FMswwkSiBVXYly0YO8Bs+eLJcEmQifsNYkJrLcG
PgDFxQ4UqdYIchYgxTVeJMAh+XLGm6g57e6NgvIJRRm//T16M2euE01r/dEUrV5J0Xr6nZ/oTZNz
jzCiiY4ms1hFylB5n3T7cOM6asIB+ObPyxkLBGqZd3EjVwxtJ2agw3S82JM/M7vFrwj/VwEwtHwg
LLGufWJ0p8BjEmNPghMQ9yNAgf7vCd8SCdtqao9lWvPR4CTCk3alWLzwzAqrjxJTxhqj8XDL5gpO
4ubPKjuC5VvL9XKpx9hhQXJ7czy73de047bmLAei96IBJT3nH0Fw2hbI8CPNqeBJZU+SkRKp6P2V
lq9BrS+GQRvh6sjFwNL8STO56hVV4UMF/uNby+uE+LfBpMTRK1jh8clCjKbQkPJThBG3elksZiXY
tvXj5PA8+NOmN89IQmN/1JZwAQztrwGlf7+SLN6EuLGm0bmlUaGsG/VIEPEnvpZ3l+tbFehchMm+
O94p+RJNfFo8XmFu3oh6S3x5grkG0qHehwXZi2e8kerzet9z6iK1b5/144FbkK/XyAbHMrS6kdwN
A2mSvAjvd7462i2fFyPzrdCycdt4CyDwJiiik/PsXCHjBpT13n+NcQ4euMUHzIQ0agi6FRyNrpzD
WvHjudElnVzPJRf2d5RrNJvVT2XdOJ4pneBUrTNGg+3V3O1UGQgvpykS+KGeK7HyDgW1ocy7qYe3
SOKD8C+HsRt16U6Z5M137oDwZsZKGi+MqUm6zF/+pcGzdtdOXFoy9OZVnlyVOvpYEQRBTJtv8VNO
SP6os3LXmLy8hORx61JkEfjgdkvqGpGFoKNjsHUZZr36LN/whEy90RpgFWgHO9ehDregwW/9+CFY
seNysutqmMiB7nZrh/fZKRo7E1WlE204TgQQJCv+07LqvokrvDhBsMTOYbK9uCdRwPJlke8E7ZO+
42ff1ihAMz1iE/RX6qvk+TXOPTK5mtAspZ74xytFT0XecCPQ4UfbgHMDWO3n9DinGKTVTgkKt6rG
8SO4S3QMwCRZe+QZ6yU13gxU13CSqXhMn6dU5YWSkwq/Q4+NEo8o8rjhKUL5SqelfR3mPEjLpFOk
aon1rheJZsirGichYMGYHjWwWuRVwTyxSzCGK9hSAmHnWQV3RZoTa/+JG1KPlLaDsYo+9RNwhjPT
xtpU9jH/V394okgLCP1Db7b/Z9OWYLFN+EnxVYOcAaJ3t6bja/CDXfN9SYZ9P/mjJMoi5p/BB4Ev
3SSaqR551dnee4EsUSqvumA+BngwccQkKSDAxc96ZtJmxT4qM4NEfrdsPJYLq3G8jRuYfo9xKp5c
HghJ4FU3usd4H+0tkjFDPFsdBuo/b1X4j15zFJxOm1PZC/VAfE3zUXrWNVvyrTdIDSo2IByHdbfO
e6EQYvXHRgdbeJkCddiEGlUKWJrIc9zFTRFd/xBzwhZpmUJRIGN9gb8cHeo/0DlJyGUpu+8rJgEU
Ks9p9/XQ0bwx14BWCcmQ/iwU9jW8UpS9akFPBcu6stMpLRuCQ+TRSjImff4OR7x91etEIPoJ4B9W
gtFNErxKWw5ISOqaokMp6sRajEq01FGFS80vag+Ntfm9pu/WF18xauOrEwgzwZ8RJ9sFQuCiV0oq
o5ZGuouNPgj7l6xD4J2DHG6MmfS4s99QjmiAISWygH4epPDM+wMsnukHoG6kbARWnbeXfgDj5C4j
bPgE4nxp73OlRJDCvwV93RKbYDttsEND/a0HBHetmPhLfD5cag2TFNMMsoXf1y574nw21+IrHIDm
6jge1YOjGHwUKI/gH/bzP0Mi15srx4W67pHjjd6A7+/UV6ABqh+R7pcP16Hnq5YScbShX13Pft5M
JSgM/nXQPOZ0tRcK1wKjD08u8X/8+mNjHrwC9qP25P1LPP0PDdmNSn3MbC6zOKzsEVJBFFUiVUAZ
WchxJRNt8FH+Tq96i0drjqte8pGHQIaoyLWeVVRoZ6cmw+Bx2BY7Mp49+Obb2WTyDhadZrdIdYo6
DUcaV83hLaA0yNMlMKaBUfYXxH4SI8kMQLk87yee3vqRhrtBwpi1kLT7I2JoySdpvXEDJkB0UWrM
fwtucVeqpUH5eZ0zwqGoKyUQFkZ76hXe2TzHJ/WgDZhyh1mvOToYCCrrn2DgITmNcsIxfuRpJpkd
tIFyOARzH1f62Vh5cRDmDpkepHCAYWYOK7xSu6PNhmenNacq5FXUtCpfVVmlKOkYz8hy7xyD3eTO
6GdXXz0mYbOzrdFGROLnq+V5zcU+bHLJ0eZnsMo/QujLXVC0UL/LTZUN4hoflY8CwKUK8x3qPnrO
3WpvMomBKTUuza5gJvijmJphRjd4pWfkxm/+iKdOvEnIFirLCyfV6icc7eLnFZsK/lJBhjLwKdGe
MMg1ZGa9wdolfvAIES5a4O5XeNlJ0y+llKEk8ztKpRlAD7XOSblI0ndGtUe0BVs3uT0Lsc6oIqvp
5G07wkkqenNuxJm2LTX+bHrb9J3PthFqp5ZhP9Byn+yxHUqbs/a3oKKcOwCmPvtKlXn0orR3dAnR
D96szuyWP8QH5PCPgK4hsJsnWIIDIvCc9XrbqOaRLSg4U/qghSUqXyOosR2TJz6v+klEd+1YbL7g
HvaB4xddIorN379z1CjafwQEpxESzfgZVbZB48JZZYIqzeZYtEcG9ji1rsAWsCQnACBe3VTWI/OH
6wbVpgXbgol8a99NY5vhfwQkP7BSR93gMI+VH0/xO5XtMJR1ehcMgD79vJbI/lu69QIKyd4I2ANH
IRIVH9Zw2hzuUgLcbEw4Aj7VJvVfkAN0gPrLFjdMqw3oupi7oRZ2XYKj76TuRnMWSejKrXrjctKw
55LzhTKT8m5rBkA1rM3lhQYyRmY0zh0HSTINJcG6DC9ITCpjwMrAvOGJlAE4O19ApTV327eMF4Y4
qumTnYQkCBTXXWsJfRrM9dKPTGBXPNu3ApA270Exmd3cn3q2b/nGheSwJXo13wgIAaIvnRcWbh69
m9cUyitCoXt37pQ/VzQ2FiYkQI0YyjXR8jEDJlrfCUdhJ1pk5XLyk16yIKBWPMYmGC2s+ErOX76X
S9heutsGx0v9p3woRqXEF0DSwvmAMQ47z7UX21g/ke/vJWGNn7uY7c8eDg7UFDC2JNOsmuLEzxSX
pCPBRrcuEIytOg/fVcc7mD+WHAg51es7Nypg+Kbm783KLMr6t5HIkM3z5zEHeUyJC7tMfQS6C4WW
Kv6eaaLogeFgsDE73X/76dmDTZWUtHaJRJ7OC6C5zmepSWXE8Cw72M763UfQog2e9CbaXxWJUsjx
rX1zHoJIOYb4wjTW1+/4T0bXGCxYHy/8z3mcau8y8p7Kpr0FVZlXZAVMpnvImK6YxlcEomojtMHV
6hqU9i/erA3veA3z75ppf1I3RFArfLPVkpgxWFcn87YnzVE5XLfBMUX7DIK0GByF3UJyC8bGulOV
+MG2BJSc1XvD93k68jl8ki+bbXbsYS/8qdsH4+0g8egtcf40KFuajJNYUSEgsWtZ6XPl5gXLhG36
IU5BE1xqwpJIgTy94qiVY69vOgJquRNjW8XBUg9MD8dECzMb1xV4xpRHi4E7jvoxcAP5qmdBKgK0
phhG6agxQ5qaODSPRjUqHA+PPto38+9TtXIV0W7mrmxJ+0fsoXtyvYFKpHagHmpMgQnhYbJlwk3B
sJxf5H9yiAPANlk6m1HthX/yu49jCXhQuSefjr/hDm3t6gx+3GoMMogUw9Vxmx1axPJTIT1J+GPH
l9ud1qzEmhGOyTVMMeHV4u1z8Hs3SBfyZh1lLpmoEM7cJ228V4OLo9ZiWZdMmdmqzDvAgfsEi4fT
Vq6cnkDxFKVHaBxwh6yMLDxmJ31rWcoRyhVs2pfnelyIDLKPS2QYudgug+iC+5IlppG8S/OAJMZw
Utx9BVdzAMbtgLCpYfCye9n+wEp7YoKBZOQwSZMxb3dTvqjyR0OQpUZQ9JrOSuqhuXIM0v2N+t9P
owIipzLmfuj5ddXiMblKj9prP6PpatXBWCfDi3EUcyQpErQgBfv1JFW6s5+hIZHoWnMaXRvPB3wC
7i4vxX+Ckjq4ea5lHeggq8khw/fMD9KitW+7cbaMXAJ90QvQBG27Vx61uu1cGCuASDlLHNQY9NX3
pApCH+sdDk4vu+9MaByxRINO2L4FNNrfscBI1Th1R4CLnLx92NHnt1p4+HK0EidoSxJG9MIbTIa0
r91YwYk705VA5+2rxOON7c/Ue3K02tq1u/4cvdH28PMF2gttWmREB9dRZMusVV2Tqa/UJOfyJvVZ
vCmNlX7wZcsoYhlI7aeAvzPVpAgNfoXvhJ7XmdwqEpt8yYLtVUWStT806l76n1HBSUSHcsHI+++T
6VnuVo0ae//VAqYLSr6WFxwbDDMl6WKH/YxuYrS7BT8TaSoT1xckoQbkmyLadjS4H3GizGbgwA3L
V6+qoGPIUuHX+Iv9yy/2xp11SMXU/TWoB8lPgJzIAhBm/HvxiXbzKxigl/4r9bu0O0tR6DKPiJtC
Pg8rLB8mdgNAO4MDpFJP1achP0qNQwVEm5GHHcAh3wAgtFN1+LSUaR+ftZyNXL3lqLWyrMAepBZ2
nnX2J9q0BmxY/VGUd2GstddenHOnLcfpQ5PL/JoDLYd8aJub8FLNFlCyabeZfenZtf2K7JoiawKN
Ai1JBBYuGTa3MnvzIH5D5vIgn0VMjxmZcvaxGMYDhIyHlKBkxtIgU3X8ZbHsReq1fSb3YIyVE391
5RSL4KYSz7Ccj/nPlRKSOQe3AnEzM+QQlmiUpvBeDOl+yDCeI5xk+WOxN3g0bY6ZJLQLBtVX0+Lu
+h5h2fELDSWR/3nNa0IjLeP2JqcGZZczdgTbOLuRY/xjhHEO17gFdCdhF8tF6q4gzMKvGHfFHT0x
Tr5pHe7jJU2GlJsO9wc4BDdeKpv2E6X6cbvstcWGIT1JOi0jpyOxJgyzsjtUCTVSQkij/oJO1+op
Ig0I8z1iyrvsgNuQmfBbRPDa+qtu9WRwejzpnICTIx4GFtQV6Y0uY0GiMXu4DC9IWhEmxn7aC0yj
H92BSPtc7ljNnUCAhjwufM2R3LQurKytcfq+GJkCAWqGvEy8H8lzxO5EBUanjtb+OLPSQNT9nwnO
0Ebbf0pfAT3iM8HDizfXg7rs3F6hDCG8HVJtuYGcgQ+DTTTjCa3ZdenPv4DzsYHMR5mrZWZIw6Z0
S5DaShrDotkFjVzDqppIygUhEYWczxucgl7Tw2c2VuvLeDLPHqlSMMTwygo3BZDIc4ENGo/w3eLd
g/NI8wNeCMgRXtRwlLq55EDUE/tjb0/uTn4tJWXqyaxc2B5dejF5Kb4JMCw7O2ttwCO7OHKW2c0f
8lRo0XDYFV9+lcIeEWFjD3E6TbWHENCH++M86IaWrVEJY28TiDG5Rm63nVpd9eNv3oq6Uo3cbLOq
4BfWgjJ4HMxFz/UzsBfzT6yzonj3jZzE3xV76PeLkEEfVB5kNoB1asb84RL5qyBtfPDEOHI+ZfzI
CchYPiBxKRqnsmLzSa5mY8Mo8Ye6ANebG5kSNCPezlW2ZuuyARuep7oN2J0jta2jiPS4c1mB7glm
KpO6jLVI4pXLnFoXpQSSqLiwFfPMxFUjyavXPHLmx+CXEEPSO+dPGIVsE4RhT1YtIlxK5pYbxNVY
mcAylVJpOeSaktrPm0zl1h/UEIzZgqGafSYemHEwEYNaQ0bJV50jGThBLcnBiIDLfPrL9CxKPhXu
Q9Qb4B19WqDPs2AZJkXvZlJTYzV2KAM8ql/3ek0g/aX9pk0vHI1S5pRDjDV6dFI8l8M/cJ19/n48
81u1HJAXErV8u7LHHJ5iK6B0SY+roKx7M4lR/AVemCRPzLtqGu0jLTyydiJZQ07LgxLZP+GdIYDV
ViHJvOE10yp9uJVtvmCYa5zNG8JHLx9r1AvYavZ+E3ZsPWcDbvaH4zH2pMBcZ08vVCCKliYvVdt8
n9tfJPJbTO+YqEN6btn1P/0Kqib4P6ZP0KDfXL1ST0lc4/8jYCRMU5UZYwbGYw5RbsWLRcK1veGr
IdNh+FuHc0kA3Cv8WLVvrjZ0OGkL1qYwDed5M9sytqITKI4WtLkTdLeuiZ2GHDctmsKedEnsrCZB
6DCVEyEoD7Awg62zjG63p3fLMXPRGhJfOgWkvKE6g4ba29/ebSWwjkEG+eYpIJCNhE/94ZZiqIv+
Xn4ttIhVsCOf4Tw2DMXt34RyRn6LFm1ATjwqojI/WcS6K7a8ne0u2BwvUM08Sf/j1XOLUbqkRwiM
DyyrBAFpIqhKBjFgQMQgj7C17TthQhQNk6pA6WmxThIqt5n6wmt5HZzTOJuw1CuT5M3Y9qhCijVY
5cyhcRhQaIskaDXJcSvL8/c/NGXlwH8pJujJAAs1TZGhx/Vx10OeKYkzDeXzkRXLm9ajg8wXL+Y7
y5+J8IcA9j64xZiuiUk0PJgB5jpfKjNeuY0MJeDbyyMk5/XAEjeprJCDzQhwqHjxXpn/x7D9P3ZI
M7LnFL9ILSHXPNziGWa0TtRtcF7adCaJ7BPNI/gaoOAzfDQVfcv62iSPNo3F0RPt1hH7SvJ/ad3r
ZpIF7YuHMS+zzFP22MB2IEE/7SwLzHFWTAJAu7mExG0Oz2B3xAd/GkE3lOSzJowr5dDlpix4UlFA
SOMTNV3Jt8MYPF9viHhL+QUhd5e/IOdDIS9kYM4gYhyA8+PYSj0ex27UcGEZcsJr9FuQCopOI6d2
8kqC5RJ14kXdp1kxog6fROFJt11gPTZeJeS/0gPL5cmrrPTeUn0PqTFFeCyqKAcJNgYyfbPU7kqg
8iNCgD5uJeTawmI+bOeYCHEz1LWPlTZcYRk9HpxXFumcVtY3cuHT5cDmF06pYaMcMj6vQc/wZhQd
a7EUjvDg6hBiiutDhwDDnZdtaLlFOEFsd8C33TsgY2Vw4aaX65rH96XHsxy1wwat8hdfYiPyUGh6
UGhhXsN8Y9u0moQCaNYTIHXjW17E2n4NATA2NwmB0zl7+JkO0HFKvj6CUyA7Bm3dkg8OX131H0fu
80KPVm3N9ryzeE2CUfjiCJpmAFFR49zG3UlX+qwrEgfB1g46rgMOVDb6Ko/UjYBsOnnUwrjnogkA
f6IhzLioW8pEI41XOeFjaiIcoVifcr7f1efRmlGy/1p9/JLMYlRASUvO2JiPG2IoWFr93iFUNdJo
IbgZA5JcFn7k5ZnFVQnjsiUUY57TwXjpbNuY8cEA4X6PePguf6ktal2xLg5sHCcOw5w6pMpX2aH4
+7w3t83K8jPr+yIDoEmjJ83xIX2eeLXO1weSAEfl5udh7IC2/h2EwpzxltdLmBnSJRfbccqBfhNA
fTRP1ZylzuM/ByqRZrJZfjFN+TNk3NWHgaJUCOVWYj612zwIMDYk8kZOHJWd3J4LgI0tTtc57mAa
p2yoKouwkfTkloWGHYiP1eW+fQd+lbkkgZeT8we80d7OwT+09bJQpBqJc4AMzBtur6AuMBvucXaz
DmGqXQNosU6PpMWkzBZnOPsh3afk2vMZuITknhtV1Cv5YXjiHG+OZya6KUForSJ5aJzEWdJQmlVv
Ig/ScpyxhCLBVHy6YXQymUPg4oYzbqkVkvIXGQJ6/fASb2zSAONoBBjDE83aLYmwg7LcmPjE4mWs
OSlC6nrftqOaBxmrdqMgXpbDgSFgSZI3HJfmc6veJTTmoqeskx4uVBmp1ae91Tpm1PjWxhAaYCh3
Wlq+3pdoZ+Lm6TaptbGuZiqBq5kcN+rpw9XbW7BzcbWmwAQ6SBFcgjfc1HtOO6/LagKgKXz2C/IB
phSl+4+77GyKGKCpi9Xu/KbGd3shtRoz6D3iIAT2E01Q4uA0kN70/hB3r4+mB8mRsBoI0Kspd2R4
rsDeVDMsoVbSL1d/aLZxNYf55jFgUSY0iCcoB4fG/4jVuflpcsF1cFkUi+eA/rBBqMVm4ehu9KIl
0AOxOAR4zg+lfhojHGPHM01dFsVp/2Tydsjvn5wfLjWkrO1SDwGZOydVe3YDXTWYQND0cJaUrebK
R06xpk6s7nSaFQZlwwHd3/+KRTch/PdguHOkjrJba77OXbxSFzmG6aATEDQrc1KR/LyDOW5qCzdV
d94lQclO2DYBAJo2SJl36B+4qy+OmK+XXeTWYURLM75TVNkRCbNdmxlffKrL1qaGxY+c/YwJr95G
YjiRCQYrjqE8uf1rm4xlLGxae4Pc7Py8rlXQGwCLKzOK9mQRsjwPZ3tBs+KriLe233Dv7Bp5GMt7
FCKi+dfsAukQXkXYpqbdVEnb9/M55SM9s/89uuwceoEUZIMkbVo18e8s429ITAsBC92H7DNey3EV
DtsmMZ2lk9A30M8F9uP575sVeGZvvF/P/Xc6AUd3q40+euc0YKbu4jQYClrqy11tAUwTOZ07KsEy
SwaCMh8SBTFDMP5AhXZPBdM+fjpp9GtAmgWn2Mx4qG9GYp4QlC2wjB3+EhqgLe7+SFclqL8LiXHd
BizdbN0PE9jVIt06xwVYlmMJM2zj+bYDNRel4ltMRoh0G8uRJKMgX52i6UEs6zHmy8scBpPvrmdk
M86P32IZQU+TuRVQFujV7ko14h/ccGwjXrmuUZlAEG0TeyrBgbhvlnt6USVDWgTAPoyrm+K/ybe1
Be3R56o/Tl6bRWCIGodeX3uZr3zj2tASnLAmbRtItJKe6G6C62qUjYloonaNAwEsCb80QbWcuHP5
hBv6+I4e1X7o6iX53oWx6jkrPonHyRefFhKblw+l0ms6R1aRrA8padXswY5LCLj7OydkPvt0WXro
x5WBqbxrCqAxArw+56OwVLAuf1ysvdxbKdZvqHUj/Ab/EXs3wr8UnzXoU211fD2XkU3GjarpLI9n
ANZ+pSblrgJrCYVVpaJAy3zcOe1WPjL/AuoW1AWcBhPmdVeF6vT9WoT0o6gzoDz6Et4IFl8t9KwC
4O/XsYClH4/QsWpKJ1wtYcmeE474Oz380Bkz2jOWfBqvDjTfnvxqVNTvqO+6voJ719Q1hujzJZWG
wnU+P25tErDkZFyW1AjFmhpBIqQT1BNWxtEPo9wXVk8kIUDMi5bmY1s2j1eRFnl9vagyCOJlFJgn
X6HZ6iiQHapRmsTFeAEO2KRhasKjriAHVpkt/epkWJ8qMt05/MahFak6AUrmBvF0aOI3hlFYiY2y
VSNA/uu9tPoavfL+qxefeEhBSZ+/9eVswOd3WWQ8HZYLXfLWMmYIZmFQGBaVeZDlryPzjkkUkEVf
O5XoBXKBXTN6Qmnsz1RuDGjV5OnzoytcoToUl2m8ztRTbKs1GVPR7unCkN86tm8XbBB+GVF0x1Nv
Byu4hBD/1ix7o5QB0dUairvmStfLu29t0dY+iSlHLFB27dAkGthlVo1LAXK/OuwMQbXW8Ekimdf2
tw94CyMP5MoklGM50IoV/KWmRFafmDEIRkb+Bmo6lj+5KBAeC9XzykuD1m43tSyO7lNd/VrReWDU
F2qoOwzGgJ1HAhOakqa+BEfvi7msbb3qqdLIa7YO86wr3ZC1zAv2TZBZf6jx0oV+cHqm9JJJxLOP
6StWN0XX3RcBKWoWn12qUkn0054tCzzRBgnCXCIw2pNgoJAqN8Qkkq4l6RXO8enHwLApTyhgSGf/
hKLH5BK6nVlTOrHUYDRXfjpO04/khiZoYwI96kOCNuV6qhXsN/iLkSAMkvpjlP9/uGGpe/KSuM0f
iFLtfpiM+5fNvpnx2LVLwF2BfpY5BBLpmj/JZtfuRmzQ0vLhmHARQQG5KOObBGy0+pT6yhCsf/TB
+dHOwucoUKZt5lxGqJdOaFvPKhwN9lJdeBlIDzJIrbe9NBnQgqf3Gazup7O3PzVDFKQaPi9ZRDQ9
tRfhHFVUsh/DwTCnbTGPK87lRHkod+bDUVVZaQlB2wrWfxbQ4q64CXBjS/1SF5jIawT2BTdSsmet
N4+jx1q5wotp3AYiK5kYPvpLzrHB6DEEYCcpWw5Fk35LdvwZZETv32ZYlFwF7dCsw5ympnEoKltg
tvNHQKT+FggDHj9GGX2CjhJWNdRlPCv4xhFao2OLAunTbf6nxg0LtA4sqLSIKllxAjkauvJYFQrw
7ao4l8QMWMFK4Ozwz+4uADZDanbPVmeuAubVTNMHLcnC+A5KRA7yRkIJuoLJPHF6Ox0prudxrYzN
uX/cLkqk43HchE0+1hGs/Njh4LBoYzExctrcsPBWYLKkZ/dMMC2zYeoUZWZbGVma11jrofLWM6/D
Edoy/DIE/bP8oEMLe0sfA1USMSGfDyILlv2VANy/7QBJiBmYf6jffymx7AyF/riQdxN+KIHENmjd
ye5ODt46lwtN7Sy6n5/nQgxtuy3beTFqczd6Ftrled3XZf5BEbK4LcFBv8YihpeuhPdTbLBi6Cf2
K3rt7eJjm0JsAUGxwLhxWiupUCVymLvzbzG754Gn6y5DPYDrjuHcGfeekJjR/pAOj68lr9TbKs2S
OBHI4j8cIbpTEiyQlTn5doiyd9DnjFWYqM8ce7bNpa1G6blW+APfX5egJYyax80clNqwLPfzWyu0
1JPr7XzbB5HWF+LR7jGiOom860zjthQ5bicVqjeJc1IliX/j6IFQ7kor23i1jB3kmklvLPASzHHy
7Nl2B0DC61FtO4uyz0aXjmcHdftOYqChk9dS+VSD/O+to4sbcqqMZ7UU5jYZJ7TzE+FlBI4KUO81
5FNVVs5D/juGFKHtt0ySX5ETdIBk2HdikRCvBQWiwNeyEUIBusVAzKGKmqmpchSgr/KyU0nbQUpI
KBXea0PwLeJwhwtyUcAjFqQQIbIBeoYumt4lCp78LfuAYnGQxcTiftkjCzs1knMjKxPcudsIWUIN
3Jfj47P5kasQtzuwoXXEQsSCLu1QCOSraceitaFgG8WAhmK/uX8iNEQ3e0oS4VDRMaWf26merJPz
zC8Mcr9etNFd5TBdD6s3a2tFutZ2pMETOKn0YVyHzuOknbdxY3uZ3uWv8fRnwQjuvEwBNRd0zpA6
7u66QdOs1vYWmHAqVX9I2L9FCX3R08HN8CJI7LIY5iDlLBmH7CLz2opYBejvpa14DOZ/pCf9iMnT
+3/+9ouIHEiq8y9ItFX4SVZIvQMtdpCho8LcjYaosEFTu2VVlkryIEWek4MtVPGR0tUhnF3mBbwf
R4bXxRyw+x4Wb+oNk+sO826MwR9jiTEOQx5z3uLCVXRhtgOZC7BRiqIITthu85w1KrROq6sTLbgw
3YWbO4lw5XXs78F7109tw3Bh+SRR8SGM8QK1gJO76hISzLEwUU8NbhWDvLkCC20X0XGE+d8W38Cg
RHMIMF0KSyY9xLZnMOuqbZz0R0XSDUxVcbP4nYjBKcUOgL7yZylQUuFS1nB937PScNuPG9i+txrG
mknOhbguOEZGsIlIuWpQjNYlDLq+jPO4hLw1ZTgv4Sva2rmFi7uD7KZxq1HltnQ50JNZt+II+8LZ
WIWMQLk2v6iXKZwNMkzhxBlm4FhvnclPi452KRRGbss3ZQmM5xHvMtRu04IQSu5OKuYUEsn7I8ME
6kNHAhag3DMuQAC60z36O1CYgMOa20N/m7LDoIiH4T3YSQuv8hatqkPERAipXF7prmZCWLRnrKw4
X70+SQbymIK13auUc+rg1r5Ev4ihboDZzasj5TPdEdRXzz+WciNQnDQGB0YVVCOJjTKKk8v47mPz
iEChELqzWVZdVly2mId0W72j1lOgLbdasXvB7XF8CetCfOt4eIXYOH7S+aiHKjJKgt8UcudxOwC5
LuZaPtWPaRoIQbI3FmpsqT18JBHw+n9tnLL/c0AQh4SmFTZuudRjX/LUbp9EwPiLJTRythWitM/G
jkzUgKD2Gkj21fq/W+sr2q90KT/C+ZHBSXUzinoJXEe5GxcyvFwT3WyER1n7ZCiqbqZrNCXRM91q
4ABTWXJImG8ZuQKyA2hRRZA8UY/Y4w1s3v0HQOt3FFpohHAgMywGcCGxiCARjoj0h5homvTbjGE3
Y5jQExsIsvRK02jATX+V2EuQOk6MZ/p8XUvpYhajWi6kkFXTC3GujR66gx1KZEzqSsWvvfAQqbfO
CfsiKyuCDY7aimPMbjXZrwsE5qmdJ7DJmgxyVeeMRSryd7AhkvOvYj6lT2ASpeZAHuRpnorlV8H4
zn6x3quEsR69hZtXQ3/5WvkZEr8ihGBiSzY4B12MgBveHQDexTw8ncKDFNGlluWYMhf04SUfj3hf
OFjk4Ecj+XHcQFzeYVbtC1vNx2xJdH2/PvRjntqDKCgmmJcUpb7QCjBHjh0mxLlWKA3NjM+vw5e/
6k3pDAXE5UKzwqR27+tI/R5yDHiiEUfNNizQgsvScSVIsf8KX4ysZzeEVhRGNgXxnUD6iX3KBigK
UgjM0xkmgh7VIIOq3KKFbnO5OYyAnGQ/eE7f4b6UCf7dml6p9mPuXwUoTF71SIgn6kpoL1Tlzd3y
mxkBEz2eh9f8G/ejlPTxt2nPssMyCPO+sz+O+f992Gd0EnxDKMlvu3K0yqEpIZ3F/x96M15wU80m
DAKHoou30dPBWy6lW9W8xhJ9JZXfKomYleQnrxJ2CIKE2cplGi2ln6R8K49yVTdiW0AAumqPfL59
tm8+yiEyC7HFpyke+YzZ+mCTrDXVQdar2bKYX7fRwf4YHaU7gW9FvN8Nnhi0gCJrLp2Udbl2KanS
SMaCHo3/ODHS4fKrajdCXPhVujqfTmKwElcS/VPFFvA7+enYn03Y8Zr+I5Pd8G0q1m5D1SJLcF5C
DZ0FtFI+wxTVbdudB5q293foDDemB0/ks8EuN17vQkV6A8wIgC42xSOFiXWnzcP2LR8WQLTHTZXS
iV9GzHqFcFb9ZPmCHf/d+W2JyPrE23DQygsTCeGirtmCmvVMIy6RdjES5l+Bq4C9dgFNwDUuXqD0
NcXl665P4O322/qPFT0VzP6K4AvSgcROUwo2QVBWeLgfnD0uBT9Hbfi8h+zN5Mc9x/9hw47vvYQa
DFkbHSKetY69teCV9K0gus4PGhtPJpS3WaW+pGlofdSSDgfoh1Rk449nR6AATQ5UIz1S9BEac7w1
GY9fEGgUM6d0BR5O902EOXD433Q0f+5rj2mgBwZFHzgFaPglBPEbeqW3WKHIUcUpD0Wet2MWWbU8
2InzJe06ENsdbtYtNOUyPwHrZs3a87vPpck9SBgwhk8NUUOZbei7djX2filL8+8/umRxzM9rmHGF
E0H2StIlgzQ0nvUayfvfQYWnlbC0w5rLknB8CKwh1j4yoM7c4yMvVL25O/5CBfdPGAJH+661tTPu
YmZ7cXgIkZLHlgRn/4cy+qlMVJKtjdE9/WXuFROmG5ES30NTQFxntDTly9RY4GTOTTFslX9yYEOe
iJNSH/G0pyB4t/O9l7CXRAvU8zSSDXqOtFsw3GyD5CHHi6QTWodbaY+Y0lsrKwhB01HOCovK3bcH
kzprJ74AhCSwOTIyG9mFSiTucga/NAENy0U0vXBfjdtsE8katgRFRZ+65SY7tDMdHHGYqr0YrZEy
1AHxzAtHYyrMNvY/0h4EN8BSnwDFzaFA/y8PHPQayoOwshbtfX4gWx8hc39tlEG8BPnqv8/voCm3
TQIAZHyY8Z0b303wCf6jSf62YSX78Fp3ziDkZ2xx643guxu5UjTx7Cl8ZE80VMLY2/a/7BRHgeZ8
R7+9V+KsfZbcAo19UC1sJlIlBkiZ4c3aHRU9SNtoAfL54VYgpc3EHHhrbpEsBXmA76jHUTAtSh2h
/ut478VFieVoblTKvFxXw1fbP3URE6KwzNKFyoKWxDJHR5d+8uQ0ukZrEJMAtVdMVlSrdNaeDG5A
xWCChyt+WtqKAaAPKWBsJr9YYL0yv/grJ/oN0SxaJ/H2MEfkRdJ4QiZ3sF8m91UWig8NcvgymvLT
UkSfRHV3J8u1n8dXWbV4I34uq6trGYvOUwkdOl+ua2Apq9RTiohTANiv+STSF4CBb1LMyQUnivzN
fdU316A0EpIj0LhtLc36VDwbKwV57ud5ehpWP3D1xkJk0qOY2dQkrzS58Gcpt06d+u50b/Pg/5wY
Z/sfx9LINVkv8qBB4r/3c3Ou7Oo02OvWYSe/AV1llpfHtvjUh/1fGKcyCxoaKnn4SWt1yvX6PaXg
ptrkpFWFea7HVZjVQBNcPSBhhzsmwLuXYTxCFyEcFM2tje+XNfmpnJZu4PT/lQ3nUVngVNYgqfMs
qqc41n2gXaXZ6Wm0RpT+86XYdKgOqRRNr87QtDkRcQM59cdUidAK1NNojswolt/xpLhKi+FJP56b
uFL76JJZveFGOPnRKnO7w+4lQ0tjZwino1Wc28Mm8u8n0YU0WNjhYVlmAY4tEjxhZn3Bq3/dkmJa
Aj9SBnVL6wn2oCoEI0FUin6I9wVVYtFh4sX0Au31Ei6BcuRnpenA0tGtvNUS7bNR8c6u4Iekgo1N
0P9qhnXdwkPguzONc7YUSrflK5FzG1Dci2nxtH7UjcB82fXH/yLeFpgbDD7WKACfCfhsgAKpC6Ro
2eAxQ57KFdtFeCBFgnJ06lWMfu0RD7IEko7d4gxyWooJ3nw3c93SCOpcF4L2Y9zOhosvPI4t+8MN
EfcOAj5WOkRll+wZQH1bM5KO24gdH5SJErrSTH7pyU4up5RnABzxl7H45L0KuuR8nNqUbe3eYnI1
R1OsvjSqgBZ8kVE9mUdsNYiQSf349UMD6IJUwgwEsDx0b7DuI1MBoxPMnCUfM7IsYsa+5m3a/u9c
DbIb3gvpSOyYFrTqD5aJbLI2NFLubuRfrNoijv+vfMhGU2k9PRcCZbo1+Y8kfNquXBfl/S8qxYRS
/ucsipTxt4q2uZRMdgqnRK9jLp/uEQcLNoXtjIfOTnMVk2YOtal+XP/qUh/HZwdaIY1EqVGsLBDH
A7krZ080a6eG3cLCB7NRnGhLNN2QoPUv5s3kNlShxYo/9/1Fxyue678U9FKSMarQQa7r3LYgHiQc
IOuWhPzpkBp2aRox0RXL0YnwoJzEfbOZhyRHu/4W8C4oh4ikyBvH5uaMFCVpL6ZwBFQlG0Sj5puQ
5YWq4YVhHIocZOhG8lm8FiXBdiVlcwwBymnpfjdJgbV/U7BJR4bkE+vkaJ4IPjBLGBHzj6iNlP1o
V1MGrFpEvjBquh6BNz7Ceetx+Qp7kZKzvciPSN3p+u9/2moqf04MFhh+x8rGmAMvk5CiPTsTSPnb
+78m+mRWiWbFuD0VGEWXmkBCE6Oq3qN+MSTuPx4u2z+gKLLdC9c5WogGHSlRAYfCJ0ITXduPaKnX
/tRcKYEcqQFa2oKBfoLOfLcU+wc/lMIQQr17jbjH7mUPtWfbpjpPFxyDh5L8ebHFDj1PXQSp68QQ
0s1kdh0H/jD1neOgkK5z/qcMM0eUOd8zMVewc3Z2y9L0PGEXgtwrErpwp7TrnO/XQSMX1EeMbMGl
rj8ZslnodsRY0aB/NMJtP4KWpFqCw87o1Lnkn0VF7oURDwFLzbTnkc/IdYo58poxjE9rTDnO9mDd
dZyaQAETWDq/zN2DlQRs0M4jkp8q0uRkQCe3GEPFjEOsPfkucd7aeQvteF61t8XHl/h8+cKgqHUK
7cYK3iIm+xPzJQJHZeCL7dARoHQITYr/UerdNIafTIVLQAxNV0GM6Z/u2T3NJKYOUU654quqNHl2
C+negJgya+uoASagFz3Qc2iHneKBlIbNGn7i8rMu+GiYf0FYenga9FI9/IJMYBhTvLAglYRPvbbj
+wdl9enR8TlmO5lhMtJAZOyZY6z/BL2klP83ZI1yZ6HAP7eVDkO3NLF+A4GQMXb9GHi7tGe/E+qc
SanFTpcmXN6clQhfdckknDEa6I+dkVLmwnoCwSdHIqKzHe+PAVKv+nZVfEtT6mTte8Jo+qf0b6L5
M5506KeG3AUEweOwyYuNRBxlBW3ZRs//WLTnmnM7GWnvV9zNUXjr94IAHx1Q+BkI+ScK6whPWqy2
Kp7GEztguJfbHO0f8LJyoK3c0ZeSry28m2E6iBFitnZQz41k+SCMQfcatl2TH4XIzNX8eunzyZcF
PRSuS1D4ZQnqz6+MdoUyFKSg4azsuWfTglVOqu/MET6/TY+hebfikcjNBeI9IZBixW/2GTo6NHoX
3zsANvuVSfz8jDh1PsCvTG00wPPX0CSBdaCCnScie5kH4e/O01+F4MoDoq3v0afmKt+b0jCN4HVs
SKsXREx6+UFN9h0lOGs/92WtU8s+iEWAFtc/5+x0q95FR2X4M2qsrWZ40nZfvonW5FST3n9ljKY0
DHG7wnOITFnHaYvahPmm92teqTYOUBBzi3Ep8ZdPhGb/Cay+xOkGjiuEWzbC5HB6cs4PVNIqT2KF
ssiPRsVrc/vf36v/u0Iu5GjtCK91p0hIvCEg7hyq6hOgk83PAqhgKOQu4Bbb7TtbENOSVWiP9vwk
VQdrjoGj24O64VrAR1KK/owzVq2iHZUkYdC+yjYzgAHMMY5gYqpd/Impt9n48u9uRzdjps2ut0GR
A6rYQoHAuAoSC4rJ/euU4U/Seq/2aeLlsjJ8UaK/PxANMRwIRAPdab72ocAr/DQwAEVjaN28PpVq
ocAlQYt7yQpskhzLdmIYH1+/dl1IziQkucu2RVLCNNPyktidJmb/KVXvNEmK+j4XYmpSeIYAp4PI
qwNjXIiUwiIjgsMVqwVmBYN10w7N6bMN2y0jbQ1xYcBkKk9F4bmhfW+xxit9QCzNBKGSyEcp97zd
mWLlMxVYprxCA6/nHzHvxp2HNN+GM+ETE988aljmAAa5kVUUGBC1DvG0BZOJVSL7jqWZeeaMb4id
44aJcMiX1yPbGI0kKLLowqwJjiO52cFtpXd99W7XAObuSF9rrMajcZ6que+bkvXZ5dHgMVUhv4EP
AxYxuiH4FiNHIcLZAuefOTNyWvMpjZXo1Pio1C3s68nlmjG102hXhpXdpf8OcYihs5o5wHY/rpV7
jDDg/bmHqS1ofH8INBZHF0L7fDzvdIHc9qPlb2T5Gf+wJNCI7bRI1WnLlXfnOLB1EloGbrxZFRbP
cWd72UCMy5fepb/kMGkgwVcqFxp4/PlJRJEv5KUi4hffJp3eDrBvfYB0381wj3FXELdWPotN3E3N
7G5YBPueDua/xAXMhNLSQ2Y2bPJtUPH267/JDXx+P663sD5BAO2hdLNnq6QpZyzeb1Q+EuZ3jeI2
ZL7hmsUv6Yzk17JKVat8kkjLgdruRGo8PNZ6oFeL5kL6zZvuKdpP29qo2r2Z3QvJex9aiRsxrZdK
9deSHHnY1RIrZnJ2lG1zGyBFNJqFkNllt2sPh6vp8PfMhKOvdpTvvBnCGf6R1+3pew9gsEazrDyQ
NkmkR7KpYnTFD39gy9Cdu/8ySXsBDEJc9DMD7C4Gv62yMZ0ozDuwOuy/vhIZXU0r6qVuIDsSD1uF
WyyLzF8UrTvGC4zdT1k/zp9OjDxxyHRU3SZ4CDp+mES0WXdhCYzC6e3Sp2mtl/F/sTo5SEMZLaq1
E/uA9eNWhna6B6yk9GldJo3XoZqVVp+3Lgawy2Gc+MrPljeaSKMIDbBMy0U0Yax1tl6aAbOwC/cx
hti10cLoSS+XcjtoZOHARex/dJofLFMP/B/REcG5uwfeDfkCQsVG2F9TnPsKJI1F1sOjSX/Pjr2h
+uqBMdzqyK6QMmC71Emgnlx4eh7Y6aU7C5Q3llg+dXpRVuuUEavWpGmSnKWW7SKVPAYPGzDnBq2G
c4ndW8ETuYqGRDDBo6YuptYpjJYQypvXWqlbXsIRp7/PE5Rkbr36Rikzk9K6vlOpPW1izWhyxESF
5ltYglngciV8ZtlYWx5Z6T1ZVBOQCau7nMXRzU/uDNlGbuK9E853rEp1HvhL3UdYyVEtTpGV0H1t
LZFiGc2xux9bbY5ibpWuEkuwFaAL+u17oi3lg8q9gh/Ed8C1d2Q00CvrbMakRfjAoG023qiLmR4m
Yv+Sa6fMlR1ZG6gtNjhG1nkdOBwTRoYEOdKjSXH03VLKcLo8Su213iE70rLKu0hyCMtzEwC+7N3v
8qUH1ETpeb+3cE6HIPZNeUjMPKIQT+Tba870xIeW/Jt+pmy3Cn3/K7Wdj9Wl8zeKRojpP+Y6QMj4
eKBwqzkNm8s0F0DCsPiy959Zv3YcHyCCmhPVwez9TItm4bpsfrXoL7I1uxFLjsxHpIptU5EUBGWo
nuA31zLcJRFGNLm+HOOIrqILO4JZxMh6sUtCbMQSn207F9iWuS8b9ZvIpb0XVCIfIokQ9pLQNctf
rjo176Fna5DgP6auyKQ9qF/TIpFGAEHmWYt+FgVCde+80UP+To6kWmykBVcWxf5UW34pqMktqYH4
LUaFXRHuJHCPkkOl/bBVqf0JRpWGu6u6n7xxCPaHbTgmItaVAzutTm0jYmWkHsi6AgS3dvBzOyHn
7Jy3NjRwpzVoA83gM4NmQORki/WnDC89StdV+kfd/ESQzzUF7jvCv97qgE3K6VwwiM8+CJxmYy1X
uou19LwHf9WQG8srOhlJvANYI1t3VlzbtQXIkt3u6IFua+3Qv1AWuVpMZi5v/iQHlQcjLHGE4JDU
3q2cEZAqacJD+jZTi+T/0osD/Nc8dzcliytMXBkmWn+IQuVeWo61MKGY18H/V0EdFCPyf+kd3ugI
v+Ma/m2fHm3+/Pv8HNoG7K41v7X9/XuByENaVwOT/zcVDC+U5XU5d2bqM6+tGZX5s5w+ZE+Rr0a7
nfimUXHukrHtoSTbXRgbqZbj4Hx1MMVOPozu40cmWNapFKyUM5jnRsRzHBxQ19iyn2RGVVhE84Qn
rOy1Z3O84//tws9qlQGmDsoMm+dk/ZZiFHDsOb5UGqUX0u4ZO8J4JLSyp4+mSTT0rZ7hC0cnIjWr
gc2z1iYlrhwuEoABcEjnJK5RfC0SIiOwHNl7UUv8r8iqfLdnfEPPr1Ud/Vr4j9Q/l2b6YLFWffAL
VmmB8NEWn77MBe5uQSo1p2TTHq9qDwBNYx8uFfs83mHqTS8y/cWfqY3nfVkWoV1ZTNmo/Elwl7oS
aNLuO9e407AcnNMnn5hrcwEylmZMh6K9oa05rK6HYoeBqkajwhg4LqkbQYVwp+KT+zNRXCW57PYz
NgZ7Eia5bYDNf/CAKjcQhts6+ecCouMlILM6rcmQ0D89tIEFhCe+aSy8RWUwuVc5/j+FHEtNmVxo
eT/1U5SMR3XDAKxK7INX2hrIpR3nlx/pxlx9I965uv42iK/f8peCNq2KUJGVD2S/GQgL+zI7/DAI
1LObGi2qND+L7PBKktqmtCCY0REwOx7PReXdMAc9WC9j0wI2BGyiU75MjGGd7TrWofm+hU4S/KPG
wrcCfozL9cG3xWwmnP8HL6qckIAWPQT2c3fVS5HwjenCc3K3sva/sFSBdMWEDzAl4UMEurkTPWsK
Q3GoBaaH9lk7NGrHIf7jzd081klvfLDSxfA52fIkJSbX7Zp+MgINgH1oMlRl2n8g91sASCKEZUOa
1++aTQbizOn52ZwHgX+FkXCFZYwXWqUAApzOfBMlS/iTwdB6GF1Vxq301YWPcEcmKepPs6aQfmok
knd+OczyB3loydly+Kr9LPCAEUE8jYIk3GzXwJ95KBNrCOHwYVV1DeJFwHniwSoHnhw/LVEMlvB4
VuHvMxnQawtefkI/c7HahRt5IaxkWl7prrFfX1pbw0ogGWlgPoQ5rRwIVFZJ6mnddAC1phfUzV+d
KFmwzYL30eF2Eovh64rdL2zBQglPXODiAXCC9ePSb6sYSpV9oTM7AgIaN93lPEJntG1AU5Oq8XJR
tIKziU/VKPC+835P9ff5RHaBeCDwtHNNlF+xe71d0jMmKyAmoewOM1nLIq2QwNuuZwCMdeh8jVSw
5pJwn9+skbYw8XVfv0R+S9woGnnwMGUrdKb1wjKwCBA14z0XFv092R7JFp1sLj+wasTHZDD4yrs9
2MursHNR9TupjgoZ7kEv8j+yREOVYHk7dfG+Cu+Mr5XCGK4vTk2AAELyDUQb9l1IoDTBNNFAaRpy
wpvOVqFFc5cqmr/hegT2UWWW32ONLiHcmZbdjWNUB0YGFMl+Ainm3wAgy+bTqW9WWR8W6qeHHFu2
/GCyqV0pdaQ3mcXSeRCr6Wf2FMW02HsT7vv2d59jXTvbmKAsVHjttXizAn9E3gAA1ZrHbmbfon6Q
Pk1Wj/v6drR9KI1BwQKNS42MrzbzBN5/unbeHFT/A4zXyzJ03kD7DxbbLwvwfDLVtajVfh69iOhA
niGW/6iI7my521rg/QWKuGvEKi+TjEGpJn6NBogQL1BL02ldcNvq6Wq//m5h5nWWauYuwd2IgxYI
TCAX5Upi4tvdTO+RU+8nGv3pZNWqDA39NCJBTnwaxtUZA83SD3NcaZES63g/av0erpsPiyg+eVsM
pv7DNmB+moFhiR0EtRa22LCvxwYg7rto6S+0PD5yX14UZU0WX/amPRWTz90IL/Lqf3p0wgZhJKIE
xuwnvYwXQ8wGtRViiyKpqUE80KJcZWaZIEGghPOGfkMXQzb3xne3hb5cNDBXaPDJW7GN+pQgXVMl
LZJuJ0OiS3obmh3RWIOcjK2L2RQjwhik5PsJNvpRcXQ3S4FSpzO2q11UtAqpVlf7ozrrVkYRyWUs
c77iwBW1yHDlkXOXafch61x0aPfLnLy69k6VVqb4VsHa1MDjCTs5ZMqTlHjrCZnUVRlQd3BG1Uz1
+KX4Y20wlsYj2SrAT3Ldsy1+xf0+N2TTf21lbJuLlILf6rX/JmNMFb0O2btu3d/DroWxMB6ukKns
neacDKKWxu/xhWiTQi1ndOVDQmbEDKOQaOAEcRgjMH+I1qT/+O3KyENmJuBGbxKzPWitzFUqz2fY
KqZrSganCoACo4W0a2qzxQN3MvCHwELIUjP6sl2k++HUXJxFTKHABZAg4Fq0J9a9EMsJAd9nJ0FW
WSl7I1kb8m8kO3isZ7GfJ2L3HCVyF9aWxuLKqok7rfY3lvqSUKHUIlAwSHVUByMBY6aWpbKReODJ
ozCK4cMBrNXnBfNXqbTLkjmUBikSrkQqGwQ8E1S4Igr7cSP0vi7zGtsGl89P7uOU3MxHCej22hYO
5aYjN2ELXfk/seGtkYTuG5GB1mXkTYcfKv8sFloFNrKmgkfNcaaSwUHUFmM1vIKPx3wNq8tpnOZj
SH3CWuWKy+e/bGvgzf90HKxAlyIQYLL1qWshKZUuVcs/VIUwyNlfsqUslIQn5t3RSlrG1LggpE3v
fJoEJszmH+b6q7gqpFWzq+s3izZRoc3jDrrs3nn3SV/CYaIAYObSsjJr0EY991Pa4Vz1Yvafht7e
hvU6jPBIJE3ZimqJWva9INOZp7pTeqFVwfpWyyaLygDIsQZfkB7iSCZze4Tj9uN3hhQcOUSYA3sm
cLBe477A5trY268bFQkQwk9dyAvtAmOBD9dbJYckP8/c4hmf0Bs0j0Zjri1xtz5z43Ub+HFNFZOW
ddaAaOzOiZkTwwO64lNzUPTPbMoD59ukrD45D/ytsIyf7ylNBIRoVK0OItwELZYUn4twie7FJt9h
WheJIYerxr8YLIWIenaZeUlF+NHo4EmQcpdvvGjaUCg4XHdPd9sayukhwfFqMFoGvJ2Lagkowlwg
53sphycEwnrnKkrbnB6DXH5QA7bcBDL3I5tdwZv4I6t+ALRIaIKYe57Nk8tiZzxdk+MQZ9cUOjEf
Wt0yagSAGn6J2cgkldoN/uWgTBuDpfB8Zm4Pc75qrC2iv/JrJNlf9V4X6HAGfoysAOWuQ7lKglAg
XgV1VLmyWvAL+9D1/WDUijWKTquK6tjLi53HGowWOmBeTxGmd7zB//lCY41cKBTN8NBR8tf6ucPh
OqiIuZYFQdi4yqDGGU6eY28X5IifMF6oI1FKBMq1c0OlepZhP7nC3yWrbFD25ft3MO2eVl9BHCMX
hs2YUIkChqcrrJAo6kKj7b+fs1uMO8ctXN4ClxYDWvacRPjmk55mKhAt0GnhOofL0c6LG6EecTNV
6++jsv3y0pQYw/Gj/g5gqUL1QPkSPiTCUJpI3vGpR7AKpIVakHzu3/COwlVKxjzN7ifIeaMbl0zd
eD5TAxlWE3e0sKOvgqdoQ9ECdVQ8GqGfPFhhPU3dAdmoyA4BhtSYIco8+FfRPGIHzw5eNZkdAMPd
2a3cz3IcpJCfYVAXY5bf30j8YLkxbnYzN88WS81d6VT0vJqG+BrPr9LgNVgX0o9Os093CCXQp9DS
XuTuCn/7xkc+PHLIcm1nxlASTWxMwoaQF0Fe6jDXiIfOiv5BZPqMzNM6+/KTruvNAcHnlHONfaaC
dUHEksUm0iu8XmTrOvZ4m4y9wRvHRLNqOV3/PsJmfTXPnklq0c3RW5vuwd9uhwR4/Ysc9h2xQK4p
b8g938F2WpcV5EnBTA7TBiYeTkfCRPcW2ZBmq4wTP3tqSKKoiQlJv3otqCbNhwaR/fq6uROFiAJ5
HuBB4DtAEFrYL+WscIJdeBO6GUAkG3GlxePuJJlcre0AOo3ex9vQu5gKZoURiC/mnwKVUQcVvd4F
8VWoIdg6OCgmDT1Zcb4nAgAMNayoR1BXYC1FgJOwxBjVVv/4rieFGIuxIHeIv7nNPPtzR3JYGLqR
hxnqRsf+8nqbb350Ph/EHoQGPZPQ/4+xL61yUut6LE7cTJdMQ7oUQUNWbg+YTP3dGpaTkatQhCEK
cxfm+z9lgFnodyvpzw/aVoQTBTnc7mAE8D7u+EF9b0b3RBRUt+/OwDHMl4QKM21X2u9AHv5+sU5m
ysi5eWBR/pmJ1Ss1pUyrmgqQnNqXR2LVk1hel5POtwfIMn2DPkzJ3kO65kpiMc2UMqtZJXw3/yYB
g8UMngvOfuk5juAwaJA+vg++QHWlwGSzJBKZCrxCBLuNgIedDpodrhZ3j5ndyNf8yPe0AP6HA9RH
Ql/rGceQl8HVvzcpuVScHMX3Jd2lOs3+HWgvXVoDlJewqXZsmSMEYwQ8xQpovG9I/kjHvX3D3MDE
2ZeXO9S1xvXQNDS4fOmswMJHJ8j358tz20NTDA8SM3UwffuWYugy8ZxxIXnlhx8h+gODlzPqAjCb
iYlEDxRc5qoB1paEvEDn2DhbJ8KYfM6qeTpPoTrodTAzgkFXJeKqF0QY1m6A2DzsXRT6S/N1rFtZ
mxobvG2Gxpb/YuuCi9ORTYNDjrJwjPODtgplxvlqP69w0IW6LqdW2FCo/Jb9iEFRl7xeahWH0N5G
y5O7Y0AvVMSUOjWWr/ICZzulT4UuFZIImlPk87Fv7lUYZoHIm1LLh/91MDxjW99jDnW/T8HsoEii
2i/pRGYh8oVvY8m29VR6UimA+GqoHqC4AmB7TSeumqWuS3NNzwHb5ojR+92QcfdV+7cL3Sr7Uy1R
aMP4ybAA+yBz8Vx3sGZnsoYfr/u3Os0sEnQI2uVuuPwtPsZoRYPk17JjQqymoa9jYSlFMMmpE/dw
NFfJEzCXrTQ/dxbYJpy7Q4ldzRyPjHxJwNbyTQnJNlMQadI+OiS04e2zjJQQjakBf8i0oi70su8F
J/PRVvMUO0SW4t6CyCteoKUNsB4o8KTtLCICJaggm/8NGwVa/FmcKh7Ci5kxwU4ahzKL78aANbwl
WL5Ve3dquYlMPnSMUIhbWpCICD6errYcQlGbA0fRIyF4cYSFzkqCdLRhtlpsWpfAwiemkaacMtaI
0tfIu4r1eBzkAGQQn7J8w0zkvg1sSYnPI8ioSS0wyLM9nrDYTlIOgMvtjCqrE4G6GGT7s4+Z7FK2
mzocHKJpWT/ecmQcTvJyB758+AuCSy/NRFQ7N+zUlwOaRKmMri+ddn2wBFTUhR30KP6uzKQeGhrB
a7AxLo+1IrEG7SqHdUdM5K55VW7MSehzXZjuA0man+B0YCZTWGJXAXDYzkU3+dK/v2Qzi12eeYLc
Jmvx62YPonMV/Tp9iTq3SO3Fh0N7rXJ0n/Fn7i8bJRo05gU2RY0NE2uPWbks74HKiYKELtiDItTN
+WWtm+YWILMDmdZUC8AIJ2ZmUqvBqfKkpY9woHDKh9/AFS8/XVJ+nwxBg7vPGb2g6Awet9dSzKGw
K52rFD4T7mz4C6NYvKWWhfu4UUcvCz9ZtgLQKFZJ8ijIFJPCCDc0xoTW/XDA11JmF0zJeZW+C/i0
5CxxQRb/PkPk6qzpbcoDDXZLdeF6vFdKhOSOFLliRqTTDFO9a0+Xr5gN+LRff8WExPBJIAYjBy4o
CYert4oIOqIj4rfceCrH4X8EHs1gLNQEENa4aM2xPx2/LOvfxIx2PFUVe9J817f23m1ALZTO/8kv
QQdu7zYmCEoPYXlKEuYdUdfzAtRDhaIWoj6fk78CnCi2u+iCWP+fr1fJ1GAcBoesIc74aPh+5tlS
naKP9WUgsmrnhcZVKn3Us7uSl6rUcp8x4+jrBUmR5YdVB6l5BAUgAtxJwVRvBKVs6CzUuQcHSYKr
yYQgt/pA6Czt9e4BWSjHO8XWJY116MPhW8mtIe+APBjl0OXB1wm/KgFsVt1GeHHhwXS0v8Q7tQid
jK4aPsIebwY7fOSDeuwWUk8WZ6hALmurWiolxwLgfU7b9DU9lLKqpe067w1ZpMzQdy4eSqvrZyr6
ooLbcUBjWqkpw2fINBubv/SXpM36UwC0z4u7T5S+qiWyC1PyUTyKDyuVXKZ9P5QgN6mKu/TmErGr
oUpyAZRKsrI2+G8weCS7KJrBV3WWdvMzUZpfzP03JPomJdac0yuge/AdnL1z5zK2/VIIbX3qShzl
HQ1EM6sqN614Cfi0PF7SmanDy4HMw3DmypkC4Lo/jRbIpwW6hy52lQQHwFKSOEQaQ6fTCgq4iTpM
6gJm7h325DItvz1+OeLxwIGCxN89BLSngtZDIcv68M9WdNxUart9uKOb0xgfOdbWHm1tUFvjn9/s
lRP3O0QMsBxkM56OcEy9+GzrTh6SpMoUY2hMy2T+b6gnRIT/7HDfkWOqc8RjcFJ4diCHeohmYuCi
Ec9tWmcm+13fiAi52oXsds91pRjl6EZ2ApaJeePvghM+IN/U70KNbxEvEk14TXFj4bIvprJEUM2B
Ky+KPMGHo/Q6k5rtYxmo9isoF5R7um2Jn7nSnRlBufDG+p/Rr3FQ6F81oDzmlMb+o8VJ7UKOTyOL
1jtXtvJqOSAEyL1N6TPiGyy+B4NTpD/xOobb/QQK/11wInSaOYZ2I88KGTMinvIxTYufiFQV5utF
A4i1Y1vHbk2yU8TXsKmMMXe2P7Ow/OmdWKNvjfqzDBG6mRJ1pFASa0N1xfvYh6k1TeVu0XIuxbbK
1eaSxyv4OtMnyT5slGihUQgoP8auKNk/+L0X5Y1CEp41KVpsOKVdwUuMue36qU21gHtH76OzLIaK
44BbO8d2Zd3PSXsoQ9qo1IcUtKPqb22TVQV/gVE8/0qviJCPisUAbVBVdYRIm2YXsrGRP4evolfC
zEoWTadcscyFkr8grBvEYy7TI13Vc6kAf+pROws6wv/cNicMnwogFfbPmR3aEfAXz7vrwRYv/gOr
UC1ILHcVIQqrp1FRFz/8vEV+V6v6R8UAKe51+51Yrw4HBP1ru0qRx+Y7JAT4O7/chS8AQ0qO+Pym
1VWsj0jHBYJbX1Di2WEqbXD9HaYteOgwaQmED2LkvswcZffV6Xv7Ou9UXjXlmQqelnksYDlSdMo+
m0wkBMJ734VIbcZunL7btZ9nt2xmf55OBfeX6WiX1vikq+QQXQyLuTbZC1E79x1Ng4GaSs1z/198
zCAYrJaVt6+/JflzUwDshGsAf+K0HHrlAyZopzOfofCuERW8ASc35NGXgWK7HRvqbdRW8shitaTc
titPX0OXNtmTHkOtWCnRSu1Xlt+a0giBW+MwklBijU9uguIW559XL5lAJ8wqG4jwQJzmw7cjFaly
Ug2hxbuG9k9BZbgbD2sErFyNl+uSTrlLK/NjkBrgcre5PXG+YvRmxqvOV5/5DNrHPrO3t+Vb4paB
VtWcL5Jc7xwhyhMdpG8YTFcLTSzp3k0C8lVDxg/79RV9nkURFPI+5DPjqsC511JRhSuX/Aq3SWPn
98j2bIQ4ZKR2sPGWO0DrKECtEYdLAmeDqiMIj/q7OBtR6nkjv3vE18uip4VxykZhG3uv+KT/p8Lz
k3sXYfmx7Hj0LM9C2r+/7um74Nl6NrStTodbRomJyvLw9Dkmi92MKGqSB2+I05C/YKzUwJVnJ1yb
73YmK81am6YhIahB7NQlZkjPoBZKoSwmmMdgxc3QhPnoMsJawlPX/no/eLnHrZ4P/+JNbMq9ZxYt
M+9leS7AA0/4m5uKM+cos7VcTrR5Kd7fTrQxoM5UJbtB98mbj56E3032J/FdLCcBFfe96Mz9JWD8
YY9YziUoPUm8x6oTIzBgfRf1fx8H4qPIoFFcQJ3rbkip3vHgl0PPWBZYK32vm9KQrmU1iNwOJgBf
H0JqkaibZw8BPbT1N1vlDspTkPoXyKFQktYrEbhhKZJq8QLDeyUjUl1zSGnWU0MsWpFqyhnp2hRB
+jQhHTDljF9+J4OzR6BZVuJMn2OCYP8CMT27CnAljsrY0hWo+2maKLmsafuTxnX9TAmda/2tNLGY
pVMyuWBH5mGI0l6DTU8UuvrUHt9u0OnY28009fZXobkw8nA7ZPyHIJ+PzPTuXeMarC8x7E3zfd4e
y8TlHRNLfRye4PfNMomkv7UVmUMVHQJ6xMeugaWrtUVhYCaA/fIIqCr67F/rK8cYRQoKyF8HvWDl
00JMhuTqZg/OQzXOna3e826Ir+QJqu9phE0d+9QJVDh1AUGesJb85IB6v429Oh/RCNZ63sxFhHes
LKEfsKyjMyen2iBgYwJq9sFL5SgDu8MBjVWCDmSMziuwMXb+e/qTpXLkRT0n7/X1e2k37JsEiwCM
WRheYEA9Hu7j5IXoTiVCNL0MgfYHWGk8ZbnKuKjFkjBPzJtaFjc8tdGqWUBMiRIBoXTUGTbewex4
LAkVlvXO+RT1FyUzfcXUshL/GOOyP+wL9gSocxd24cE/p6OMofpPmwXNxhRe2EUx8HaT4b+Cw/5u
QX3Q+UM0YDjy720vrIDhNzy1+EX0hmnNjFdQMw5zREWTa48lWenh9Bcqz00xFOWBtvtVGTCJkmlT
5F7j6B6q/7dxL8sjrrLaeVYuF1RAPWjZ3H2XV35OBuimpKYoCGayVifksHxEPNP/Rx39a2Ut+7Mo
fNg3Lf+jBJbQAyLIWdJ3ZPbMRst4cw6iPk7Y5yr76aMqojWDC5uTv4M8m5LeGT26nUpDQWZ2X3PH
fxbQqNcwreQ+cy45zsfqDuVh8acPvtnh9TRT2Q245O5DOU8wVlZw9AYdFQIPHYd1tIvgPVQ10GPq
+nt+e+ZpX0LqfsRII6wTUevmdBT7/zIrsyMUj4JmpMG9SGcow4tkBZ+vUu06fJ8Q6j93r0d30jAZ
1Zv/ot9/Am8fGypsLXLG/+XVU/jGz7xbJQxAHpuO+AnbmpdQDOBQ7bLjWj8e7VMTwwsaqSp3hrmr
twBOuP3j9Pq1qJJ+9zAKnujGnleZ1BfcgUJu6yjG/1xWe+20+1uF/nHB3soKQJL+o1zbamSmxrs3
HKh7t/vjm81zE6od+DZlVJpad052Q0gCaVktulDSlj58dA3grV+ad0t3zcgvlzH1DWFd+Jp/i99l
YJQfQYQKw0gO6/8A4T/eRmE2yxywq6reFya6nzLLpGTmcQXqyQbmErGb1ZAajRdgMU8XL9onXCkL
jrLEFDblCNh0yAVIeb3odr5pRTInpMNIVGnkzIECgsc1bpEUEcQgYHvmgLIYJoNUhVZaNOa9YvTG
ZW6xu+FatTgDSLP05zkFYZKh5+QhluA3bKfVhM0stb+WhKoGtTYQoVqSpJeVVxof6qAHdO9Qg4K7
E3rN9SxjdGpoqO5bvTZ7sxc88oMlEUXxLCaM8A4yOORdwYUSiquUMq0hg2nn62YFV4HnfhhobvWQ
+M6Ly6lYWSLb1QrjZZXUQDtkjkhidO72kJTL6nU9QjUJDaUGJhI0CYjW/1lG1TXmPiQIYjTLv+kv
UX+NMzOdZBS4iEZkwI61iOlHp3ia3LCRONpxqsDB2iMUukzPSwm2/6YX8/tg1ugfTZQlFsS8K6yR
V5ugKLt6aBNWWWBejlNL6OUXtcZdhj//cNas/XpjaIHR0ufSb/lGg40cs3uF2Su2rlVsf4o3JSRY
Kb0RwfB7T61gECiUwCTMnxSmrE3cURnJjFLQbTM5W44QeUO5BuPe+PHId/TM5kP49O8Yk9KJ8mei
J7P19C3YfBa95txsd++huqUAg/X0H2cM6GfJ5fcGdLbjoIBvpkM2zmXO9/EmnRZRHfvT3T2UlrSF
a5Tw0GJEMb27EwHLuggvNfUO87H0sck5xnAqi6gLMwFvJuzr1gD2T70FYypTemc9kmidqMKZUgdI
RQ920e3ktzLgRsMbcsgCf0KEl1k09LzPXPoev1pHrGLwjzFuRwaZhksqiuKOxcuq0/0gEuyND+dh
+UHxHmhIVmxiiOPn1rNK33EjFaSBs4+OXH6tIe++U/GpeaPatXPM1SUC7+um3SMQS2LbnOLGwpOq
+UInIqjjt6ZhumDamvkLItsAkm6XVxaeIMN1J8UzPVNsTfQ3x2ykObLX2q0rvs0xYhxjuENo6Kwa
74im0tTVvwd7Q5s3vUFzx3DCQSMDRl4AG0GRvR+Dr5GmbqA0IKne1j6+dwtfdAi4KdINMBGnmaYP
4xY2R3DGpUhGbnbVidLg7TErfgdh0srrqiQDqL18+9pw7mSLaUEv8kNjb4iuN0mP21/slx/JZmq8
rFSGmY/zRApy5gVfpAhhCSIwn1UmWO6vomZiOyijFcjuriTh6lXYqelQSndIwQri6ZujkAh6nyOV
IpK87ydzI2zmLok2JnH+bJatJb4l6GR9HZ0D0r/EpLGAa/m3wNdwfrszsssuVhHzgRcVkP+FOHGF
s9fRlmfvl1jWwPOqHalBjyphwR9Q40yRM6Z1K1M8P/D6pZKgAH4cSpX2MSh4nDCj1kn9LK34CNTZ
vQIMjqS7ASFgEWQXdti1ypxdL8IfCf8aXHzUzWNfEayHdpvJGm+8HqH5kv0scOg3rmPRnKrH95Os
0gs9vbDY+45CjnEMuKwxlIY8qk7hWruiBcP7KF0Pj6nhvSbN4EVwM+T84GCqAg+tRBB4ebNhwMwu
z//DkB/a8ecpQzwxG6QRF65Ur7XNK9JFKT4//IYgHCxRh770QbUrTFxFdyCdpLSZHMbs0tyxUda4
Ce208ySi3j/q1BOVx/efci/QNZoifS/oundK7Dr/yC28/4I6/wtiVbfoEtrPQkUE5HzBSq6MaBJl
QHBhtTVccjBc1WH+yoQjHmTTG2uMGJM3gGcz9OvhHWvv4BfZVFg6mTDsPUW4vieOMMfJOI1/cX88
3iceZ5S5O4m4imo51XEXoYPfEeXPnIb9uSPVji1kubLG/YK8pRY2qMRpg14aK3FLjZgK44QyeEjG
0YvvFE2KhjtpjXk/msaMnqtwnNsXcwF27HGHta+UuhUZM0617OABaw5perGPVEsp6gemk8QOnlLh
gp8zMwBF9yduo4cM0+vHfsHgQwDq/9hVln/IKna/H9YbHuTEJadIAfQSJQdjqkSwNRuCooaBUzrs
/v1bPZphMwYEtZ/JxJqc10JefuEiVhmfv7qRIe5Jkrcc0h3hYb/w3JMNZj8+OjniNQbnFti3bABa
gVA+R1GZgubiCXfti1PNIIb9AlZa0ppPlFZZQY5vlsAFeqZFEIpZO0Xasud+snI8Yg+DuxdFxveI
GrSa9gQ+nFVG+1Zkgr5jVSGfM3jps9FCN5i6TQ9yO4mTED5doqep3nK3Ec94bZslL7EKjU0y+Sr/
dfxjdRkhxF7NqOU9su5NhH1vJiw7zYRqJnNkA7uJQta2lx0qlT0EJFZJuB16l1f71pMFXNJV/rNK
hMr+w+UNsRhqwqOpIkk6GAbpCFGkgroe8E4iqkr3pWceHi9gp8TgAYlu6ccxpmsLxBVDAvjVTspJ
WlOVAYRweGrdNA8rqGFIBKGS41B06FA+DtldkmlwP4obpus1WcVriz812DwhAZDSY1Tl6BGgidyj
HtqRIG3sVwz8XVqLKTKAgCARpqOKtj9iElRsC2zKU6KXBuY4rTulkrU5Y6r5B2xwwrPkNaXPfzk3
JFtee9mVD+suxq+rfjPUqyfrrTRAHqYZQYxbnlrkezNYlnkbSKRKmn3TZZfh7ZP0k/A2DAo+IVLX
t+jl1ADWxecDa4oYgK+AiNRpk0elyIa5tEB/cAgTcwouytvAnfTiZsntikWHG2H1Zr0HMI73Q3zt
2qWROgfGV1S+fvif0CrtvBCpGthhNoL0OvMk/YajydkY19MRWP6NtWR5t7NsDaea+F9PSoQT88jI
jrYpcz1ZsTR5TiroZ0C+2jl/40WoNwwQIgtN9Gy4AHj8vWhDR5/tIm4y5MkObZyqgKQiVadqazS9
jpjhVVb+bQQtNjO/Iflx2jekD7jkAHlu2Sv95/YIXap+1K0IZORKdZmsHKlcxwt5PQPJkwo0WNuH
cigRttgo7Yx2+KLugp0NK9DtXuAZiFQcaj2HkNiXGQ5XuOID6Ea+gDVoAm2jNoTip1WlkcEMuI7y
c+tsynoXuM99Aazaiz2/JFZ4ueXXpLPDfCcjv5eDuR9+yL20unAp/FFIwuOtvObMNqbE2SUoF+Qo
B4xa79J7cMJaQAhJFmUz4t+meah4YykYyI4z8rdUgp9AMGgg6jBe9dUJZG36tb5DqTrjask/aYD5
f2f7Z0oNUC9thzzhoANSuooiX/3GRn3b3k5wuv9VKZ+X4xH3r5wbOHbC7dzFojncRISHC2bgwjER
gNzvv2mWybcLuXMOZHWgK07CSO/BZNX0nuAcO2vBNrtd7FFC4173zs33INYYvmIpx8u+Zo0jAk8X
r/SVldRnGgLiFgCZJFOOyaLCn2JQa2GymrIgIbsGD9pmfg+0BEVHK2WO7puepvStqL4zCkE4KDz/
UP+AUA3eQ0nAtavVOq484xkk0aPbs/IQXIzko/2hS/RXXgUaCDErAV8RndlUb90t5q1nrsEggaJm
gbFhPC+hWpe6MQF4LFe1Es3UjEZhhUgJtRrAJ2INq/i1X6WG8XFORK6YtQrjn+T4bS18L5kbcWfh
iH/ZMNGYGG+ZB9SYYvQNVCXj3WDYM+3Qm9/K0Nqap1my6L0lIqcO0G2v3B89hjO+lj2594zaDPyn
fqeZ6LLbJR04QrsqgbQC+GZyp4eXy1oNWSBX+4lCiEO4mlcQ2Fj4QhZhwa7jXj05tP6XT89hJDqp
TApeY3gLv+3bIg/b8rFJj6hxxwb4tZC1JDj5sbSmq3OpxKNVxA1FPwa1TcXvXrshwf2DdyDln426
xTyFJeTrvB83v9Vtws2EWhPhsm8vy6NApbFpZeUeZgH6js4ipqj2MDv26Na2yDxt0QClP1xECwcE
t9Xe+534z4IlOLG0iXYIdRZMW/5/L5xV2jTmdmX6Ceaw9+5LTKjc0TzeAaeN5spwdk1IRkc+NTQW
WXNwuwgUAM53ucQiZSzzZ/vXzverBje+ia4ugCNUAyzKmQNCYLahWRngshaDEDgNi934O8cedKbn
6UT9/DHIWegEDdZ/S1M5OGyu4nxscOYNYR+i+d0FuuAlEaM++f5EIY58VD+zuTYDXrI1WmznWTJE
0pVsSHiOYEBOgGpbMq8z/63B7FTRVynry8UJcrzxtDNYCKTs/Zh6PPo1V+kTDJUquf2ZEcaX/Ri7
a6GeKBInVkClavmJiyJ3nsmQF2OX6giW1ps0YdQLKXxDy/yfzpHeCr5MK+vaYqMyJ+5maVoAkceT
jVliwu238aYJQMH1QmB+TfMZ2HaF9OXgSMNDKO6PjQbS/9u0iOzPBJU2Va0rAbHDjBZahZEqJCOI
q+7UqX/gUq92SquY1KsXRYWX0fLOOOZdGpKO3uvNX1WS6om2KgApu+IzBt65xvYShi4TVLcC6Gcs
7ys3+R3aNtnjJacFW0pANAI3u47hYoDcGCjtAe2bOv0IwNZMZQvHRgzDMMIa4CNxjHgKZP1ZX5XZ
Xhd7H/wmf+UvNF/eKU8ERi5wZ7Ti1uYOppHzu8wBT5rqofQr+f549GahbUFFFcZELe/XGKJf48Ep
B4LvTN8wbZ5Z5j1z/MNSXnANDJGraIxT3/kCj/TtK5t4LW0Ky2h6+SfhhY836K4z6SkvycYGWyuT
i3+FJISbzmcqn8skLaWfrk8sMjDBv6iV2wFN2Q85MgwSQnEZzxnexmA30OBYLknwzNDY9+2qo8Z6
mJilF2nr2GYtdAA9YW68JEJOF0HGYgNOkqbHjtpm46qubh/6rWPlhaPWenVKxrAK+jTdnPP2JVZR
yOdB7W7IQF//zndnpeNHBNViaFpS2Ca71doJvkkf/T0u8SAuz8XO1FImsfnZWe1KXhBCstp8jlOZ
Yy0Ss82gJ7quvuwcFX723SXqW98/VtbYpXig5wEe99Izf/HokOo3IXDMbwQZjQNB3RJfIApiwUFu
eepNw6ei7dzx8T4TkFirCTWfxyxEtFlAphjBkQNG1se0Sq7nex6hPv81r2GL03gGC/mm8BaISdZm
oLQg1NrsA/hV2No8t/gK6rOaUXCv8Edg3mLGtI6nWHksgjSKUTlmR6KCUdAGQEHOK3jHgq6R76Lu
Sw17mNBMrvHAiAEMZ13onmknYthkpU6toP+BsB3lSFzo7HAOSRrQznantqD/XPxLf9v/F2/He6At
ZZfzXu2AnYAg1WTSonVFrDJP+k74V4YwowS/grrrsyN5cVg6rhibRdZ1hlDn4RaOxP4+mKLjYfkW
I5gRJdzkQWyw039eYZvS0/QjIgV9XwEoOeolEjjI2tvceHn3GPh6nZ7eZsI4JmKDPDhzzhzWgg48
d9VkH/xiDxAfVH+G9UbMdEjB58E7/8phO3etzVUIjKIGbRobVZd5KxQLQ5qIRNVrO2rRkN0GpeSo
ASEGE8SonNck1Coac7fGNL0DOj0EZb513B0IQSGLgT2eV9/8PrEjA8UFVR/mlzuMS592Kup7yq+W
xKFnbBkgWCTg+gwJZgMq2UjwLz43aqpi2+bQ9mnZPjdrW6Ut/NbpMo17uMXL+Ya8MFuTUBF2rPYY
ThHE9Cgb8MEJXHBEeGjC3srrxTolzakcRgKpdy7ytgBj1NpovQHQoAi32GH0zGa89wK80KzLbAQQ
W7DYuDH0HK1eXMbYSr/TrfBgofqPYY+OLUJk4nJNckswx/KzJLjxAoZD8Z7r1D/LtXr3WZHN8Ffv
fcDanZzfzEvdg75l84N81BD7nKcua5yJECdX6dsOdmHuMLG1dJL7Ls/6pTbhYiZbkbeOISsaMmJI
fW+2kQyLl9E6Yesy1Mwg4p5MVK0GQIjyndqFzUS29I+bNIiLQVy6jf7e4N0FAkAzdonfcPowdb7L
pi/UFSNakhFcRwAhmFKAmDgN+sgkJHCW3Yiq2XwoSVLroekHYfx9vj1D4kkeXfTUErdVODWNZw0Q
Wk0v/8iTVQcoXRTjA5Ub6lhbCYN7UgPAjNGElkenq6udOzz89Wshj5g3FxAF0yT9sEW78orX7D4D
9RxLS9iyLCc+Vl4zNxjfUEkwzdhJxmnq1WaU/O1tohNfbK+6W8DlGBQAK7lKW/pT+c8xyfpUu1B2
QW00NqKVcO8h2dQoW0jLb5nmAJ9azYxy37KRENPierCeHnaNdkodLsqxaU1ZQroXbiUQSdi1XKZE
u/dIWIAGLfJlBhDKw7YYDzaEvCCC4ENFrQ/aYJv78YOn1xmFOcQjxkw+e03v/WUixpNPFVByK+G8
+W48EaSFkRK0YqOHNONw/BFEVVzmolxa96xTOEkKtlGNeWnJ0wg2Y5xy+rvG1I0ryc85ZDNf/MaY
yumwu40b9/DDeAH/Py27f9VK8c4bSDtiC6m7mk/UE/dAvMs7WDCp0iRdnkvQ8/iXjJu8XOtArIWC
5+w4bLhACzKYeZEegiSmpnRCoL1BweP/ABqSQnUxIpRqVGoFhp5ZVM5yU9kdDZbqXfPkvzIDj46F
bqU0JEg/TSadewxmlgV0xuYdEXJ9gbeVL2/AP80VUbDUoVROrEQEms+peas3h5BpFO8ivTmQ+5qX
x2LcUEzICQHOMkF8joPja7BJgwd2hi2t1Yb4hJzL4wDVNP32R1y8Xl4rc2KU0G6G2I+zgUtR6K6c
J0GL8mJSb5fcbtSdtUbaCKq9VHywVt4KT8XXCXszdTiYM4+8PZNxWeEwrWPP3SWMQhD0WlEf9Ykw
VAGnYZirvebw1CvSdNYtIE10axUE2EAJz8+YjUVr3FJfRLP73mwfBPQ4xFzTr3ArAWVYk0nftH13
oYMqEkvHIENGYa9swsXzjvp13Utofc8AlrO7A3xWW0ebuaFIDTMRrXD3bMLMGRQxH9ME7p7e8raB
j/3Wue0V1kwtnd03pWpZxjK18dKO+/Z6SKEU8pu3Qh91eGiNW7oXgilb0w8eelPrtuoGF1t13smv
aivSTOeaHkH8NVGMQmIN0AJaLblz42E/uhDFe+vUx/UNWc05IWZf60m2JucDh2dammqcbXn2l2yv
CswWUg440ncL30l/phj4Cn3YbfcsIrfY0TYNpvYJznkdtA0yDNjkQnsZWzPweph2DruklCOZev0F
bew0JZNyaY755iMJootgV0ws/LXgrU5yr/LBXcl1ObAeTn2P0DCDF6Qf7E3XF2o/OY7khLXukbLc
ASh6T5Eys3lwgwYmR14BCSysTObF5YEdHZbrdF8Vu5XAEonHoYPytxkW25CmN9GLGckb3KcKAhGU
igBg+PaHDsLbVbKE4JO4pPZDKWt20ti2xFNhCiyh8bV1XN8dKX01aRPstuuvD5alMOgabtuVfT2/
Y9tDQWFt38xzrNAq5RxToTnSe3RpCdvRzbRK1F7rGp8DJuSuLu3TzA7h+i82Ta+u96/chvENoror
Y/yb90qhTTE2/A0wz2wnP075/ciDst9zVXaDCGORTC3AboLlYfjQxyHKGyhvzBVmeI5Z7ZrKv2A0
f8fPnkM4qj+BOpUUy0GInf97/UwWbu0yGHng5CvuHGaV+p+XDeZ5cHy4Zdq+2XOireFfuBVDQpZN
MDa2ljN9ifTyGPFHQRmF7NzV51SBeQ5Erm2G7LCFk70LS1R4UwhlHWux0MuipdjbuOHk3zQxug2X
v+dOEqEOjTXzZoeUdBFbxA3xKdrgfa0MqTH1qjTl8J24g2cLbGvUNOdbR8k6QDSo7jX6WU68STm3
j4H+zGLNErNV87zW2fNkPZDGZzKE4dqPPL3Fv80+x3O4M6I1bHW97senANK0X72NlDm/2n84eoUl
0+W/MceMl4H7EX7pwTEp2zNvMIKb0FCnnLKC5fm91zW/DSSEne2+HCiFEZisoBl8kHN4Qy7dghck
r2nVBQTpl8l3JMqEqXMox4I8D2bZ/usjqXuSb/cruv+qAhVdSJv5fqpJpBe9bQaBwGcpAq2IUjJS
44t9iE4Hr8b5pdxD25UEuOcxqsZy6jNmSNB7MbtcyRkefRVshwxPt2NZtFxeG+GccoUOjbBqUxKO
Dzme7ejU65l3v8DKNijqijutPr+qxJRcI5NpuVOhULq6p8al+FE1GX1WhkU2OKyLr7vWxOyjO6kA
FQsVmX2dm03LifaiZDsUT1X032AmPak/Q7qOf8tC+T9wCNDWuJRfawjllCduBN7Yl7pd1oiwC48h
bG6fKpgx62fOulf3ZDQjKYnp8A7l44+t60D4PLyv87RqsgC0oYGHf+Vqk/LIoahU58mG6CMeAmg0
fdIQ7EYWxWNFu5dZC0TeSBCrK0n27UYZUUgCmEICQWCadXi7RopL5R1Yah8CkU9JdG2vNgrDfpAL
vrmEgZNoflSwWgyy7PPXtxPX1WFQcpxHNTtRZy7paD2F8TXLJQfuaDchp0ThySo6WiXktVqS7ADu
OUItqlw8q6P6/yqkOum4PJHd5Fg/9/1zjwAbfMbRvfVVGh4bW17U7yOGXyx+Lq8vV1IiBrzPf1VB
PwaMKygbD4SDibcE5kg3nlLppDG2AmqF91f20a2ZLvOh1+SVdB1/Q4IFcj9EhqlcdyShRa5IXNMI
6GlSK+3KPzaR3Qqk/fYtV13UDQw7LDNH8krbB8cuiZTKaOJw4AIXpQaIli0yqod5IMWltC3UexK6
AYMyGlQoed8wQK4U6Dbxi3Lzs3m68I4aSNFRTYX0B3IP+XVTBoi9IGdHW4MtPrR7s0wXfq1I9K8B
nfZqT3hkLJ4Ovi9h3wcTUly2TxajvAM3biKD5kzW1EXipgRjNx6oo6fxamcfsVVWj4HmQnmNI2fl
8tiwBjdpiPH/cZ/x0ClhVJ5bBFpHOXZrtOlbusIQPIqtLO3sR6J0rR3oTb+hl/QOt1LBwt5P/nPO
85cwvCxBVNryLozA5ATA7Lqr8U/ej9iDmnipp8kCjBXtlrjcW+jnF4ciItKwfFnB7CHqi0LZ5gcP
0VZMaO3xdM3jbynUxweCnPV3bwnFW3nCDee1BDxAuSwUSmwVoiRNxc2WHzTlTtLQcrFpavqfmsaR
xZK3UIgaZ8wnbD7SNGY9nMwO7aKCNR552x7TcOk+grCy19g6HbYx5pxk6OkyHcnEVtpvNHSrmkWf
j7/u/qE44sWmN5Nhw1L1MPRBqWM/rf3qx3IDxy6xlzOjn2cPt5wvgxuomyY82sbEGWRs+VuOQI1d
i88OpM84HYf7wzWpZcOLKaH6O4/NhCzqdW1dFiBc2eQTv61WU8723E67L2+xf1Df7hD3p0FsGNXO
Rf8UbF/6FWc/qhavlAn2cqAhfAGWGURgLrdcDvE0eiQXp2fpCvif4ZLO+2vfBYFLQgZzHdI3V9yb
aJBzLTCaMXpPT1oUjuvMkslGjHZRv6nCoUrqEMOAtFliVC1+BtPAbRbg9Qcnj/m7ZwpGZHuQ2nlT
AeTuIVk5NlGrGYsFEjgpqckfknMJLJKryLp2YDOlDUZwJeEs/iRZNIPfmBmuYDyjcdLDynymGlAY
56/7EM53J90F20uA2AAqB8TD2482yc1Cg6Sue0McTDmHJgwVgVvjD4zkjLNi8Nc9qbshA6Yr0ceA
Oy0e2NIaWFWbQx9UEx8zNVCngVWC3jWyomspm0406v+1eVHnwLXW8BCCRi00XtXXWCqaf8NIwEc/
+xh13C3En3B0BTecov4BoE8qcKwINARrFcF+ylaq5LWNQop512PJooai6EdPMesiOzunYujmg0jO
7hAnzcrYHAOBI1zMhqinD732YO6MsHNjvutlMLgMcI9TqoVpK4sdmlPcSDQkfRUbLJkiwj9ELl3O
TYArr41VHSlCRb43ezrmFxfNlL9jIDLS5XkHjeAHfX8j/KRNRcoiP3uOX3j/AbrraEN4RwpqnKd1
GyqHojGMtOpRvQiUowvMSM2eP89D29uqmQSiWt9bOloBCGfO8MNj+lYNg2RHB00dNRF7TP7KHzbj
/ndLdm4v954bjDhuHbjnKpmLjaTRnldNskmurJZxoqv2mT77AigI9skN++s0cYDBeEQj+ZQdmm1/
I1Y+40+/zRPAx0k3IcfxIEocOs+Zz4c0C5ifAsVcH1k0gL2hP+h9JPurKC7Q3zZF2UeHvXBLNxNQ
NpHcZXww5JDVxQ89Od01S/MUeCqHIFFROdasJZ6cNt6c/SBOzQedN+YgiOGyo/Ouot7gas+OleQK
1zrHnnrpVWZcSVoYhfef75oIdq7mxnbNAUexxNxX9tRzoq+fGDS4fY0lGTpjiFr+xHc7cbFKW0+R
SZuR3d9GgrwM2T4klwc3Ua3Wp6ovX/6zVWE7DmUCnY67P/If8n8ZFy+y25B4MPmnH2rEjHHWE0wW
m+H60pQW0bVfa4sDljTzq8GMoFZyVDvlQGwD85wbWSxLjJAdeLgCxk2yS3SLaSYG9ClmLBOl0tEt
CpQvrSBqW1x/2wGZb4lHT3zXDgeBwDooYUtafh29+LTqIsLtF/Do16KIjwN/CCWM5smMAHoy4LSz
gDtiOtzAVs7yWnQRFyJSjJ4lSE5IMPzXwWMq/DUIRtYFjHnUaNwSU+6CUvlu4bQ+5TlKjNOwOnKC
EOs4K1SHoOwdJi1UVvjo+1ENzC6zwn9csEqbpstw4IMJlnjrt2JrAeDdGMmgsaTQiy8uzVavZcVx
LpL2EoZRZu75SVf+32lhwUaY6BP+PikJt2B63Hoa+YHQTPE8ulfg9qAAAWoh9h408namZP2ulsmO
uOoGKmHcVsfEEHJRId01n0j6xdStx3nMfnS1w+XPzTUYkpkuRgkZZelph8W22Clk7jQPJh45+8EZ
VbU76PSbGlgKDu6h+qomkDhSIEhItwcSlqlPwQevwTZxAPLhi7wCgsLSJm9wTlzw6PHW/6FoEqWf
T0PrPIcqZ5zkqJt3ThDqD0zUqQ3Iihx3za0dYBlTn8qAwrGOlf4gnrlv9LVTlvKTXNiv/RzKe2kO
4br6OkCNXw8XMMdQfCrFEqX2pzqDk1LQhCYEbuewcqvgi3x6ykU/8yZdXDuBtlWqux5iIvZF45BA
kZ1g8ueBaC5ZcmNnx3Tm7hDPXetTHgrwaSwIGO2JWHs8HyS1J3r/KsajqxveZ6KQcUuzzrKIWNUJ
pc9nM/chTK0za8k8r5Km29HBa1B6YWUBwRvCVFGHHiaEB9RhYD27K6gjXJ6VN3QA20y2YYjsV/2v
vJSeu+iB21NiSssZTHpfld9dOE/8pjhaiLlwOIodNoxT5L9Uic7VXM6HoQhPbM91aX8ofRFdnMdX
bCNooz02B6sw9VnRQo7oWSBeUV72xkC10i8bfTPE/kfox4cnaTW+FPSvKf6dvk5k82yYpmJlupGg
7rZk9k2uRi8S1tqz2RRcK4sLdNA2EoHlZHFXi7lfLB90fSSi5U5vsIR8n7VemxV8Z7Lr36E7E7PT
V0Q9egFFM3obO1RjHeNObikGd32pElpcp60f8rvJIfzTQfk+tDL1djtaox27kibhEjynIpX3Yb48
Tpz1wvOOM5bGBS2zy5IRNk3Cl4B5DBgr04FNEe0adpZ1wCeOue1MtmrmeqamMJ7Hp9Qxb5DxfQyu
xVWP33O7JuTNwMFYqXmtbc6TKj5uYHeL+8YFQvHa2vs+uuuRwzGH2wL8I6A1zrtazGVopPHzziJd
EAZ8F0jChJqpzq9gJiBt0JLGmx8rOWBap26eyQmFmmOOu4vM9WHH7NOjIjcCoRAnGvuY+vjrerSM
bWvfej4VmMlK6JyshoWLhA2Y+WhJhHmh50jmGPjStE0JLJ4vljy43Lm0XaibsmMHar9oZgkQsE+Y
z0Pf9LOjpv1E88pB5h6CjgIG0gtZWqx/BMpHrzSD5ro+FhTw2QoGV9L9rDmM02hFHQjMjh/35VOJ
zFENuSatDgs2GSlTXinjaE4VsQulKAr9JsobU5sdB4uf7x42vHNqIbWhI0XZmHc/W8cmvH38vUCt
p2q0wFmwfJld4cQUTRnp72PsD1/0LStQEGoNwuySJAMgdlMLvAxyBR7ADuCOL9kS5ntH1bx8dtpC
FQJMKUdGmjBKs3LR1EfezwSq7ZTH6poTh29rwVnMU4Doxzb1brkedlwa4Kup3w5utET4wbFH+cpH
GlZqOLFLaXFa+xsdFQeimACsad+bjWz18Cd25XZJau9Kaxbggj/r52+5PguReexmlOKRC+OMhJc9
xB6e+Ouge2eDmHzYaGEw34KM1BJ6ZBol43M7S4YIvt+eKai1Ld+2GeQbFhkoxY5/gFoK3N67QWd1
+VdRuuwvl1513VbacRywhIlLpDYFXdkw7rkDLASF9Kl5JYUWdRM7up82jlHcawkbSgubgiBBKMsB
3c7uj17zTUEiP017n4fKinrdhA4KuayK8LNVeGP9y63SxX9yq606784SEuMrJ0umoaJZA9qTssXJ
6KMax41jQ7CdDNc7ibD8x6M/HHgiMGyJEnrj0Coltn0BNo4SrwiBYqKr79AIlCFEN9vNo1javnGS
ruzN+cAPT9cQ0zd6MwYe2PggDe/NlpZN1pXVuGEqluqAgJP0rHyKM3bR1l9wj3UMjuJlhiUz9l9s
vizyVYSmnDqB0DRdaEVXFUgtSWK65WXZNspW7pP1A6KmGl/Jxkdr0+ekuBqYmvXdQWOkSnwhDdFH
RMjTtPSQrNjo2r76+eOewLfrt1PA8ngcNL3td8emAT9I8SGInjbu+jcjeyC0DU7q7DAPP/U9rouV
ghyp2TRC4GsM7EtMb+hnDB83N9dTFltPjAIP6KgK/1kdaMGfJwMu2+A/mMQApZ4LjbA2kEoHxSiA
AHa6eCXTr+n57Ym7U9IX5kfx0KcarHPHfSVfyS4Q2JQ+hjbnlAG6n+RNH+vPoahSFKwg12B0o7AH
EKkrDt5XApod4SJ9j3xuxuFGBNnhE5up6CMO75aXQk+KQBnUaKRpajrejeDdVf7lHUlqSZE9Mpaq
WsyyfDQ3a/iK0bW0ELuPbPEGIzh/jMOpAfPNBfr/9k5ebqidIsnDEovjKjQIAUsvyLErcg9z9Miw
WanuFPbaYiapwKvjMzz3vuqIag/kxx4zEobU7eKG2MPD/Pl9Gro49t4qdxorvQwGB2hk0hEwzI/v
g6QtjUmp/k4s0MAeCi0nfyCJXScHXgTnbXTtTgKXleHJQ81OpvcqnizemqN+/343EIUO+38DAzDf
b5iaqu1UMFeRJoW1FIlZA6oyupQ61Uk+7dKXIJsJDMDpyzeXzb4/IpqsU4AxZmWgNLCPJn3PrSlo
p4ewzdEgu5cOsdGmFmRYb9njLBnhq+M9yTYszpwSPuBWhvdqNjG7XLcRysnnCoX5+qnd1y4i3ng2
bywXwrrAvlQPkQDs59dcVhfBsphKBz3v7Xk644ZiTwt9Fw9o5FXOUPwxIvlHAzjozkoEbk82ihGf
yvKRwPV6+pgdJzCnUlYF8n+8aBBJeT7dHy5/Il4S5TfF1/gluhEbfr8/dwk2CXGIxnGloCtOO4rx
ZW86aC7ideTu0Mzx6gf6rs+kD8J7wG7gKRB8evAkLlaGtpamD0mknFclGDCFwkvHDOjfQT5rnWej
mzM++w+o4egQmerdq9SEGGbLKVwBxHoa3iMDqP4XjNT4i25eLorDqlEjXgVPyE3gvBRuzyWcvcrB
P9jjsYdmykx6sV4thebcuEGN7y+adrXaJ+unlCFwRl33OtpEwQ5TLqk53laLyKE61pibRl0+BvMT
QWLdQNvTQHtDJln890SHBYWSNIU5dxndQZ5GnrCzv665hb4iiGrB44sNdqk/ZrO59xr/a5r4QSFU
Zi0bz1DDfmkBCLr59wNu20sOZHA1qD0flbk1JTSIw+l2IzskVK7XifqHmfjqM1YVnZDjWdy85jZX
A8dfBDk5T/yOKZV0+Je/qjw3VdvSNbJQO4S+uYguydfpYlInyWcxjRxVqSkebAhfcG+NgXcxKqXr
2GOgpkYyU9+m3yWXCgzLTPGGLpZUe/QHr+9XrHVkj7Afo3vU4rTxbhmCQS3o5bs320/GR5RePvky
drjYYPy/TKCFXDC2olART0GQs+7NB24kdB9Ffx7B5kW1t3QSICpxxaolgFCZfdfH6n6/99QwuW4n
I0EZVjczlrnISY6vYklGuZA2eZp1HkOhKMRwa8m0KwA0g7PiyPQDms9P8e67rcCGe3/NPmI2HEYR
juYmJ2ceLlKMRDavL7E9TjKix/b+Gsv2nOPhtBKOj/gdFV+hMLh9eGVnTCQ6FAdQAHICjcy82980
3TQj6I0lar+deFMo+Fo82UTo/i1mh2m8dd4cYYLdhuz/SUv529oqDpGCdTdxpz59kijSRI72P1em
fHd6iizF8aulARw96BSGblnLGqe16HSLBqg9EgyhKyFjUZtZWcVoahHH6YiaPFjjtyH13ddnDPLB
atdy6pdIy32wW8SAEDjRj43rdJ/PsogPdr8u8szMENQfE7D/n3aXu6H8HXTp+zR3uK+hwT92bFxQ
3ZGG2uxGWg6dG3IoSYMSUNGpvZbv+TdO30p/uOZ/FA7QykzsucgNSlu8dPxyqq67+ZBqEnH0g1jO
2p1hkoHbN/t4tsDbb9/YXpkI8vt0YBYdGxZgl8IY5zZmF4+b4PuQPx7rOQ8jqU98GVE0Y6eUNxLA
KVBqPTHU270nV4ojM6JhVBRzdY0RatcjcHU9u/hWgSV9locU31vzgK53ajut2c39qMhCEv8nh3dM
e0sGovG+vpPjhDx9cKVmuGLzztOgDZXkOtrNDRVWKQzz81iLvskXLo1tn8UJ5i9gXwYorun4zEZB
5X1NewlyeKsQgYXfwxqSPJ0jrqmz32J7phMtYBLo5YpHXYstbDQzYhXXmmF7m4sE/icarywKchB4
U0/y/B9tU2NwdFzFNSBUw5M1HzULhIYjBG4QunPz0AShcZ3cqzVVm/SrR8/9YvWur7LHUQ0KUKB2
8aYssmr3jL6diWa1MJ8Fa0wH+mywn5OYa9ltw7zpYCd3wNEdoY3x1673JFr480TMbBpH/SgtPW4N
zyAVqiVGyFyh3ADd3p2jeNOYCiKaqq8tkv849DqnXqHKrnG6uo+agKxqvNl4DqTQnezUvrZyaZRV
eLFGn2KpNDcXUQejOfj0xOgfHc+YweWvi5N9SQHXmO3MvddssxGtbb0H5pyOlTWtQa5GoxqjTVeI
HoICCkSgz0sKiF8rkLq9JR4im4aedYUA/gBDnHCB1uE6VcWsBz7x7GofUeh9YfQikqueIHYaRd7k
5tl9sAGdmTks+OQehUqgAN0oR539PXHrCXVbQNfuKGo1o/UubRB3gfGNWC2zDEYhlmdQv9RPhHAh
/ZAxQ21YH+6z5sxbxtAaoUIKrRo8EplbUi0yLOu1FbWz4de74o/eGWcmi665DxMAhUwQb1wZVWQ1
Iy4xWd5kCB2XZg7rXPTYAOm7BUoYpNzNK6ntBvZ7HEp4lXQq1bO1qUMB1KN+a5AzUqbgCuToPvwI
0nyICa+oJVewnRe5hanKXbJg0OnuRdYMslHPOhthU7qNQeU4ElUIzBxPna1xLNlkjYyg/GFAxRfs
cvbrRc3F1SDEWN4qKU3j8WtVX9zgVzOVTUGDmwjzfFfnp3TE917FFKrMkQ8i947A2MS/M9RJS5kc
0bCAiVPfUZuY2/X3ijRRT65EqdEM+XjCw5+r6jQQ087e6BWm0hfRPvyzYf2Cmyor7KEN89hmXJY8
x5tR6bgtb05QLsE/Sp7ZEIMxm9dqRQh1AtlHq+lCPmxgyUeUEMr9uCrHKZ7aE/0aORbfv/OxBN8g
Qp6YNW5klqSpx3/Hyaku9nLCI8nEda4xNZUesHoibtDcl0poFxi6WsUEjIFPWFt4hjXE/NOaEuVZ
Fs9fdihQlEAo+uJsDoemWs1O32tz5lZhfqojyjk1EV9lmp/gzvHAFMk8NqCPgcHQqIRhb9w1Oi63
GF5riiwWTZZZIaq4g/Xsb6kOdRe3a3xn7rhJHejbc6A0Sc6MZcSsI3+ZYnEKQ1kMxYFTcRzIqArD
ifSyzCIIeqbUKNXMP3NeYt8WIJdhK0wYcZT3OPv1Uembi2etoBBSemXgZYnwSfvQPAJ9T3q4wrzH
BmsOgulX4xASmpBYg/zojkiqwuv8AtZFpy+OnTuNS+nfJ43aSfIkXSJtURiBuxs7Ba4A8iRHfP3s
OXe1O4TRS7K3e9N1tmPuBGu0uy4s/y0j7NZO/K+8R0D0OjKmNSeeyoMyngXomUmTGsuUpyVWYdEj
8m8fpnycErbKYpDKaz1ulSTqwM2c6/1mWzIev/gKsLQFbfkAHN5uYAdzXUX+6SbzNtRpZPW594bU
ypFSqcD/8ZPAHyRIcADCaJySONttcQb2qliRH73Oo86J9l5AOCAoWdc1IfBtF3l2sfvvcSBaP83n
bdipcBw0SnVUPxZRj3CoVF4ng7+Cpu0zsmJ87ka5lx6kvUdOYYMuPlWCRD2/c3FjvAeSkIoJJKtU
o/JrauTzQgCH2k9zT4KjYqy6HilmBQtM2qgPAcHDyakEDO5wNzRnxtu9NKpmESwmD2Ie+yZnfon7
ViCSKg3PHuXczZFn6q7Xi6VEPSe/53TXOJQvNyS9VwVXMTO1Eks9H+LIEkLas28ij71zXDkPhwT7
2Tu3Ymy0zG0DGLB1bGk4/bQP6DVbJFYz2qkU3mzxNjTT/kcxhGidWLZ3ydYfuW4to0FuZYswEZx1
vw9LFa6d4t41Y14EtDerfGc4w0HYRaMJPZIwqgJstUymp4iwM2o5q5ilFZjBXh/By28RUIl1TJxX
4OBLS9FkcBTNUpemdCU2LXDJvuRunq7avqm6M2T6EwwVyGrAULZDS77fvMYJcK1qDlrpLGzGHsO5
oKXQ6tyylc75QxJh26/dTCQ0Hd61mavCzqkOZRc/kbPuAMbURyWk2OLGAa4qDcNz+NGmDfnPYg0E
+Iq2nqldLCiZYPmof0MTGaHlNub3TynCsd/ZQe/oeBrfdw8IToHUg+rdqbWCN4t9P2DjS3sROvu8
HMk+b/akQQQRpcSeXEO4YMRH7aJA+YjWqDy8z4+v0zgs98i2ea3vdjyz/7ppxxMDuF1hYwWSpk3p
c00r4XvmNcUCndlGyTNafMt4p50zQuW41wUAS8VzDGsHGBTkZ073U17JlAxQrTv3h1l94S2c0GwW
sq/ZP/CltsPBm/wVAHWaNmDp/j85kikUluAUkFtQCmafyemoXCkvjT5Qgx28DFrTYxE3afWV9oly
Lo8B9B1o990W9XHj9up0dPzY/qvmlj8ehD4Jv7YwnwDY4Ekqvhyit7OhIBw1T7HpqcMxWCBMJZKh
RUH6e6fukZ8jSw5+M4jC7Myi/TT3giWyippz0oIMqQSJ7wWlqLmKuKLVL+xIZVXCkQqAsYTCepoW
ihhiqATVl9Xr5RTvNrXDRWjOz7BmhgBdUOM+x+JIHzjOO4lZDxPO9c1OaCJiTROrxoS/QCZjvlfo
a1RQucLkN1PMd/mjhb82d47YhzyDW/nILqgqC5JPQlKlgkHeuVOGZ50NhjH7TsUnVYy5FYOR1ZVk
Mbygj7fBIzTVQ1OvRnXcx6IJ5u2RRzvjhw/SucISdKrI97+CSCslyIT6VJe5GXanN7XoEVm67vS/
cIanhEuotfEtGOtx3J1shkg5A7WCBfcCsLrK1sbfKzqncjvfYVqkmUjiA8gh4fPDHFOIS3yXAT42
xjGhZxAyMtBN7lx0jfWr7kqrg8jodA2P6VrMBtCY9522VetVv3mXCvwgWUSKkWJ521w2OaS58dvY
BPSC76jbl6xCB5E8JVyRSYloAt9AL5ybEys3V6YJhMbWatHCoQUOqA8tuTIwJuwJY/bcaAgNIKAp
w4avMe880iIKNq+00iJCXtY1tM/e8IrzlO29CmsE3JUI+2Hyp5Bl2WBtoteu6m9cXNWUQVVbmzdK
OX70AE11Vg9SlghokeCV0cVD9jf/cuRU5lXiYmUqAX6So4iqPpv2Gr/ipfa62t0uXZBEcoUWGSQn
v5lSAOY/HMJTo0TG5nFwU42oi/U2sSOoP9SuF4U/vWttM3Ar4U4dF5BYoHCxTd7lzuE21TNubIfv
yjf6wYdvixamTEM171J+VAIc6VI76lCiPdFCC+wrsVAnLNPvmy/Dc+SagPyixetNelSDRym5eBEz
SLnY8u2+/VMP3bimc7bW39729rK0S5vltBnGRmDo+BpaCnp3Z+dCGxzEXqGjP0CrArbDn2wDdUVY
AQnChO+X+hCs6YMh2FgOw62/zwXSZrJUKzXkUMJA6kstM4YcopNYKF8w/7cKicjkUIdIu9wstCOx
m23rOybvVTwwYWXLxADwsbUO4x+tFVVL0Y2l25/z5x+SoulmHbSy418j8IXzr6ELgxQb5Pjd6cwH
TBCZnIxbt553ORiD+V8RqxRYdOYrVtESt6RpDAuQhwDhCiJbc/9vuSK7LUD0m3MT5VMDzEJIdL3s
KveriCJRApZletUxnvCeZdcBSRb5GGWlK0hybyMk/SVr1aWCCH1H9h8krvfi4ueAf52gxERFAmab
pb2Z6CHbLSlAccx1lvx5pqZ6j3GTKYCyG7vqewHC7sA7Q56xODis/USt5bsRGCaiNOJ7/JGgJvQG
lYq/aboqBlwq4e4JvEW8SxT5woajlsA3f9tkPUsLrdEuJnbUhb4Z9ixuAv2zDFNiTyGitY5yUUuk
IWikhaXsBpEnsst1+SyC0r/Wtc0pj6pydcYpNigLUi9ciVVoL3ufmKDmyq73TQRXGOlodmDe0ByW
BGBRWK3d4aNWoTU1HL76St7WuIMmvmHxzX5j8dVCvX6UU7I7ls7jHGHax4IrNW0KjUTkJkHTURAR
y01aWE/qEsPvqiiwUhrl9CelsDlAnC8uhgJ+IrM5/3U1oOMzvefZYykXU8mosRp97EwhA5bkQRVN
T6dQakxctP4dqgIX0u7f36KjydY9Z2bdCZ3FRttrOwmaXi1q3SHK/ElJJh4mYA51pOQmG27l8tqI
3zYxGBNQwBrv5zD/8X6WM/b34kxsgchhhcI18fI60wZRr8s8zFk+wBGdzG8yk/ZErGeHYWJARrmw
rQw2iZyl1g4P5wzuibld/x9aSW+wlwVSC1FdIr3g+Mga84Csbv4eglKCRghfEacgwImq3knLZidV
jfovkcBFoBsTdIQfGWRrw6IyfwlPSiLGq2orJ2bgD2K69HipkuJDj4iDmBElwRzhN+g4QGTt1dfj
47rj0si8SgNQkAw38yAPYBrTZDO28wtqfSTCwB52qfM2M2SBQx3dz/s8j2vr3zoCfjHEfQIByUfX
kvEPDDBevgmR86Ubr6OZlhSxFEH2bbpaxQbvAaA2/EU/qJrkoJ1XwRYeRJfVVDIjBxXoknkZxrNT
URTfZTg3B9YCmroJEBm3OLFzcYNP8+HKiWCDK6JC9hv3q2b+qgGEeK56IasGLF7+W1VTgAdQXQGF
9pMFolXBuD4quik09bwkInXsceEwoqN8pmen5cpjaMMsrsA0cB2sItymFmRJ1lW//YQY3t5USXh5
McN6unOmsLnEpvCS4Z8cWUZlBf3pU/UcBSWmAOYa72DJfAc1bmzCayM79T3CbrfCksFHIAxCSqcC
t/76C+xrAOvDi2BPKkstYOLfabc4FtiC9zEVD10HKK5VPPcxp1otNaflCB/gYPj/jgfKHJE4yJz/
rE+fB/OAQVA05BnPcthQ9YMkNzIbvi4HKtvLJlCA8hEf+7jZI/MYHs40uKoUOUTq+wTTV2dHrkrO
8bkoIIP1eqVQ/8XFlLh+31CaqV532sDaKIHquR3k/lD6BBIrVIPjqtVCfM7ly4Nc4ZLe2oHKLpL5
u4EMrNfP0WahM9Br9uLE991Qmf+vbR9Q5QFSki51N0jwFWSc1WhDDQMjumkdYca317BAZqDBFzwy
TOwjYZ5Fd3A9fWoS6oL7z0VSiheVAKFtUhXj6JUIaZp8618r7rKhaot114nfeGmVruGE3/dm5r07
LoAry5MS0eVEy7rk4IDm7SkTwmfoyrNvgWzBvTSkObJsLIw+3pB4ATCf+BWakuf1SpKnDpVsdUsq
6oFBQMa/84rWbuZmVGEl8YLtxcuVcn+JhK1cb7Cnf/Y8jJuq4E/q2L1ec91/1cT9Je+bJVxvOaK4
vNGUs+SO9T1Lok4s1KTocwxsWRIz/PfWqg1XpTdMpyQlz8M2AMUlUD0jIttaLd2+j+gQQhpkRN56
DSjN+g/vAi06zZBCVxZ/1u+qX6o/yADN3mZXKEf5EeVnxPaypDDjzhqbAzAIYpWCSIJzPOCCbZr3
jdzRrvTbdWigkRqIhdP2LHk9IHi7TMMMfREu6l8NnRIOul4UXgmwkNKbLZkPA2SGUoy/eeMWJ1s8
SDSP4e8dqwsxicsftDrIAUlDXx/oVx5tpQ8N5HSLpxwsdbaEmNdaFP0qJjJfPADnl26SBtg8N8gc
ltz7qz54wRUc3zNSwHRGEcvg8DvRvh0Bzl1Ci6awac8Bf9ERK66IRVL5Wx1jrPPE6P3MUKAEH8JA
aJ6k568kbzbsuLAPWKmXy/v3vVtVLyjxOQQPW3F5aIoG2kUMQo31Gk1BY5leu6DO5oVOds1OibbW
zg8fV0WBaXGKlfoGT2qrjPHNPO3g5UdIKuvymUyZ3CRPcGmoPzftT6sTC/64XIeLg8ZDlNQzI1kh
8/Obkn4Jsk0m4N6dxAU1iCdcaz5Cn0G7Wjzs+AyOVxmSNnHeZlTy+LVymYAbAY0R6Ub5QTeEVQu8
tCQOQRs34d90/63bGnSJs2ZyZkiwda+kzslKC1B+vfyBfGjfXQ8k5fp+Pf147AqEk7o07KzhBGpq
wEW/Cizg6YIClGhgOAPjA0f2jxc2JAPs6chvL+lx3RWrlMQzyPR/L0IVxLOaKj3MVMdnmw2nm1JW
lpCCNuiC+mWZhLtAP/eUGH4Jtt9pnYQz1f0Vo9o8VXUl53+Rg1ku2kg8LLtGFbWxWzpPQxomQdpM
5VyN6OfoTGKoFY38FA0MJblNiRpPQaJONM1ZtwHjZz8CSOw7JrJCJ9Hi4yUB8zKBvD5umf11rGqN
wpUONYzAmeX5escjyicGGScGOIxteaYWkrQbOOzmVGj9FHmiXW3VUr4kPZYuwE4zmRPgMzw90NjU
3dYcA69adXzD+424bf/jzxMRtmwSgd31jqQ3tEk++tmISIjwPSNBtN63ZyMMtaKtXr4cQzGUXlhU
Hd3w4lxVPKZfygqJi2gj97fPBM/7d8tu8XlW7B3gXgtRINgS1SNxK7+IxqkCr+lTj65HBUtSvRtx
CLq05yu5LGBGRS9lCdXeOZzWPryF8ECdVUU8B5Z4C+SRREWjsZJyF+kDREvzXohHBrmngm2Y5+/N
O9xI04vAf2wvtqG2gN3brlwlNoJEFMkRSH5r9HfrELoSPab15TpHP4zYwGdSB0pyDmMTROAbJhXP
cMifs536Eih2D0F8mLwOa4qEZ2pePYyBZVu65P1sle76bd1K2zHXbbDHfvR+bUaV0x/SxGyYfclG
i24cjOlp6otZNbX+hb/FQ1xQM+ZMlBhTVHUiVcz0fgBUEFAYvDw9X249BDbYA6L8txIOnPKj5b0K
1AkqFW/Uhh+Nx64mD5jPFcnhu5PPhB+cv0C78oi0RAKpH3261B+QlGL4KacqmmIcJa9qGNmByPKw
RlGHVe1CbSjA4OLOHg39xFcglzBkNyVtcof5icudcRdiNc1v37wG5mq1BCYhP5z0vwgzTUGzCUM6
wLtpstK0GUK+MZCOpJ4siXknoQxH1No7SOPHIc/9EvfFQd3+Jn6yu9jWb+8UnJsl6OKgtaqtgkoL
9dtaxUZsbTS9Zv9Zobc7JE5rQt6QIoBx1+9xgqv6DMjIujXh32naGNKNFNwQffNQLplZzpIse/HR
lgsRC+FEi+VHm72ro/MBykdjvutXATmWI17DoC4WPlB0FRV/hygVv0EUhthy3Aj6Ddh3oCORi79f
H1WaMegDp599QR5LWuRQQ6wA9qMD8ZM3Zn1eGzRUVNsX+HjnGCHJy86aa3IGlPObx6axpp3UK1gN
bSrjSSN+93OEBkVWvmsSmmfSpHjSx33xnScX4GGjTJT+SFzmMz6SwzsnKbBsuPvHVAlF+wGARVe6
OF/2oySi1TvNT/eQArWlksgoielXVBhOCzEpTs+1dTpWGSkL540gZ+mrpECYVuWd5D+12/dLrPBN
splP0yX3AnnLKaT67/UlHaqqVpkXRXkGcGAZuUsTIG5eWT/QJefyA+17zmDSqiT5yZBHURmah/P4
Y/zBbYZM0qDpsMQRjTUIz4uckpKs4SE8XLUC3SY8zz+/NJgTYxKwGFc/eYnaV+yseRfBlnNJ32MT
FACHbaabLHKbd37GGl5SOlT+XIfl56nM5V+ICQqrCwyy2r8+CTCoik9se0E86kV9qonII5EaIEhy
2CGzgysAiIxuFLs55Pvjh5FrgKUs21/hjabnQcoF2R1IItgjxIm0CqFOM3Ob7hB4DDE978vdKV4r
kyvJNmZqjpXQNYhxC/qVq8Mz7b1w0oC1NwR/GqA4aSiUyOudxtybDHbhUGJ9h7eAYZmfMhRBjLnL
ANfl4gQMPxgYgASVcijhPMTvvWKnlHUJQIEDlFGugadFBzakdP3v004pz4/zPhEptGZz76pc/Tt+
gy1+HJpkkwMuKXnclaGz/IO+2y7/6acAzD0loSm1Zaa1fkYu3l3hra7PUBKfkrFie/HmLnjb5Ven
Xr3rRhLENtY1t7vDCIJGber64OG6dgae0U9FhDNDzAFpvIy0IJKm5XHBYC3132jNgU833bYfOx+6
IFGHa35BKrzPpN1uSJHknzOCxAwe9tJva/4cJcTay/9fqglEe9mIq4UqV4Qm2EWxvtKdvHNm4G1Y
UxQzlq31S0rJE5e7vow29brue0gNL7RdKDQwgzs3XP20mfxe9RiRVoxIT1AtrBESGXNmcKqvdZh0
vnvMNm70O71H29NYRtO9IkNTUblREWqF3r8bqc6hqSd268jgAb21F2EYxWTNNyJknI7dBcuiIhqu
6rDsWmjMf873eERkmz2+9WIiDehPFx2zW/8WfOJNOn+lTs/QbRFOoaoB54LoEwy2KtPtBxfMWi8w
8Ldhk7p2etkNpYJUnzFlvtP+If/Pbr2MPpC8QQWQxzj3T3/S5r02hW3ZRAkC5DK8Sz1OC93iTB6T
k1j6+Eby626/lfyulJATu9EF9G9FzHyAk7qM+WjS++ww/FFziwSTRlRYbl6VjYU56/ay3ywBhFKj
BYYxdJ84CuZVIGBoag8P4Atc2GOlDz/ZRa0EexIoCc15t1LkyLrFzZtYNriAGJs1QnFn31ioZUXs
PVoKbRKrdqpBmhqqcLKmQFQN7zFYzdVe+feDQv0Mu7KBFWSrM40+DM34mNSeQ8oh6Kykvnh+eB3X
D70yskCegpR9hbVkucZJg+PxNN5KKa/v+r6wGbJ1i1Njlgl8eL78YR/+exp7gC1l2mNbflXmR5Uo
w5EIHzpPDU2f1fx04RBVeJHUqpRA5+B1WxqHuUWHhC002+PPdpZczr93Npc3slTyEJzsWYAnfpBn
sG30QGaWy9wb2orAAjOccZlG8tPUBm+Rcd45XuTugQ12xpuiml99cmcbiNbEdCxwJ2S5nk3Z+4Re
N6cj6bX6lY2RvbLMRc2R0mE74ICDH0rVlFZGeJ9qZyH1gHTHhWtV0Y8yBjsH4zNI2kZcRs0VJgTJ
nfZVSiIwe9xBJxuL71mzN2/mvUAkLPLGfyfNkb7f5XhS/NIbCbY5F+XxZdeiErYii5Kcf3zmzMLM
5cGRFi1oEadLUKj7cQhjdezV3j/aMXGLZLiRV9zyZzV9WOVqj2e2iSaA2qysT8loKTLbCUOE3SYi
DHP9gdgfCQi6JArbpV5sMbGcYS9kkmsc8lwHhugDF5LJz8oDc+t8jO7fDHHChLHRmJO3inotTuz1
RWUL50Y4FCTMnf1d7nsntyYpiAm7wNvvLGwi7acsK5PLmHXbKpNjHHPLZKU8DxZgg1vDpaDkf1yQ
pjPmODur7TS3TDVBhfuaGQGpviLBBlIFY2q+fN99cOhayIGMIL/t4JreKDSep0ktj4nWlzpG+yTD
BcHufkN1RN4B5AfApOviBLygOXIqlJPWLGhxGqmwjE6Bw5B6XqxaJJNPRJY2xDo2Wbyuhyyok/W4
dVr0AwrPWEcyQiN0HXFsZLsFl29w50i9cFAomE9UrKUqXPw/UC82N6jir+enu0zPwq92k+NsO4ns
7oWBSdYM08IOsQIkn/ezp8HzfiUIJTOAIfuuE4yklo3LP/hMdkRoJSawp1j3XwWkZWz3tnHHkUds
JE/mYnKV8xplJVDbJraZr8VslhqKi0CejlLOZb6i+7lpmXpm7/okC5NaJ0IKtPX0GMDjcfeZmf8f
VcPxBqWz6XSiBmmYKjqONectmywNFJ9UWMkxulZey/DigW1IAsM/uu9zOnWP8X7falbk4DsVdVpU
KT7nYx+PrsEljuZVQYM1X5eVSlBTHycBRIupI3VP7HyWlBcl0ChIBIy9yjOAp3Cmxs6/AUtH8LXA
VXYrry77xK4rR0OzCAhl6b1Rrwucp6lz1dn8Iwe9WJ1lBOA5CdtpmWFa5zfqy8nLw24HXqARxLcB
03KnGI772Qvc5tpCK51RnBbSL2s0YfLwTANr99ltofDNljO2UWt0Ua2SuYzzJk6+8cObfauUAGAk
e++8JJB+UjnfXf8dCuDftLbjcCEwl4zp651Uny7surnr5apStljpy240Qah5HZl2euhKir7YtBkJ
JvUT2EADgqUXX4afeDGH+y9V2Ro8BSl5nRdyqmfp3ntmRYwTMmuL9g6zqongM/pqjqb4a+illgTG
8mpKgzydcbqT4GpC5SPl+PqY3ulV4Yg8djmcP48pQ2punGM3VjFMOqqrmG9Io4/wNRATrXcgwvWH
W00ss416MVOcHM4mRZ21IS64AvwJJhsg79oDK83BCu67YWdYRuxJFNzuYcOthDo8xs0kFktqM3mR
QTTmbnQKbCKEis4VKx6oI0NW0SgGiLNqiD6I+GFauciRxl2HPrCDXtBpIRw28mm+AFWavB0hFWye
VBTUrYB/4rZkkjIiyXOAAXTYEB01efsHrQ7Luwr8x3amEWGViUXy2lew1CKGouP3+Rt114ezX7+G
o/2dxz5qR4v2+BuphebfqziCjbAR2iJF/2hBrgHLlfkC96cOu8RoXXW5XVZSQC277MRDUKsjB04j
p6ISyQMJgJu+aWd7Oek2+t4EioCWKUPJK8USLGP9YNxqY2ua3m8dLq6ZVadSffiKthbL3p5NstxP
mgNUmvRjVYejTNmlHIE6hWsCD6ZC4EhjLU30Bm0G793DTfJaNNeCn4ko+3P/7LvSnRAMRf1zXN8b
ZRpa+cohjc100R3xzPA2VHQNgdlRpA+tcVQUzU/HMJ9JZcDOLjNsGT/ey2CaY9H34O+fY+gHOM0w
mIpftnvLQIUUqHguAloAQomx5Z+bS1Sixru+jODSQ2iIovWbARleG1ogvLllxDt9ThGmWDL1VuOu
J/cpv5JmkhHQeibdWkWG0+YmmkxnI5MQ7yqDnAihODzW5Lvr5ynfvIVU3QHgrrJVHmt+rrE6muwy
Pns9Lqg2hqpMq7ko78SBdCildPCRWM16QQ1FasL6tzj7AAfiDSZztc3Kxp6sJmt4ALHdkz0dw4q+
P04EnJgLXrv9facOvoJ3D6wGTJdj1b+cyn9KObvFYjR6kxUnbD3m3w6ov5h0+301IYzfiHiuH91q
/rFQHFmLaFgUh1MfX5NL7x4ECKOxoVsnXdzYmUFCLpSey1eBC/RXJnUKqI19zU1IGgh+N8WJMjq9
LCRMRHDWKMztDdR/Wj88g2mxB1P+Q8ch+aoJv3ndsHF+47X9SToCEAxfokWLZO4RoZvXlV0/3XJf
RFuEmNMOQb85HUJXaoAyGsSuiHrKND9QnZM7f75HAWQaOkrRoYK7BSqJbdxF3LtDetkkVLyTTGqE
cZmsRsyIw6aG1r+HrPNYGxyDT6TlmsyGlgQAHQ1iwp4lVPlGAx2MDNUeH4uwSpGg/LDKq6olUKJJ
D5hWgKbhaj9ytvoSoq7GX0YpUjPxQLQyN2BtywSY71wxIBceLCk8iyQgWrkPwtCY1f66oYSIrmGn
eUYw4Zd20xM7+GbcaGIFcN8j77OtwYjGXM1m9HUf3gC7MXgkX5xL1LsV61yj1hf5xu/u75c2Q0V2
fqlVdfR6ut30h8gR/R1vuyZj8XqOoCb1CbvL1IyYxPeTa1N5mxyFQiPrkeSihHkZ7w2lHha22S1J
YeLo7Nv+x5qdjSt7Kipb/aI4ZsG97hf+HO6ptEf7+VdhwfHIZhKv9kNmzNZ6NUu4mOVy2fDA2HlR
tmHmgbf2eDlUf0joBSmypILISbl49J5WD0uvJZfXPEk9c9OWkSarpE1AHT26/aN6XOZ+IxDY/sIk
tVMiGI798LdVqBeIIuQ7DOzmbTRqlmTUSg5HNqa4Q0Ktr8HiNwCSpHtVqy01mlWzkvYW/tX/fb5F
6xuU2wHM+pSL8ANFDqgaL5aJSizrF+hmg/gQcZPjuXihd10qvCdsvulfyO30X8YFkkuRUhleWkJp
ZtTtT1fL4NPr6cZmrpCBBrzjL8ZS4ucAu+PyerlSblv3Y89TVBqFvM/oBFE9uGJ2Sms6VgkSSlvC
7MiaEuC67mjmfofuOXZzoqbiMaFWu0EJ4DmQysnsZifTnZvxwBuuON4B3kRVIUIN4Ty5TtN31rQy
mAi1riJtyMmcVNZ97zRDz0fxTbuSGokaJ6PxPIXqVOAUodoyygx93v5uE9CPDUXHfOmbclji9MU4
qjG2BfZZdz5uUwoCN6McGwyBGBgiSrHZ9uyaSwzdo/mW53j63rxUJZEHmKgw+nYVHVA4l4GY0dd3
x01PJGCl5dSl9LBo34Rj5FZu+rj01yHz+6Z8RDVCkq9mVe8gtbP3ulql88/lK9QIe5Di8aJAbr7+
zq5o4Q/CAjrbgpvsKb97TCMKxESFvksPBCuxc1LQKBBPKm2k0YKY/iIRXxww6cEJd6gxOUE6yI6v
lZhTFc0+dhqzqjcjNpHlzkaLwOifJWupnJZwfPyBHMHNsEkpwz+YEcJrPYgHtQ4IjWQZMbr+4//G
CxTm5eMFwG7sT/uocSphb29ZyTR3YvUUNu+99uFW1RPmaitan9ToYo3n39Q6xscCxHQEUUWqxmbF
TsVX35uTT+3CaKDakXhYSAnHbz33+BDyquRG5fXtbcOy+Lo0MInssT51vdC21iMd3gEanTXxSd5X
bCCpZakxlgB6Wnn2Ta86SMKo2ekyKHczzFT2zje+BNI2Oqoi8WqHmrXu7m42vr859xNIWvfo0uco
6ppOrgH+N5dKjndERSgsuQbrypiyJpFTWZIrKr3aoReT8Nhf/EBmyXCGxf71BuEAQLr67eSH3qgH
gunuSYxVZU8sAzDwIs4R21phCcWdqvNOnPUd7wHLra63ASvZ278lRKFkL7KyzTQ4Cbvaw0OP8JcX
wuh4mA7DktKpNljX/6s7wsUOZgLH9Mag+U/W9K1TsKy6+vF9coF8B6nvqcrXSOgyqniz8A4/kTpC
s/0lYYTBZOHPvdJXefhwmwlgFGx6pwEnOhhR+YduURe0gaNrkmeo8mYmqUSnWozP49r5zAclg4kR
aTyHYot7m2g70ACYTKuHABrWVhoF4o2dJ2olFwUEQ9uQRfrEwU0u5hxMwje2oOOh97DL+v9zk9br
b4q/J6yO/3LUi1v8t5rVq9c4cqXHtTXdZ/mRWDwYkCxqS2UDHlVrWoGpXq4rDo+Z23Khcq5MH0Et
D43DDEQhpPZXvtpNbNxPFCTWboDsm0StIB5ZmE+0qKlO+qJ3uqyrIxJryeLX2VlPzw3wWiibFE6t
+3HUlQ/IqmiB7kUvztyvTX8PXX82wWHBr9SbfyheCjLaOEnFmjCuEJs/9r7DDvjqb42DvwDqC7fB
CSpAHR1rFQdIULn4XmOE0PsGcaSsWqYquk0VlmHzdx6rHoepWIfaxmgYxolzceHWOrbN4Gcm2beR
h1csJZQMoFJrV3TNX2fxE1mXoWjwbiC5s3N+51CpmVEm/Y6N+O6jdur9b9voe4sJw+2sy/va7eTK
/H73jJi0nnc9HK6tcm+TFMBEm+Skpf64/bWpuye4T/8tSaOJOkxY3Mw9CjBH4zrDgTAG3U0IkN6G
jrzx7fpnzMYJ2Lzw3+NI6TPFPKMd+Ly05cMVlVzjv/QEiSxZP1OrXvGe2qWMkobvILiKYWy/QeRY
VJ4iWEYi5JcWPtkWnhNVCIKibbpdC+Wr3+pwZH/e3azsrnab5xDaxPBw2F74h0zw+MzBIeFwl5Cx
NCI3oC6JSgCPi77ZVIPzNO6yDmrO1ziyP54OeCd3q9pohyF2G/0YKfJp1Mhifzp/hyxlAE8Qth4x
GaKOgLch/qVsVNPmrnxyiQK2BOQOrAM/qtCjMl+oeImhGht8CeWw1hjH4Ek/orf3FS6KdcVnTjZc
wRgLxkS4m8TyeSej99AFWfy68240OuHSj5EzBZLlvkXgKvCNzdLpzUCoPbfCVWpiq5jlu8E6LyXI
fdMJUUuJtPJRqyGtD3YRU1CiL5mZp1P2hdB410wjd4IIF3ZJGArLGataig0j0rzEgLjal7y0c9I5
+xWKbVyXoS5ZlTtLv0/mSb4wlk1NxKx0IpI8LMt9P1/gYJf1lzod11lReUgZjDsKxnftspw9deMJ
y91dVZbbBYmZC+1vhCv/EiqpFZDOMkeKH8dKLGKENXPFZisMXUqBXJNjvW8qoxKKUbXqE3iAF9zy
ihel16fcvITISyCNk9XVrKXsaPNp0PgTYvdHfPy/v7ZypRDg5FaMHe6LL//QX6hLP9fdUb4o7klh
T+KAeLTqB5WeEp8u3B2j/HVrB0MeAPuJLQPtC3CH/9SuPJJ/GTSTG/MPvIXe2XLE9cyVtmWO8djX
Bo2N1ITXx8r0xXYZ1HBjxFtqePlhEpXQ6FLfsS9o2RGxrVObvUp4SvlcZX8V210x8OmMZE5wwUfX
fbitliyBcJfVm89VTdSBEMl+CUHwQOc5IY7lLYag2bB7lD0Att+TwpS9r/5UmLWYECjtggZXKSVf
7N81f3h7/diIlmXV1r8mfnLf5dbjZuVdGHoq3amclXmJ9iQiFiWPr7/H2i2JlMX0SfPpxf1HaCaI
SBazab2GNKEFpKAut4p92qwJcWh7vz7ZEB9ewfR7fDI44igolF1KFTFw14dBX0Wk9oed4safDGW3
xpitgmXMNz3SECRS3ZTLU+Om2AC7Ycy9U/09a505IoLLmUu5AVAmRBcVGmNLka5cvPjAqEjOvtf5
a+rO1PjgzSQoEMKC1qLMjx1ZDR9nPWJWGByMYSYCo3oHNBQ78tksGtMSw/4mbXgfWCkhrKKj6idS
GJt7vPZU3C4ZEBNtyFr5hjWzsnYpmqqNPCDhtQqNI+UxLvOzI12c2/JzZA98cThEQjO1efb4+jSg
b4kmtvEq3azBZfDSYWQdvwyEJJ57m7v3JOiUmld5CCkzAnIa1mC0WGHjrQwZcSBTCPAXO8RLSdht
FvtfGV5555M1MMGk/1GvQckI+9Xh55P54qq36mIig/NEDr+4EVKcHkqaKWDx5IDM5lyE9chU5lRg
RBZ5eMeth9YdHSAiiZ3Sjou1nv5aQ8Sm0mejUcusrnehTPwemqBfpS9B+SNVzLek7NR5sQA2MyuM
zY+LAWsg5r+sbK2U4W4F88ncoK6rvC7UU1HiSXdgAieWYYNcGgCRBf9VQhdWWgwAkOS5SQVhd1cS
DiePSsU4VN4P2+9pDPhPekDOI8es7QwjPvGnhl2Jrz1rwm5CpY1Xfny8JO32goRqndC8CCZ9oyAm
SlPIm/8DsYXn/i/R4YMHlr8CR5Wi0378eIRWh1kquxqfzsU32Vdqq1ZwsJpz6xnIegDhPx22hn4b
D2x8iV/aNDaw5e1DaaEJ/9uG6Iar828qs2WAp+R/zYNBwTggNpHU4RhgwDCkbGQ0Ws4xTVASq3bs
cDxFpKdy9CtrVperM5a7f/bMSOh/N7fSv6e2+S+RIwLWAbBao4hVsbHphmpHp4m1P38vvqqTgG0z
3xq3xG7T5jS7oHSbmmjtseylSPzBQnPw127fO55naCmeUrMqmzHB6+YXw5iIj6gdgNneLcyrnCBb
0vQZTrpJJ0SiWTyMs8QwChI5lepTa/WSb8VFlwKVdhI3yUKfDc1qBCswIlMbxBKFEoqJmeto2DI0
UFBzw8ts6kne1Wip24DZyKN2RtNft/qPJb8nqPBt9f0NkgkedXys1H60UVAMf1Sa7pM0thzUDONz
udIqN8wYsJG9JlQXDjBKoad6Rnff6mbc9LLBkplw/DaVD+F+VqoN+BMgeNU1otNXHqNrQzONh9G3
hSt5UYvEiE4G4AmhFsBPffGC9j5exjhRM3K63nZTr2gEE4xBbBHk+CnO1axdYf3Bf8zQyoTirVWe
Oo92CZIKSzOvzmxcILNUO05g+9EvEtgg+QHz1REZ7DWLRjkTMSZe7q3S78K2mEemXKuAHXvdfL++
ICp7K/eGkC/ostI+sld2DROEW2JoNVk1ZA2qEfdwR8gznNTYSVz8FVF1l+WQClCTgTjVjZ5FdetN
JARsrl2LqhR+IhCJYvBMMWVG6yjNgnFcvpflA8j5oN+CRBJ1qzAV5Hp/SZI3A19uHwna70Rp2hwA
mNOTxGYZISRUZAW/Hw7eBRcTldui40TDoAK5f7zfVnzruwJSpFRa3frQABNGSDu7h0Ca01pimIky
oT0dBwckW0sbgO7DiPb6y+KysM5rZUyvzYFfC2cdWXjO5ihIHIpgxeuBHKnBxYIMTcyeBT0pm0Vh
jX8qaoVNUL7f1ie7kseSKsbzwy/uxepQrAjMxvkmYsxPxsDf/Otsri5W8yHqAbhP2YuIQq6dFYnh
OVoIj9Az5htgkPuY/BJPs9QeQhYbrnVMa9A4XcSn9lY+hIRcKZ18t/yEvCsM/0bdeBMNeBvnu54l
oaKdUQkPFvYLco6g/YK7nQKC4zbRXp2/neXGqlTKeSGJ3lMtxY3LBfa8X0hiVWhP4FED9rdmR65m
puzlyvnHxe0MI5UHbnpzwx6rLjW/BZbUhoBwmmSe/nQJXb0HUkCSGdw7vwgCWOnq8y90ylH+xF09
vwPsI9Nnwo1cM+z/CMqf3OINZTqOnHJsv8qIHleKYWY4vNZ1sCdD2XUNrUsLPsKaXlH639ewMGR2
efJl+RbVLly47JEIUx5sR7lIcCJH0k49xaS6OnbI71BUT4e7Jov7qaHzeYLjzlb067EFHtgsl9Rz
jR0q8Ds8EkP9B9/pZ//A0qeOP/ljL15gV9/ij32fHiPnflaa7ihYNvuDJegug5ZAv5CHBqS2Ouk7
0Yzj54wENwbWg/iQbT3D5eEhpyRuW8PUKCVOyHRPFLqsQZ68qtoedvy2yQAqKejT2zq5jHRkShfq
45kA5ukQOOnQOSuOW0CIkM+iaBuko1xQDgbNhKNfTT8jZWTnOdJJFdnVAG6Wg07mRglaAbUzWndt
Qkyl+x/j4+HVaJe9Aw1nt6/vFTZpIRFiDTDGfMz3RPiMfpNEtn64fJccggX4cwm4txlbD3rRXuNw
hWolZDY5frjK+ZYh+ghtLxuulw+WZftcZHlSOGh7A+8rYuD8/5ahlDyk6O+iZZfKC/J+tpmldfl5
34q1/LOzTu6Z60prPJRi88xdzX95BdNiumf8zd94BPNm6qBaEP3D06ep1BldJ2xn400oNpCKb0Jn
nYMoAY0dH+kU6g1tK9RqaBShmQoXTiWYCGVs89PXDcyyoL9J+8aYg51AeJ8PGbj+xbDBz0sPeKW2
1KHZGIZ8QQaWS3SRHRLgyI51OSfpRW/c6ZTqvNiiCCphZzOVprOHfiIZ+5IzkAfz0G5cCFqnNBT/
JfmEr7lRwEAVUMTz0Xe98CugqirypQxb7V/VemGmEL3vyyaooiInRHULKHC+rWvwJhKx83FmD13o
tcTVl4cnU3cgXtI0uPtTIy4ljaQ7ri9GzoeBcXn7N+P/1eGJ42neA2IcQzB+6EimZdE6XXzWWlni
umdh00Ny+iJ8cCEvo3sCPjMLAGozmmYY1R6ESvnnt/m99EdiakvQQSf437p0xKdO0M9SRIZl/zX5
wH4XilthozTMl6BvAN9j+zCygpcyRQeYix6nIIVBI/sfqJHZsDmS57We8vSjmE+VvCm537hKqkOd
yIhqT0eUdjJ/dGA/WyMZrN8E/NRXz7wglBOT+WB55dMuMwAhHGr6deivhZ0R7JgXQLDtKX8rtAhp
QyW6bN2O2YWCBWYIppyzgJ01fkjX2ViaSMB0LIfrIgrbRtvA0cwDYtwZj+mFOZwSCyiyEP2uv1x5
BfeAsA5iTbCBdJVuqbsMCkjWq6UamCXuGUUFepDTMAJVMNpzyWuuuToKefxyW8TEpRuPRDCmj6GW
/cKf75DJYN2bkmg/u7nQoi/1bOwdRL243nFPoXfsRQfJhR10A4F/v6gxGaEumY0LspYs4DCd/SDy
4InP/d2Wq0OdlqXgI2N+nq55w2rlJanFvxqgcEjB2PLu9o5F7foN1l5RC2VUVZuv166F59WVMKJ5
YRd3RKy/+wzLMlaD7uknpxhCkmyedh8e2BK+Ar7wqWAVzgqsmdoAAt8sME7Xlbcc496DtAK2lwO4
62epgkyc6Db//6nQtK9DlpwA1xOHXhqVKLjO7Y5eU3mndtbYYGkyLzlTLOl0OniE1lJa+WtGhx8Q
/KRZ7dJcJDFlNhpFIoTjsHc21o+j/TMgt0DBjN6I8VuFmsEyF8qU3BMyhRGfYMKaA5twUhVOJJW8
Yynqwcuwpl8IA5BsJzGxWtzdqmJ97qY3IT6/763SuI8TJGicBh0w8BocW0suvjO5bvijSThCyiL1
ptIIm6kzfDEs1iIkwTbKUS9j+7p7bDm49UNciaMTnV8XJy0ZqxlW0xVeuhX2OEhLA63uApbaUl4p
icvh0FW+BCunRwYXdJ4tJnKLzIVdKaHzT9hXPivytWqHaqh9t3t+jlXS1P9N4UpYqxlgx37Ngqk7
X1DlbU2R5WMK/HBzZfMgx92k1CexAjxkipNX3afsG/hQcsculeNvuZyuKz6hEvk1JMOLchqK7kxI
3H0tbhvKbBEukfz0pstZaN/OU+IUM3FM/iBk1sJ3oRJ9UdwGauC4d7xvyf46OtKa3ngT11sVTyjb
gzovYkkgFPfT+iN5MAswwG2EOgJWdjSrSnrjRSu26fKkNha8Tks7Ccxu2kCN2NwpN/XDWeh/ZAMB
cGbLO+QM4FdfA18nxLC/sWsuhhfcZ1nALQtQJqchGjBJQ7cpfyoBz/tVWzURwPP5PXjOEfiy76H1
R3wjeDV/iEyPeXHluUv3B0oXG1vrWtHxtJSd1iqPMQYhBw9Ej3Yz0KACDuulU5mECvW0ra/ECQLE
cEswZgMBNOZ/3aclyRQuX2k7Sgk5kd0Zajb1BVQIgeSGOC9izfcsqKuKKoPkKEWI3VUQI0F3IRVJ
/Xsy5gewC9Zx9x7MXj1bxvezZECwIdKGJjPuk6Oyw11qKbBio12+/KQBPZ/4pgsXJPgX6ZEgrqXc
sgTPQO9JJaazFrKj6mVGFoJrnMe/7rvWrTvHmCb7dl6bdmCmEg2jG9of1DwMNY4rbIPv3yTvgqva
aX1uThmEpwHXgudgl8yce0vr/STDifwWsckBzy0GF0L7Yddzf3BMZtcf0Yuwjj/UY0ut/dtAeoy4
7gGo7cHQYjZX98HCFJlJNZp53XBoDxC0n18OZBe0mkyPs8s3agkZkpzDi1Bi/sHRJKe05gnB60/P
nBkzCNc5dcQmOAkj5wP78vMqbaAagoE/YDMcn5SCKjnB0TcGOH4yvUAmf9ivcf1MJSYt64Jjh/rt
ZGpcoWjGivgdkt6hngCLpZXCwnIuYGHahQ/FpM/l7RuTaHR4lBY4CChy7VfKcktm5BFCK5VQzuLK
F2pkiDIzgdocy9mvKUpx2T50hYg8eHYVgc8jeN6FRBQD4oQ6v3wh7pcmMA6FT3Fpz+UR/2YFajMN
HUC+Qe2nO+OZfGK/G1d/s6lSclqEkn+VKNC+g64jChopoNUT+yd1NG9BcgjQb6vDEoBp/SLNHy/J
6TKMh6AYCMJZf8tOftg+KvFrxVUl1IvPNhzC7Cw6PIC4NuqOAG3A3FO/4Zxa9J3t4Ja7T/UyRLNn
+smD3Jlz8FTeGEba3MuI9N/xnjCAIkvTkJFW5c44Qe4lH6u2bbdjRt6L+bkpY0SX1Xx/6cCXm2Gd
Pz4mAwiNaBRBiOQPC9zP4af3TXvMY3jgVi/vY7T/kFUVfJApA52gKj6GzfoyeT52WBxoLpcxxoXu
z5rBgXozu8HN8NFmUBTWsB5u8qzvBhiBO590gJ7/qaSJAB6vA+y8qn8OyTyb6QxDBJMkCfRKuT9M
b2ZiiQtvVIl6JmxY0PyCYkgXCVM2Gz6DxVTrAzF7izoEJswjNKBfAACLKtDlk3Uod8nPBmGT8YrG
ApCbO8UXiWtru+zHxImhQmoshtytbXcoY4qkhE/grILB3ZbLOwwjn+qcIMGMz/fuDqk3uaJh0PeT
eCF8vCnGtURvAPx6CJ5pH/A1jfw8w5YoAcKyGNNOWjUJMTbRSnEt5ArE+/4JFQcWB15bmNhBs+0n
p4sLfo8iMKC1N0hQIMeHyr6bZB7NL1TAiXOlPN1PLiu0/Qcx5A4UGYkAKlKXSDXUUEKmOkWF81hv
iKr8guLDkgpBfRilhpbhi+cppkSoilvlqHRhv9ZgczZHmN8VbU//Fe/iM5Fjj/E/dyeYeyGlhfiH
+tkLNJues6oKV9Lq3g7c4ydC2OsJFWtltZ0lhlTQaFSqDEhnjNNgQXwRm8gl3YUGFlq1mcJiT+CH
qd7PU863/uevj3WM78fd45yDNscwiDGdEAvgXCvvcpRSNLCMpWRobOng91br9+sSa/+DPXnIYQL5
5+np2aLYVQ97sGIT3cjkjqbdXz8hT12o3IZ2ZKv6FgTBcOua6dANom/33YoalxAVQv7iJLm8RF6w
vbvKKVN8xftzRbqbA7BUtIkUcmzuF+qdsbhSgUgKNQxOem4zzoQ432WVALASH7xf3HeF3q8ZWRVs
C1jAvfn5L3zMbbBqFkmhyQCd+lf4N9/zhKiwlLTUAtYKU9n7w7x6236d1qZcg9dCY+r7NT4EaLgL
dUHZNtEdVU4cjAhT9u9X1bQCPT+Cm3yLv5ffYPCFFU89kaVZbeZ7AXhTeIzMPsCffX+Nt6Wali5x
fPPO7W8XP3PR4VKTOgE7/GFIYBVS7F57BMuCApAYSg+yVkPu4v66llMfW7D44UjphyMxoyRH3SC5
wbb5juuZbPrcT2qJzfj+pI9nWGptfdVSVxEtfzt5FZwR2XiXXHPvMEu5ox6SgWbRJHPJ4dPYim/X
qFwXADs6s6yzdNdDUohACqeTlkY7qfPgy9Fgi4vqvO/ZJ2NdZHSWsYYCpcfWEeUgwfZJ7N+dh8TQ
k9wk/v48cT8ZhfugOvTfzMoAnyLrdbxnPYmdRoD67NdjDJMgyt3Kry2bYrOpf4qbp+7CqaWX8NW+
WjLN3+p5IGlDeV2sK0y9htjNk99sHVX0vEkpT0VVQXSGudE4++z7Ti8PK0eMGG5MtlrWqE+6cdw2
IYnW0qJVkzaJpgyD66zSSD8sG+w59Zx1SAZCeiQ+MVNLsSUOx0Qrr7KlXTKcf3sgYOyMc7tgd3/z
V4vF05omCmWeRES0sTvWunFnv8cjc9GRSF34llr2GCWj8UwDPfSawvMzdeCjja8ZU4GGQ1UuHUWT
uCODVbnxSDpuOeFlt/LOJLrW+JHtwDgvBl4Gutuw8B4KvaKK8cRnZhQeTccDwBwFLgVgryelzrIl
F77QbKkfDdW3LjfXl8Hvbzbc2wRCC+SRkb3wJukLPz7jJjPHfdXv7IoicZhDwTI7JblRlCKYSV8J
6j/C08QFAMUshiQkwZYxXHMYj3kB1fA5XjJPpp0O41uIM71IwCJpTq5pZGE5DjMqV2VeGq/VjBjD
RCykSO85N7UODPtLonnLXsYfScZQzWxxFKZt5NUMQ6FrGPQU6TrmDpj/eWNk5cMmrp2vDfmPGbcv
NSByap20+ZYR6Lt1LNcUkvN61f19YVBoxjOnWuENZejo5A94xY5wIptQU/yMe/Wywgup1GAMVx11
X/bASGxPCkKiYEWt+FtfS0xHINrT/Y87q6qm3BtR1PNOHoaCg0n4JX0a7QLDpNN4AmDjE7Q8E14k
gJFKQNIOsu83v7cyPG59LBA29CfhsFPDBLwuiHfQxsvMcY68TN9dvE4spwgC4Ih78Fu0Pm0S3S2+
06ygqCh0br/eNaxlo6LaMQvK8e2cHHVcqQdNMBbwDGw6PsCTJGFqrpk71qGdtiAyo36hioIe9fOn
Nvy28H3rXzANUkD5kcdFdEX4MBNACdHEKzM1lxJ7WLuElqUW74HdhrVegT52toSRVtG/DZYC7oGe
bjjhhveXM+5BAB1F65zkHD/lzg3Luw4ixYuUqCOk7uzSoJtNttOld1iVPygqeQE0s1UYsu0OZ4Xr
E1C+gNvCSsKSaNKXJiPE6pIto/5+PUYjROGTVlPanRGugW2H9xyR5Qe3bWHdoy9CbvzZHtZK1N9x
TvcP4h9wqWYofgbLmZY/U9W07I7D6VBofi0n8dTx+QTOyiMFp2dZZcZxBWKm4xhD/luwhk9f41XG
uPRX00tPGDIMSBcjTMuNzpGrOGnjOCzGHVSUIlckYbg0yi3f8wJix3OT3bc5Z5s3c6yU9V0m4VXn
QVBgSdPGKxtxyqBmMCDQG7hmnvDw5TGY0sO8iXLqoLY7HR89wOqYh65a/9/p4yR5h947WgMXhqr8
xQdGoybD0nYFA5yoOC/4A5h4xiI+PrWl/0nQ8Eh7exWgbVKz8D9+IJYbKVjkG/LRz3l38P+VH9mi
d2X6Oi3l1eTKd8q1OFY+wwnZoxDx2ytNk/oXobBvtSi4P/ggaGVwV3/A/OqBDSQeqah0iTITiFR6
twLFeNHv5zyUh9kLKtu47yWB5x25DlFREP4oj1iNrtrZE5Fobryy08EM5NKhEcjaMg8fdce0fi9E
+yfZ7YR/wB+GwhDcy0ORy/V4AxAci7IUism3dfqZz3PZryUARy84hQp3qzNb3lcAMG6l+1E1oxwq
8DjmBPFnFgZCkig3dznkaJApg1by5o3/VKibTfOoWr1EJ1uNkV1tfPgL+OlPlyNv7mhUHhotdEvG
6QZh3e92kQY+/PFp22hvlWThEf8F04RHULrNJOxDSQPXZ32kDunzMnOQG0b7dZVBEolSUAK3fknk
TkKW10eAxp6nNuthpZcbRnt5js6Ed1S9i5FUE3x+oNOipmDiaYp33/y8zlyBd9kxdLZGgPgLSMJn
L4Kcv10lYFvGz8Lk3zVD0q26GB/7gu8RSr9m4+1rs37Bf3iloU2egppfk484iumf/qrPcH59XExx
6c1RMKJBzW7WTFB/+gM/tuk8pMO8VrYWzHjDH1fe8+datbL73+hfwQ9Oax7qokYujsCrdFr8Gcy/
VrzgDfnxOohniPiDLqyz8UP/TNYcl6djKHHvWV+93jXA1ZABIBYb35pcco9G7ezPst3sRWrPQsoe
lE2mFQq8a9G4Ja1iE4aph2egepKHVswQuhxd8TSGTlfHnkdiBxWvlStILPykt0mcRvZF4hEypGVa
n1wFfttNbW+4bbut+NsbVagNVMY/B0SvZ2YeJtISL0wbmBWDjBOW87fzjTyYRORXGFyUM5uWAjlg
te20ex3ZjwJJwjJi3OmtRW1wG3E6f6npQrtRr4Espxpx5kDw2kPGp4ZhafGhuOWu2H1Au8J/87HM
qa/iZfv8024CaeR8BBuzJ4dGLUbE6ngoUHLy32bXKlFIMJYte3tvlVDdmRpIFI4BFYn5xup2yT0w
EwLQvXDIgZVKZcOaYy0lzeH6m8gE6D0hzZgBpF1+LIuqPr7BmcjIiSiszFPX7YrerP7PY68oaCb1
Euljd4s0hEQh+WPiHHPqjKfagnHFZfg6wl9NTg/UNK1fRaKyHopBlZbuD5r/fwQhiII8TDRLI2lS
QI6yMLlPMtLEmkVuCTljUFP/HRrL5wulYjuwyWQVTzsR1Q62WgiU6wb1LX8WW6Sj724P5/GbezED
Pa61eR01ZcOWvKnMVHyYI4QuB9BPsqjBG3lYSNGHD/6AmxnIZV2a1gzVSAMeX3eaEFWGHAOn7ol4
hgjUs0183NRChOjfL5CbvdKzB6+/ic+hxsz8zggqadhJ+hoPycNvAA3SgEKA9sYpbgx1QXO1sLvV
EFBBZgDrFtAxkajBpk5cdOv6iJgBsktietUZHSZX4OvA7d9a6xlCcHB9w7blEwntRAXP/c9fX0yP
fjqKwH+bAH+k61PnBlOfFyMsXEF32nWrzcu2RKE92NHUu1sMFptvGMo5krXrH3l9TsNUCOIM6oVL
dY+27ddplX9o8L24iPFor+J9p6xGoagUV+n2V2MzB3xWVzO8x+uajFTEa30uImED9yYpe43ASZGE
/c+VPG8mkYjUotBt94W2bH+bj9+bAo2ANpaZHYUcjvtO/IhVoNghxGloO7yhG8qHkpDvDXzxVZ6N
nwiC3okGdqF7naRRs6QMDki4rVeUUqd8iNCL4N8+ht16lP2fNW5DBm+/Edrh6FkhyuD2B393mgdq
a46Z0895N0NYE5f1TgHuG2sinVF/MSHs/r7n7fG+sxOqKlVjkGXRCQffElUMIYTAkpPlDnQin95L
o6yk8c5D1HYarDUyht0ZPjh6B3PGJ9p78RB4mXV1m0TtMSdJSScp1IkicaHIrlYJK0nRAH1V62Ur
a6SeU1DbcpPqq+4zxMaJGPkHIZbMFfyh8zlD1Ib65XdKykWXXx8IbXn6EAt2aP9+D6Cpv4ES3++L
l8+G5yj1GnjfYWRGGMjg3ZcloWJ4iQDUuGoXMd93l37S7dH3tQ82NG1dji5uMCWb6IP2u3Qkjr+U
S0MH1earrYVID3ChzEyKkFV++kUb0TwMsVFd2oCpqA2ihck8LEz5Exk1nNyl2wiOdOYy2FtORig6
YV/eE3frbOaQEaWk9faCx8lCgxD/KLEYfjhY6Rq1blhDhb594aFHq2jqTyFML9JaJlfwg9RA1bMS
EVHOkB+Rl80dp4ZucPkYZm84XGZFYpdwkdpIFbKlpQbW9SFj9bvpyR2uqSKQ1c7Gi2MR8cB+mIux
lur5v+YShhpypeWl/qICSYKeDjSwCY8xIhIlwIBioFH3dOHn69j8dwU2V84VVfJCv9w3n0Yq2YuI
mrEmacnsYW0VW2boKWMkYMnqlRU/uU38Ah0S6y9jkztP4FeXjpjD0mzP4Hm/9MdYUDkiF2MLit5Y
+Ocv9tKyxQgUTZVMUXEc01dbhC69DHC7mkGITuu8+qNX2N2Yw3CqPP+adUBkzY2CQcM5JPXIEluz
5E9qEOjgfDkzqpbdMF+faC3gmuRdxWBSr7+1gNuIyRN96fQ94EI27cWJtKhuJbJV5BcmuT4sdTSj
yVVnqRKLVTAzm7msBJe3GTS1Lm7kqP7HFyLqt/2v74DOPpC/aM0DO/TL5+nxZAJ3Q3R9AJuBWCXs
6eOUw1dNGCua5jo4GAX3N+vRLEywDkmvUzDY+FZWOwb4ptOFCgbM76x44XCeFGr45fFlopfyvfS0
fR02olsYm5dK01vjkW+d8IYuRmEFUpjzhB+fodskcAGfuVK8B2EebIIGknNKyrHum4CY4zyi6gtx
SAMKTrGY86M5cr3iS5c/hAIJCIXwGJxWXi9CoHkjS0fiQy7pnydNRif0UyOBo3qna8MQcnQWzAC3
9uEUmHt++/gUu1R71O+aLT/lhttQIajUjxMO7buWwrrFyfrsoSkPiTWIhn9tf5gDFqCqGPQgAkml
DBvH6h0d9Ko5lnhU3xrtiE9k7/1zXNGQVJWFzuO0XK3nNkV11ZojAKl9u1X2xIvEqSZSCRyTOQ1R
VI0J9mp9OoSZLR1hYKux3Ach06BZ5N6uqxa7DVzwU9Fqs3Nm2WAocUOyE+D5Ht/ztpMIClJM3GP4
ua+815OpAAPBrmg7SMryHFKF0cJ3Z/xiPaHFYRnR4NPguex5Fvm8bdAKs8P3Nq14HLqfBIRvW4/9
GKR59vc7A9ZZIPLJelazkadbPlAZL6zZhv7TLxVXDJdZw85zussmIdzrVbvmNn9BX+mDXYjtZQS+
rHpEDzlqX2ld5xcqakrFQKRkVViZY9YEKyurBRspXdM9GCn2Ka2Pxk8OKgIn7XJ7nKQ3tLFCdOWj
OolL50AuI2rsgnAUCRmCI7GYW+n+2aDGqDH9Gf78I/sC6HlG5umbcJJ6PcTt1G1j8QrDh5ldkWYh
frWG9UCIsItXuf3+NIGQMfAsS0gzboLw/aV4NYibvbGGQItTXHHm+cOLl1yIHET2o6VkhTrwpAOx
N+Wx55YsW45ipaIxiqYh8OnuXkp7BU7qg9JWayFryvcmWF1QsoonZt9EqaXaST4YunY/4VZDQcKj
gu8RJfm5HwRwPJ3v20XrDjsvi7csqFaipcXUxl21kFEjGHBkCCUgNZ9yianh2PQV2Af6RKoW0Xjp
lxTAA1Fr8Gc8HVN83gByuqSIy1+D/QLe/SCJk5ck4UNomQroV0+wrbH5DPqqvPnFi6FYsFOWXJra
4FZAk6z4+Dz8jtnZ8rnatyC40LKlkL6BG5QCrJ27iFddsKwNVqnePpG3LqcgMhIdyK0rayuKY/Pl
eBa7JMSubR/pPiWcmIE0PPzCXuSZFCR92cSDMFoB8ZD3huDLvvNLnXaDx+0gFx0zX+ZFqk2DiOUr
5kNQXpMC6be1wNxe+Qmz0zRUXjc7GjtgKuLR3nNmUch0tL65F1L8SURYgFV3tQSZB5ECPpk0ifcI
z8MiyiETqPrc15iGYIcIRx2ehYf915n8bzMpEr3scRvZPDqOAXJfP2ZwIMVdkwo+nvLb+0H0okmQ
Ps8XsWbQw7eJAKYTWEPDRm05pM2GuiwVL6+Wf7fZ9572inJ8U0dR/tWDqwfrTo/N4y2u3Qulw0cA
BrCyGXhFxOw0JIWbFHJB7ioaMq8qBPuDztTn+4gQJ5Ahyww8HdmcTZqrKheUVG++VqHhNcD0i1dU
d8EMASBhgHCnSl9eHBZBN1qqqapTRAsn2+fKuNR1Bqj2ogDWTR8yRsYQt/5BWCKhxttQSUjZfgY6
mrP1y5ISNGz5ktuiXB2bgDC8Sf1UJlEZQjFJRrfrPeZGgmKFluzLF5sn50Dia9LnVMRoLTuWIjLE
Ui8vWRv6bPy269ueee4NZa41OUy/pk5kvY4ofDOvX66MkblAIAtegcyjPShXwXS4K7NPBhiYGEtl
NrLRZPBj0ZJLdHqlEOB4QqqTzkI7MkoYcsmdqQa5Qjti6vqGTKtfGi9IPqozpy3elDfPRYgLRthU
Zo9kbdTRWWSyh/s5svUkZNY2nx286nmUtCkjXzBrFKg89iCFLd4J3og+orsRy37xQSQy16yPTYDP
Nb6h5xUSmiFpMeewYx6Dy5F+699PO6rEWzC3gRbO3WXqtIts/Q/wa9YnNhrW7nYXTfbsftwrIUSp
aQ9QfEo6rWwkqdPmRwHlDBRXb8NKaNPPwas6KgI4cYJYOdPQ5k/XPleyWAV6TXx1uBHtEgQ5MA/Q
wEAGWpvGwzgc+DgEuKa+NjQv9+1vZl7FZYjtNaeNjkeIcxUFO27d7f9Dp9vodMn98gsN8pu6dd5j
XQxZ6FkD9sXFM0boAgRSPo+oIf7hemZfdjhvZQpn1WkWI1785y+495vsFeOx3RgZLzVmvGyXa4Fc
wRD3XnhaDzppvG33Vj0apdRQegVEY3XqV8XLiqw+E7ejJx3vZpJ/V4ejTTVSrXm1nBZKZMGlCRfy
slWiL7wPjREJYS6vZZCKscisgQ7Ii578AZvxggwSdPn1AfBBUIoBoQCCAs3TnFX3lJyYc6T88Njj
xNzbmDYjByIo/wILCjWjSL2r2JBlWCKkIGBZK/LGYZYKVXfSDWx0rdpQlNptmlxT/N3R+eXf6T0T
QwiTQOhTioSQa0Mog18bLx4qnGWAAlFFYFd7ZgHhpzs6qUAsW6+4CIwCaEzWiHo+VaOQZTQOdghb
kFcB3UTmcUx98gmw4ynzObkvU3WiUByIU8xV/FY2eteq9B0ys5FF2TpWyAw8ab5eDRbtc3giKo51
fwJ3ZPCRFUwFYhC05aQjUGqWDSUuvCm57cL/NHzpH+AIeCTknwKLb1BT2g3BxV++REpUTX+SgHNi
v30o9+7Hc52IDNfiyVtcJKiAmsyFqkjUheoXHHH0dbHOtIZ0juH1TnX83M58zbgOtmBbxVCb7rLf
B3N7jHh8tj9BVJvNOSYu25es25cLBxWpF6o9K2PF+maAjqew499rHWpgIGmQoeohYDo2pzdu5kI0
oXIF3gt69S3YcUUginjnTv4KvDD0b19J3y+y6ReACDBQCz+oiw5xM9WYGTA1Bqd/yEhdR3intILz
SaJWvvJxkfgvLhzRKjx3hHMXFFn1e6o4fNzhwWe7nUqJvKfY5h39dimg74wtT3Xnt+zJdjbaUoSb
GJ5xxhSHfmtFr51Xfbptqoaxs3P+lcVBXprwfFM2U0tjPpzq8vcmBlSoF1avTIkqdcW2z05TkY+Y
X8yXs4kuxXudPlpgDOKpChfsK9X+L0hLJEfVc9mIvYb9y/hp2UwA5+u/72ChKzMhtCF2QW8Fvdnp
yKX6kuFNwH/GqrvVeGdO/UyJYyEeBXoZgGKydeLIpjj+fS9Zxe0GBoIfVvX/IdBC6q8X44Bkg/13
gxYRh+qP3p7d7HL1SK/TwPMD2sWu6HW2Umqc/pMlnNvtwjoJwVImR5FaQfXBiZsM5t0ozAhdcPBy
17kXJrjSluBLrYl56DFUq4QT8nIZboNZjJawo77snb87DSiFebhDyuH0FXhPueI/ODkdzLJd8ZWU
JNBxA9wDNII9UNi5eajxFx5eypbTpDV7rDk83AWKW4uVYPFuePPMfY6Ww5ojtKcFtEO/Pid3z9Ir
RRQwSrZg5gZpv3dlgHT/k4CCCIp+MYd5ZqcAKV/nAHtqKPe/is1MDd727W8JMh+KmNjHc3QYPwv0
UsEBWLEwboNoh3byqnR7ZhjWB9fmBgPPcoo6ldc2KZQB3UGatGavBQHWRY2ANd3FMeNbQYBd8p6/
ESrXrrPrxR0/oIy+K4ssREFKXm9Bv8YqehUhftEAZ3jsz8sVbDxAmmF4HunWUCbU5HcHkZVvDAF1
tOGCSKsnvtzLZhBQ9n5FTXSMXacGGFySXse3nmO+fuJsBpfh+qKQl5JsVTAik/exnUSgkBF/5QAu
47T3MiZd176qrLy/jcG5orniw1NFL1D7yczgijHLTWWGn8wuB14m38CFkC/e8MmCYo5LoZBiTg+J
+e1S8NxTgwWmqxlx8NSa/wUoatrOhAxgKFRPuXk7GJI7pqOBebjzk8Q5Dv+rh/Bs6ixXIndFN/yg
z1ztW2MQlrC5oPYqphvDzJA1hNeLqxmvuO+EYQLjm8ZdA+yGSU0q8VQ8Bpsv92RU1PtkNu7OGh97
ZeGhc/e8+fbPPhhSHIcLKyguf6GPYx8ob8aESS95J9GWUNG/d8PcU6TD17/Zw/kbwNQa4A1tMH6/
xCvOLG1rq3MI6DrNNc9Y34OlvPCICJaZEC76fu18VyWNv1w3TGqGnstolVzeoqIn8Nf5fuReeLke
ODQ9MbiQqI72aBdiPi5HOlqAEZuvTloPvfiCDfsksbs0+CqGYT1Fq5CkxTinTz2SbixML2bFvBO2
16ctpE9X2CzB0cEMduTCKHNXHh6iXSiZj5gNCMoF1NtK9ZdMxET1Ms3Hhj57nHM4cm2yoTJYIhvd
zrH0MO6YlsGCBdaaJYg3GZiuplnHmeGyihdNfn6FJ2b4RHWww9Bfqs3VSNcUvFBQbnIYpDldV9Qf
q5YJaZbyfWYdy9y6kSAdMUB9HNT1rdKSOtCkCjQ/fgu7HOfNP91cdt6YAw2ExUcV+XgEQZ/MxkqK
J7TLWC/gDv53Bb/zHda//4/fqkovdNofH/EYlp1teP/ob552NhyBhNE6sdHtCPDn61xXRJ4aJekV
eI7ZFaqOTeeFvXfgk26V0DYX1idT7rzj8kuvUnbrl7mH1GxpWxKve3U66bjh4zs5n+XVeV3mGe0J
1jvm65TdXfxbAFJPPZ1V3dsKdxW2ox1RIQFm68F3tgRDOgcw76T7OQ+fGCraurJHHo3d/ywsdApn
tDkVv+cVSwI4YWXMli09d1xPrIoEvY7hXi8Flfb1HASMZ0ykb9xWCZUxSLZ/eVemJi/M0JKvfDQA
k2f6rwjdvgRKVrCt8SsY2MffXISSKTPJ3IX769Z0N5LOQBH5hp3KmtffNRKUEJOWlgWEgZHjbP7K
T5gqdZNZtbOAoHXbw2VlTa4/1KoMaQnvZvey+u8bTfhKFS2dSrJ2JsfbERZfCk/yKo0/uOkW6d6i
VwlNU3uvr3rqse5BsBoUgn94MmovFBHoH3M+kPIZGmkic+AiIdaRjEiFdrIK2IWi4B0npErDfS/p
u4IpnM74Nkf0X5SlMjwKCMfszssqfbJSkof39x2eGpEvGXhj1FM6ZeJxyrCc16MAy5AnOlO0ob7S
hQWgUo52+uxw+qz/OG2uvwGmgK9y+TsmhRXoLM3YHKrnLGNqhd8eCtmEPrrFdBLZGsmBinvptij7
VDWTrKGsld45zB7iQn8rCGvqjBSIfOMoUJzej2852SareljbqfxeVISoqsA61mbJ3u7WmSsi1upC
AZCOXqRxRKAa+1doETbwy+50nDrPxhAA4KSMbClrf+ETWXb3S2OwyYUKSunI1AkoCnvPozWIGjfZ
txKGspthzhQ9JibiS3pKo8jK0L7+NFv29oaFq5Hf2MX8YgStH9lNsNOIKyeXnCLmrzJWuU2Cr8kw
ZuWtORBCroQ5P82DKjwS7AJLRbPoaRuwqk0eBVJQv4rZrfqSBo4rL4O+s3h+El87PBKFM+K3ps4+
LthJOdzcj8d+64KmXfo1djOKIcvKIu5QxPPnEuoV5tnjIwupzlgoXz3fLjUjRSdC4510toVDItty
U3BHRrTZe3sarpGw+0BsHLAv46QSNDiz1tcHLpU1mjgVA1a6IwOJeTrRN3VGbvCsIfDboGK4uiDI
oSP51Vdree5nRx3lbfH7qclluySDUw8/9Tja/R/0R830Qd+Iali1LwsOievC7cniSsqCcsYg/Lci
9x2jJCOU7OuxVqOXd+30XuRo3lqYxc0Zu17fEz66vHDnwnRH0KoORQuUreJx2EozB2QwZ99pBkoz
JtSJLrdBzloAObgpQce2GOOo6OeuO1GDRQWWjKxKiPyo/Li/wh9Uja+pCSSyFQw5/opgL154vQQy
st1S9huU2kTx5zSmhsLaTHiJz2iBzD7xYD195he50187DPaH3g2QpmSKw0LhLl4eTLXfwP4Vfzxh
XhNzL0jKaKoh2mSj2nFF6sOMlaf0G34YfmMNokObFzhFAZSq8LcaqDXvfPYKZfE5IpPjD6U7WKw1
uXvi1gytL51iBbo9/w37mucpxhcd9dN6lvZO1DTe2BzGKFV7/ZNSskSX02XgVCrgwDce8qtpWmc/
KrHDo+NybNu6+ACOaEf8oEKSAByZ9pSjgil/UaGtYMrCRpciPDZ0PXPqQCudAP79ag7dSxMFaQQT
kbKaQDlWMOsqYg1Qf103TA/JRXzGoYB+tInQ2I0OgCZtydnzqJqPomWtDiol1gVyANykOwWnUsup
H0wFBLa0DvA7pIbJSlNrfdl/J/2Uzt4zTrKfyOLcNmqIzEU78UOlm+CuD9bUcs/Cg8Td8IBOw32i
kY77/pxUtIGgvowDTuHvNMsLPINLIZRS07NZAnVpn/EdyVO0ekUtC9ctuqOCnXP8E8FVh58lQMdE
uD+htiy9IlIafx/TP9CysBCZtlVqIKl5rNslSn0X50cgc1VjjaT0zCex9zHNJkYZ76LrlNJ/Lw5I
uFE/sMz3twRWM6I4S1OdazGoZmCf1VwJjU0R/vAm6x0j7fDcOnC+Qg5LyFxIsbOsY8nt8ZnqACm5
57TicrxfKUpRYVici6vraN6ooRpOazUlkwIkLbwhrKbZDAz53mLdLcnrFwO1Dbh0VUOEfC0kJsO9
J1yQoQbkVzP7jdUd4F0NbYuObXSTp+VLy53urvdI6yQgWwDyZIi3OXAWoXh7f4Xed5SnTXV51Bjx
qiCHr0s32rY7UfJQN4fGPAajvw7YMjWoP4K7uAjN8qJVxuBHn50spdbo8XdA0gLN72jPy0RCyC4k
szUnMmOX2Y69TIOsIUp13xGg1J8qWgi8HWFg048H/qitLoqBhRALDYnGDehmE8mMNm5p0oF7Mf9K
DOYq1KFA9S8fM0aO7ynumYYRrNinHdVAdMqE+urrWVaYKES9twg6Gebfc/+2gMx2zavtbfMFFNAl
aYle7Mzq3x7m+R9jUmh330uMSv/f3nHllfzpE8vQqv1cLS4IDTNqUs2Fo3Y3Ap9x2SaXwKKf7iL1
5veHajbVh5ONgrZAPZtBgflMrK3UFEpgxqbmwJ82+4hawsq3zceVMrR3Pf5QVId+NkNLDEnMF20x
FjGy9I//4eO6Qwqki2x+CcvMXfuNpVIzwa01JVB4YsbwebFFLS5HSdeNs7jhyLOETu7Imywb9C8n
AYkZAmJRa4QZbOMJbWAJuj5PFz8DnmQqATaLR0UszlnSIFKzj+L9pGF7Vsz5f639h6eQJAVkpkHT
BaPQ08kd/s4tfXpDkGvVTuDAJQCz7fFCaGH/Otlayc+GIg5MI/05TUBDAEL4UQSNIapCLvtfBMKl
a3j4WwpAKQ8+rF+jlKuUihbeVQ6rf5p3DXxNhLjIIGv1CII7EUSEdlnVQCiMdEcdoBgXUnZ5FZH+
MJA4TyzvA+6wfqjzLBiLLcQvkO59qxuzexVX52OwDX9QTDGpoRc8xrJ9IufnZG8PbirVFAEY2tZT
cyqfNz053BRnGEKvJY+ViTbh931RRA+Q2mlwGvQkWSdCTaAfjoHQGJN0BMT4bKoawId0jNNHfTu5
1HqEAcSq0L4WE88voWiJvLOY1GgIOJoQYupJWtOmXWtFz57bKjiksSxvKuLDb43Nf7QScxkfCcaa
H7yWOKIYESKf39wz8bznXilh4YxLJmGvbjUsL2bLA5t5Iw7GcmUDFWPl7UENSLsUwAP05J3fu7JI
r8uyUFJKKm6Hm55sIUyqvBbfvM7a4bktI72YwPwhtsMWd2xdrxUpIC0jZk5+cpUDt2O/gBwgbIqC
+jjf+TVazYEe67gr8N3ZE8bRd5mPFizjlvcJNy+AvTGIjPjrKJqd3tQp+qk/7svAeAehIgjqs44J
1ziWD+/ZUkZg1vCI1WAiWQLyu1c7Qo2ubE8O4WwdHumu3Wbv0f16O6WTAq/gBfCxX1xDhghHATgk
QiW1/YTQNg6di5eLp4RcE4maxIK7Mlvo7ur8QrbOAzm7CZNx1TRij4wVxBgz+BPTe/iYbda2gfCp
U5TkKCQW98La2M1eXRyp4MAjLgS/mHgFoU+HqyPLljqt0k8TJla/ltebSSHLHDeqHJL6q4qXlcgj
/cZdRbifIR3gImyswGsCA1TenumLVYA38I4y/IubMmADvQ5TORJ6DJ4zQ9spipMFd8S9IuQFCFaF
1QkpRIdHRxFeVT13sbhI6iRmKSyuRhdY80NJu525vGd7eCmKcha7L6mLGR4uCWFES+YkHIyt/9Q3
zJoJUY/KQ/3K7iAS6aBRgMCnkvof098tuwV8ri/ceIo8j+WqAO0fiu8nNtpAxkB5b89cICbrPpw/
79w7YoHVPEW8n1XbZbIaexpYFk/7h9B3LbRwM9fzfXvutd0szlN6AyBVWBoWr7YP0LtIQf2ipP60
adlgLytR4FOMPOdqkqCSNqposKATZ/EnbO+WtoGbJjvWK+uM8I54JOp/PrD46Ncl4ETJD2eH+fME
MnNBcpcWGQCMnLShElKpcFDosOlC88Ngz49e88ntedFgMphGZGoSpiCyRCqdG7kCQFRJ67SpVfpS
uliXh1/NCJKRHtz0wW4nzQnqEDW1zF8XVKukHSDQcrSiHHXwrJuhYYGv0KotF28aggGLr6so2Uts
vitDtbt4W9JYvrddWuqce3YU5wuI4ucrkjA/b8FB7Npeg+2XEXMtB+xAVG7Te1d1zR2DHX2IXcx9
tLi057F+TTUFgGO91c1VBVVUulgh3iGFKDLSu0sN+LYt+bA6fNlBSv+acr62nqDSD3SiXAl2qPoC
sgaRmzSv56QcaK383Cpe9Q7Bk2Wg4R4aF33b5RSS1YHMr6wRAQ3FQjlgcsi4J5PnmNEKtor0ZWZ+
HAYSZIxTo7RYZNR65TP22nHacFCkuD07pMpc6WxOq7FhOT9fo/kxYl5Kc6iCWsPoTLWZdUIJdFPv
kZFAWjJsk25MH1Q8m/ZOxpBHPvbGkvNkFFd04VMrl43ZIW/F7/M7HKUheM/Yg8Dt0OZDJoz5RXW7
VXQIEwRJ/dQ0B++d4l4h31xsIn6UTEKGLRL6nhbUEWQilP3XZnJl5Xfr/gbuevmZ0E7eEK9To0gm
4Ymo3p/1BrDf3oyTjHoZFpSWSKzjgV+qRjI20IXjC1dXPBGvpHMnmDd19W6CZhOY44KpRRhRTdRB
8S1TzAnmm5jsDI9r+IFLJJxZxZVDmI+F2VaKqnAw7+3TdEAFHFPIJRyRMOvIOebYMHwiVMy4XOvy
AnRoFpRQRlILHsQxT+t+3JV/pmZm9ymTwqTEb5aDp15OOSV5kd+09oYtMiKVB1x1aSwin+7Ku6nA
ng9AxrhyMFviU8PnMxdwS8l+BoIjFoKWJjGI7zYVREdEMbtbfvF/Q9JSqSlsWuoFaP2pC6VnfkP0
sIxwvNybsguhvMS/tYO1zq4ITtU23M2O0zG4OKGXWfVJ+fibDYKZFBtjOQoNao+dAvXB8I0ENNe5
OgF1yR/ZZnRwlDeE0Y9gs5KSi2oZEjm0u/jdUDJIFK5gdx37JT4Fwy4i3cmau22GoRthosowjeGL
5GG2VwMWf3sQXjOj06jmaUtM9iiMI6BRjyveUtkyfvCb+Z38aGKh3ANdHqcEnLYireJ7YHF2or+m
erTxvjFnQhuLOsBRdbQH3fQRVjm98KQdyfiJ5u6su8U5Vr9DiZMNK/IEE1mIFgavTgrYU57/VLe0
+eQtBNeyiPcytBzxEpP3/AdHSCXSqo4J/bDzU/7cYb8R0JNiBVPPz7AgLuL7OzNKPpLU5OQSKs3i
wAOK3DnMPmSbsjfu0lHy1V9VHHnBzbEOjOysn2g7kmfM2KflHujMX5PDvECcreOF/9onwDZA64Ef
piVagHhURzEKN4wsWXdv7TK9TF/vWSd4TG+X1UaBVPPIODxMnFVr3L9E9V3dU5nTbIh9lgApURvf
WjIyUXORfu5h8HnHYQqYZMcSnylGh/+mJuwIRC2Nl6XmU39tds1lGcWS3m7jvBdZxOnfq8LJ4MG+
QtpyhPV7mnTNj25UZZtkRJbjyPbsBOWY5Los4aHztRJZFO+y+n65q+I2hq6dKzU9Jw5a0fnQpSMB
XjVggTOpQZ6qpj183GIOjozkt33sljRMn1rbS70GnxQx6IqIa6OOSBl580goPNZv4ddZwgbCn87B
Iufvj1FC8z+cBFR8flVaRS38S+gQw7VNGGZ9yhJ2Nzj1xspgDDOQo6Cb90ICVuFb1ieHSNvmNQaz
cGbIeqZkuacftd7WLnp4plsOQPZfTYlCR5gC4mlmx5Nkk23BxtUFzSx7ZQ5s4d4RNTRjjA1p/Ppp
oPZXIcy3u9zuilq1EY14m0EDxW/B8bBJPKeJU/1I9kFkqHsgYm/Sp7GIfyRgOzt+zaBun5DBdyhl
9t9n6umQMI6kcWhufkFxcAMx+W61RkOMk/HFD75z5AXT22qHxxDmhT9QEkEmYpkAz+eMPrHh+hUN
LXYOSt9e0bbM8jF0oX/x8ZSf89W5kuSfk5u2lFxMrbmFdakh9TSOO1Bbas60ATp62n9rAOJm08Ey
LDvLsVLLFK/W1CYxCbM2Vlxpz5cY8SwXBs0FFFs+FPnNi/xqG3ZINDrTLoZVcHLroIxQyZTGPCA6
/i5pHWKhOIinlnICvqpJXkF6tPGY2mH0L9H53g4YwKT4kamJmbt+wjdJvH0JBn0oYqcT5k15UZdf
Udi1pDQXYmgGmIDhnyla7YoQx/r7arrIpCuhUIwlaahoDeCDTy/VrNy1bJ2tyUU39jObbCE2KixH
QhIn3D0hv/Zsw8JvIlguOxOeL8BvjpJOnC6zEnP5FVEYoJxUQECs+UObBKQJPX6MpexgGtMdhEyM
iDzLQWzkg1hjsh+F2XqBswBOALTDWej5DKplxMacfP0FqSeLASF3nNe3otfuvdYxKhxmbxeuJPuy
VAy1vYKV0a4eOxQXSiXjDiCho6heovtqCwDxuVC646L5PALPBtRAoeJp+Aw/GZRYHxCMqftntav5
2y2vaTJijkp3C3lqsimsV6CTA8adO9EO0xDrgmrYL8OUSJAz1HWtq/PdkACjwIMCGVBsCklHBwbM
/zlcAfFPz1IO/m2vK+SY4t4vp/xB3vH23RVuMPBq0KUJBaKKEjENT6AzZKzzDRQmhUeKtx7OPkK3
FR91smwBs8M8iHwiDsw7CV0F+6QbAvJhxRACuGSz6KMb9gQt9JW/sUOE/zmFn59vVxJhCf/+b0H4
p0LYSu0M050Y3phRq8fQma32RdxkTBvNWYUwAP7smtHBN2/mAZqciYGh9AsxGQ2wzXzVVfbsNlu2
+92A49M4aXLzj7fPCd7XWUksrf4oKeA0YkZCXsa0F7g6xDIe1xpK252QrcZfeHWeTwU6NLNk/GB5
/wHPQkT0pPmo+nGGyQQHxpxkVV0hDuQZ54PQEXPbGlhzOzfz6og7m4ZBKFNJYo68vpnrJciF21je
XzDpX1GeLV5rKFw7kV0qa9Vn/lkjuHAoEvwUQuf0bTmRe9723zzlrWTKVq2vdirpbgdkTMYmUAYh
hqefJ8oMxlYyuo+UfyyYOaHckSZepbdTEar5El12ggnO7ArK+LOSt0Ye5St2qYMn3gnnqO9jOoGO
JdkgbNyIb0/Q027S+O7pM6ecr0mqOqgQ604ykEnQHtOcj8HRSwvdGovlzk2bD+QZD/NHeyOQdre6
ahiWW5Nbp4puSQ0ZGJjYd4U32peFDZjIqyarzO4GspvUZKNwLkjo7igCBBxO7IuJp8ZlE60vurZ0
gF80xIkd1spAIVKVH0dr5K28DhYm0CBw6iOZLhuTUoUhRtU2uyoQF2F8GS/1avF7kjplAjHs67Qt
3bi5VN9AKg4pXeXUvXLfQhQtGhKQ3o25xk6SnToEC8p/ZPoCrAX/6BJqWgy2NlVDeW9TLCcVn2zn
HeXp4RazGOMzfUNA0Vl6KOA4DP+Kjoeyd6MLTK7VOHj0ArOZg9vo9LASxbZE4kdNhXOTrBcwQSuv
OuWqb4FDs939ZUp6qVpSbD74z5WIcb01N3hG6QL4STTwrrlBekVpct6Jtp7lZ95ZvyOg7LCnMJrZ
tMGe4EPPmXmFhLUhCguN2bkmTxooo5myVE+Nqn3ePn7W9BYHrmtzcVR3QSKVTxnNMLEZbry+ySEs
WYAQbM8gVcbanC7dnAl+hZaiKBoDVbGfJehZmRYqrvlSrzLzbiVqNZnp2fpfkqGGBxlc3NpU1yzM
OuRqmudw+AVVXpRVk0yTBzxQH8Ei0iqTdYUIZjmEbqa6oJT2tjmGg/8es+3TiJYMPbyvxJKxrI7F
YScU07Y4g6tKFdAtChBKSl9PsrdjHz+8GEH9P8CoqUoT9619l/ggIpq2rDs1XnU8w8twnkusVvkI
vC98RRpChFHZgjvcDw8tCfu6N0dsY1mx1CtvuiXAiD6HVxrhD9spQt6J5tmpJZFR7jXAxIPRkB31
omno63CDpPZcN/CXY8lkyIWmNWdVHkhrB6Q2Ma3kJ328zlM9obTRidPl1I3CFGmXhtEEqg6TFpvR
PZpMWCQGi3uL31+DqSB6rJG+R1IXtFvV9Q5gzD5AWQtwRFkWjB7kT4ZguMxDTW4QAcaXvDSoAd3x
lm1sxMNS9eDc0VMNVVmsD0MdTSXjz9AtaV1x6pEdz6orTQjorfw8yTOeLtgX4YVyfPPHIAQTGM2X
BxQOv2CdvP1uvW+KFEOuCnMLScBBbeBUvfldZML1Kik3Rk1aipPqv0cBfYgiyvFuzNCFs87/piK7
MGQw8092dFLCn/CpTM7LQGMQgjElgqpeZmxEYi2Jo/CHGUKPuQAxsGwv1MIzXe/dDujPvFyjIHxL
itta1shAulMRD1rwZ6iwujhKxr28sgPXrHCMMm75gUpBVSti2SPEGGZULt0c9qmjbe7elC7zeeEf
YGLj1yQyN3gcOfuClqgSspTHjDLWyC4W6dwAH0SBs/LSnIt6YdgyA6Hm7mc+tQEtWCYkWqR0WfKG
w/SwNj+pE8PG0LNvUXgCf8irl7xnVD4lfBoCzURLEoECL5kSahzBQaRnp8U3lKtvIA6jbwZT2frX
z3NQ3aV9Yuux++puniI3vtG/bJXOJjOsGU1zy3Rc0WWJTPBU2/ibobkos95mGleajOj5ftb3c8Qi
7x6xn7I2gMm4vL5zjezYf8hjQjmQtU4Zgg8tTMdV9vE7KCXoWFrCS1EfiX3ZcEue++4sDP+Lne8D
wBqzwAIfFTY15abhoxLp8WiOTHjvYmvoiYyd1/a7eU5rYAhFvaeZKkADRurcN2ocs8QwgzDT33AZ
izUlhaKzTRPMaBlscH97+LpMQ6m80haVi+znUUebi4AnfS/Ff7P2lLH8fm4uFlb+nN/FoYlAyycP
+T7IlAcXPWF8nesgTHlSX0Pol+kAKmPdce1XFB+0P2b3TIasnEgJ1yzfA+m2ntlCxhCkMdB4cCgE
cxoThCZX4MsVn8FVxeCTEEKSWVJoJCIa8wvoC3Ym9E7gwJmZUfRSN9NhxHZNnTu4RWJHL44jEJnT
miQitBzipnmkwcIUqLkhhYX3No6FtrGRmNzMCzcwQcNz9HGDpqWBktO/J0Q406+5wS6rm0bEjx9P
D2Cwvl0FCMnrC8Bbl3CehKrtlpSkIiuXtPg4CDKN8fi+EXkoGFg8w37oQRQACiKecO9tubBSq4T/
fWsnq171TiXHDs3zC5vb+nMstKVDNJ+w61bn4Hb+OxF67jQJZwuJZjXwZ1kw4jdUaUsq0by1elRv
KBiEuURB29k4kaLG6DmJ43Swlu5ps+3ecrGnZJ8RETOIifoHVJHQkcF69b1Wsr+c7nLO+BsQ1e4Z
S5xjkRUou5n+/Ql7WlFEKj/ka5i/Xoznc+BCBXaPftcDd+yzIcIMOB7msPVE7BHkfp6RUrGITE1p
TxCqvjdhJ4gxek3LkdgrUUNCdsse6ZNCFJSRSIzi6Cvnio7G2EiJG/nbNCMn4QGO/701Pmchq1XL
bp5wFekYQrgxTVIurwSSvMzDHHMpGW0sLuClA1pRcFrHbof5BcOSAN4cRHhpHIwW3Qa7qZE6rnmc
UuYJMvPgmS2tZN4qDaUPVU96UKMmadxHZi0N9sh9NhDP4luiexJ4MkVAhvS8CXs1OJ/yG5nWmNBK
8YpbyBA+pf+VLIvjuC50bDBSEDjQ5eX/i3Ujwlf7l9SK3kQYQaKoHA2CC/ntr6gQs1vhlxKJPuBS
+jhNIO/DvvO+2SatwROk+L5lqAjuxWyTyKtxqYywGU4oJahmYyIZkfIh3/eC3rqYB1NZsvB2Hbx+
FXcZn6GWsSsg+QY7Fnq91IovnYYVUSTYnyKWcBa9rIoImOH9cqJONo+Dt4RsvUjIL5X6rNkenpzy
ZGNH9R4MHcvUFGpttROarmsWv44YqAzJW9hG5qAHzPUipeQz7xrdaylhFxEW+Z6GGK1T/0lZTRTy
O8s9b3phVjoojzyEw4XlUN7/42uJTLQpG1HPHWbxdw9Hxg16unOpqGuE7+B5cz0VPYaTrBpW65DT
XBT24x1QXxyaLV716Lh+HQoAFsSueBWhn0aIKoj2KDKYz96H2kG0Ff36SDPqaZGQNKLj2rTwHhWa
gVXO5h+15D8LDxC2qRzW1ANuzkrJQ/OgxWiXr/N+EMLkWIEDQwfXVlpCszxZ1KnQdq7lSafw05je
/cU258Ak5NOrDHwlZzuhnPqU+FPoo5YHNrgq4YnKg8A7+FWioZTqE2wpDQ36YjG7OBMdvqFxoxhW
fRN1B9k8PT84ujAasA5AdtDZ5St8/cSykug6LS8CM9X2MW6n1Px8hn0MKU5ycsRe4X8eh/VW7Vg5
NrtZBdahzfqLG+vlWxKm7nk97A7KQnVEejrK9mKl0dVm+e6j5oaXUcpbsmdC1gSNO1wYZeHKoqoi
rXNA7Y6DH2cu2nRgbIiZzZ/v9cjzNxmgQ3ZR20hMKFZdi4M+Q3F/84IGe/nDtlc/ZP12EYgCUr/6
B8ddFQX6SuW608mQftSd0bxeQQSKvWCPxoDgMgfLv5EbHTdlcbhDuGsITLeeo3xrFBMCJpy2bLC3
hiL5BA90aZfojkI4nM2N70LkV7X+lpIVEJLJ7rNBHKbh7lyHxIqDIIP1jKXoP7J/Z1npdUXfZZ1S
iwJOhshanA1fu9DcMew+ZhaKus7ec6eEfoeQ0yah1IcAxvE8VTOpFf1A5vLqj7cD1SNpSgCKv35e
GpkIO3ANfWGzBa9JthyixrAYDhPh1Et6+mBlY4H2wk1HysjwVn3v9Ym6l0EeW3VyPtLjmV2UJCGn
+ZwRJcvUZ/X9mENc45+LFg6aCesTRQm7UVtPzEgjdUgbonADeqnYMx9Q5Sb259MvmCnkPTFZQGah
Dl9beQ8chXw21Cyb/PoSDhSPVYo4luAHhxBCjMSQtrBWpWW7246HZRy5k2jrIUOUEybN2B+3FO/r
4CSr4aDV4LACQuyeN9NBl36ssqVvyaRoMGNpsOGPVjChYw9FBDm3/3fmXQBfIODRNTYvF4JJRrFb
TL4KPZu8haW9n/4mTPwrCsj81EeJy3cLV7hMKBFtF5jmWrjZmDVLycOg8ra1zf1Bg+V75V/1T814
TtimuTZRPzKmHVvaAsmWFRu7Xtl/cpKJ8YD8mDp0JGEVnglI/9PtFnsuG/1BO9Wqy8Ypg5p4h5A1
clUhdv1HpIOS5CaKEtHzmVzUnimdSF3nKPyO0exp7qzIvgrFBsrrG4NCZGVFl9a8bp7LpG3elgtd
uT3LoaqbdBlS8Fr6rveYsrgJvglnJU3HMYu9P0TnA2PmydgkfK2CXtmdp7jh5DeCcXKXcSeQuvgA
SdeddJfzYZh8XmwQBEBY0ht7dT3S3rIrzU/0B7szKhXTxql4MiU6ulC6LODoYQMWJ+UfXEx6wP64
ZcXWqeNEq19gAcm+UgeqWuktmys4icTokW2tFunXxXaj/dw+D5T6AA67AMS8/m1kP78D05uZDZ8O
xF845++onh0FtrXIHKI/zk+g+awoVdebn/z8lzxqY+kcmOZMa+wHhVtss9K/x00d4zW95xzGAUzB
9bQGtFf21u/Gkq9/Iqv1umIdvgs5SjAbgnMCyv9s5iyQGRIa9Uob5wXH2q4K90rYeS590YcEeb+m
4HMN/gcwSdZ0tElJgGe6FVDn8Fao87c5nhuDY8X1Iifj9vITIiaRWkwv82GFVIRi14Gaf8FOB+iL
6jlp/to6LnrPrF7IyBCByxyJ/vG4F4AK2QSnIQLMJNmALZH++xXS/tB7rsDDZuHbYNxVMgzPLZj5
V3LhHcESrsMMUW81bVFP6wCLUqeTei23FUq4VRqfVN/bgtvS0aj+EHTLwI6Y8CXVtIZDR5KoXogU
mFh9N1itKVzDbIht52Up1K4gFJo2On5Js+BflIp25g8JAEledUqDFfcqdPZT6u9mU/QCGn/L2EDK
820dkSWqS1euKwiQXVP6mLdSmYZV3chtPCrj3R/8k83+DLN00gQltGz7W58BNCwJvTnvNcLCd6H2
ehbV0liKVBoTpyrrCvEumk2A0IZzB6WZsBDiK5EnlKIESII0WYl44TZvH30DEFtilMonQkJ3n3NC
ysTx/52EOcRY8TNQEkTwM7bgccfeDkJ9JWe4Go1VXbD53MWHD8lWN83vJjBKX6aWtugrE7O9t04i
kfdfVMB9e8doNmveC3grZ+swyGyoE3TgBFDHePb88yyTZ6S1KfVcg74zLvpUhIPnpZr1jlrSiTND
uY7T9Ajl57DhEGSch5suYPOtVtr7yggZ5eN9pY+UlpCmpa6xiI+Vz7t3J6xxwscnmAR7UTnd7v2W
l6tQCt+vxnADscdW76Zaq+uzPvJxcjCXZVI/hbyxVFXl2E2EsTlgHGzdh00FTMwoCaeIV8pV5UJR
3sqWhHYfy7x4ETGrqu9hWvrp4VwRi0wsTNwiFWaZAJWN029fH37mOy6gqabazduObrfuiFrdNkEi
RvfRO+jBpaFahEOdHKAVN0r3IAxaLtS0m1i40cMwa5ek9alOz5E++dl4zeRYinvdGx+ahr+oHDSc
+6/Anyx9WGmXdqt6rctr2Hi8GNbNeUYvdCqqlSFQmjrfC3ogAwOKFZr1jIiecW+2YmUm5qVk3Nxq
7+A4insBJ0BU8+1OyHIS8aUpGLUUym20K/0DVrfiLIxrctZ78tvnCF3wkU+7n8a4xFmRHYlndW/o
8d7NAoonBF3yk/YmDOdIiumiDIS9Sr72Suri+KLqhLg4lR7Vd2nGhvpd0T1rOoUzR9Gc82y5hLj4
NNhHFQbS3nPzxQjD3OZSk1fuN++fc5b9Gtck64B30sXQ9z5Tu/eg3xnpL+hZwH6gSNfp5vgBTAIN
/sZRraG+n5uKdC99EO9IGWu9M2oZXf/1Fr22/1LnPwnDeJ7+/sgGUYQjPxWvKTyuCvjmmQL90KLH
1oSRltWKRYFYC1W8wpij7zf05cI7zsF/K3+2HHE/KKOI5OtLfZxKSfDROANhjSNvHOionp4NVcBo
nAVFoyywzwW9uhYrnHAyUPEDImCYKzNvMHSxk62IdJHubCZAXGQBr/GO6eXlqTcPDCLJCRCztgGx
fXj/BkisBd/pbw+bYeEuHGF+eQF9sCukEbCnHQskr+h6v4GFrx8V/cGimTIpxaZGl5ipGp+abM9l
NWs6oCC69p6MZOSQy671dBL1wyzbo8yTfcQu3pjJ73vIU/OR+nyvgk8Px8qriLGGXpeuF4uv4WQb
uzRLoW5HAlf7jLQ7VTUg4irtyf0jkNUCMqAT9BDCHcmFOvRpsO4vxIeEXkYE9SVnoZmu4RJrtutZ
hE8wv+cbktrdrv5gDMM3hBskwsCdfs+5J00GH4609Hy/Skc03m6BQIrIb5CJq1ECIjahto8/EG++
AOqmmzbO0AZY70zPLNsSElK8oWlvucM/g0+wAijyFKPDyyWSyzIYvHYiJM4deFnC+5wEH/DVidui
P22rdDBbxyVUSg4HHg5EUEw8THfcITxJDP8RFJF3eKAustC/UXM2UM+nSevtq0G6nXm29NLAK0XY
MpgmVEH7LVSWOB1tKsJUUSY9xcXxxqT0BCkNP2bZ2mGU28Ct8uwFvFmxA9Djrx8n4q9kNODYHJoQ
nksZ005L8O596KaWm10L1Cp8NaM7KOMmx5t/+N0lNe3LgLE01M/qLf4i5x7hB+uu4arX+TYszEe1
J5R0UOI7fOYrNYdwxVAad1hgQL4vW1mD2xjHmGgroCY1XuysZu5k3mJjhQl8IS408lA4heYpa7JG
xwmNGjv2ByMu4LSmwjtDT3kTscWuQ0FKvOib8mLSzobFXlUbS9xAYGZarWzcEPEyMojXunqn/9+y
gl6moqNTgCGtW5RNsHmuf64q0OrPslhnkVgG+Rz2xGyX0LlMIKxRC6AS2tb5QGToTPWiL/rT4+Tz
rtnH2BlR24RUZIM88hpJ4scpladFaabYJss3ybls1lyLEVSUxZaJsPsiCS5Ssc3akyLUyyNqv6dd
eeLDuvbRPglgqIKJQUrSaGTAdcezQemOPYxiA0xPRaYU12eXb9RUO4YFxII4LMgUeazkKCQc5GiJ
Awt2Rd6N+J1md5I78Xk5Y+4uy/z+iF3yZPbyD/rd5Uq9hcs+Rs+sdkmJY1himFoctxdI4Ev+T8Q7
njK2QPyS9hlR2UMXCYuXgQDZhXUollCEp7oyXQ0MxFhvBH2Nq4e57DA3nLP6mAR8YNQmfLYydlgX
sxraVODhHWtktAbJ5UDNHloNVNy3fG3NnfMOQafMlbCK6aUUiE/Td1fM2nOjxwt0JAR33kCfx0aI
PkzgftIdN3jMB0QKnZ7l9ee73yPQV6vh16MY+Axtxh8N4S9PJeeqc4F2rNPd3rmS+R24H3s5ZBCT
Pq+s+gdIzQlz9ViNxbcTagTIkQKkvUnLGaRRzmFqFRQSUVwuxdfEKRg7l7aG0rjp5wnMKS48kVsv
kdvURPcbsy/k8U7mlVIXLml7kYAvOjJ8wlCtG14I8PJYOEiqobENT+veCYd+HcSSekZKmtehtr8r
VyO3YP6qWH/PXo9H8jIyfX7VfkBN/UGPE6puQaHl/phXMkiCVGLF4O/cOktDYttdDQnTrLV9pOTd
04qNQXEVMIQZk+bBUu2c1nYXMpfo1SRTrEMR8nFKyqL6gMzKvlnL6GobB+rZrlIMGLKToHBfQqCC
sr32W5Jj8f5KBYIbzww5tLXAAR/ODBXYNAcw6DJi0oB84ufE1PWc9UsPWV8JpL2NvlFzXe5fc4ub
ji4WDOMjHUPAjqCLH1xdkQNUuUxJajH3H5q93nWAz9sJpw5qJ4QcAE3Wch5yzoDzOTAk8/OoulGq
qA6fImMddSlh1QQTtD7AsU+6UAzZx/NafmAIUpN4xDC6NhPbJFB8ESeqUqoF92XP6hUFMBl6J4r+
fQsYz+qFvdf5x+w5+xOfP3pnI4WrpWh32OLO3hrlL8tV4Sq1e1+QIbHjVhA7Q3p660WYwkZPwUw+
PvxKb4+rlIjxGWMIjF7tDgB5/QIsszPgCrycUo7w8BmSfKenrXVrIiA9DoJSl9HFyzGkgtt9rgrW
FRFvoqw/6kLrUx7b1L+PM+rmGy43OkG3f3GRJXapxZgQuVHMAbKiLV3fkuCy2omZYRaqCcym1fk5
jaHgFDV+dfxBP4rFlNwp/pqjyZ+sh5uuwG4cnibtSO/9FwFbK3EBfzqPv3LADL3yWqZvNL2CaMAy
YF9AXHSU49JhdptlMInhVbVlEWOodch4VvxyOkXy5SojB1uBXY79XNacvpxFKr9pJh/b6wUoxTby
IU+iwLYED6n73kehFSqsvvZBt9lza0PGsfNd9zUqXENkx39sIh0HAjQ6K6hO/0wa8HIJ4OyecBjS
oKHdedLFiyCGtQweXmH3wacWodwhaaGlUY1fwGQF1lY22RVnD/qKPGYuUPBmabmmHovpwM3fagP0
KxeMcApo2o+mR77gsuQKKIpQC2zNQgmGfGjOfeW+tJ7PsxOfjmX31rEeIJSyG4dX3hLwpAiXPGDy
tisgRH7LOPoQ2yIVrJclKTkSCQ00PYZDOUKsCcN1j/msNgDTfprDNUG3ca5oMGdee+x2yMwEDEt4
HRiNQ5W9neBOEkWEJ3t3ASl9kF9Wsz/TL/21OWp53xYpybYyL4I1v8FHtb/lm51wr+GH3elTfHSJ
MGJUz0vJsoTm91KjmF9WjBzKdbAL+zKVdaZG6m7XW5Ba7/vp1rIXwduUO1HEQFKbY6+CrXSTg4dT
2OTTWu+paKzxrb+LWzPh5vscvgZ5cvjuNhyWBE+zRxDp+OxraDiJc1asbG2Ki0u+u67ScKPW9yla
1s2t0QxdQhrBPq9mrcUZxOdBDZLaptcVJDoHwo9ZKlshRbXaT9IKC8CePxX9J/GLVxBkTbplu9+W
z7DVRjR7GuU59g6cPYmlRWw9KLDSp3XkRFRq4ZjlOBT+RC5Ftl55GAGl55XCO7xUd3DL5o4pp3DY
pxZotixjQWCI6bRcx6ZefLbWZsGZOAkuvULk2c7i5u73OrGbXrc5B0UU13lnH3gRiw0uth3L3Q/q
QfI0mgdJJjuMVyOCS5C5y7ueMVmQ9ny6Wx/rgIavGGSBd9HgfsDlcnICpkUC4kwHOlXNQ3MpomA7
9V0Z46MWWU2PhViVBNiZgvTdaqe1UDHHeO4vh0E93RVOyBKJdvvoXtEx9RF8WovmNhSsiEOMxawF
ym0+dom1TwGGfwW3TQRfvg347BknBEEYkAr2SUJZW5nE+gNptGT6JPaQhdhwWR8V9vk2ige05Iew
xbZyI3gGyFsgvTZbmrJwF0VbwcbvOz2nCHFlQw+2USNxUFN5cyrfBUkIgo8azWVp3/FmLJCuH2vv
p1ZfV7vAPzFh9aV6+XFROLcIzuy2ehIpgujPS6kTyibYqaUWUsLKqK6fUfl+LAYrTL6a1OxcOXVI
uh2s00aUEdBvjpTm+Atiwsj2shAEiom8Kn4C0RNdL8Ti7MVr+x2xy6ZGwHmfysv+Y8SubGVvTFv8
iHU5ouiv+cHx8yKSCmE0lOCejc7J7ytLC8a8LtByUeujhdZ+Z+8AaFeUNMuDs31E4hbM36hF6ukx
eyO9vHvxyhziYEKW+keeb/HXrJ2PabPvB1z49GSP4cXgJkc1qddi+3CiqIBxkpCjDejT+lVWj2t0
cqanboIpoe4WLa1rCwsTOQ5CwhXwSTCVJQk5mCKJe1T5a8bzjpRqU7DM7QM8anfyIGyVKBcAFMkm
2ZD/RE8onUPaMQtdcVex3jnNVWytSa8krS9G1SNevPRSUFuL3fZqD5oLdYsExcfPoSJPPN3RmQhb
P+Ug/Yph9sfOlpvCtZ4v6CcCp5c7XSiJLHgOuGzUzyeAQcY4RouHZie9OW0UpEXUOvhCw1v2Weh9
oCsA0/GLbHEGReDcnRPy3c27qc2QGgJuclaCfHzGUiaBRYvWJyoQsi1cuHER24LOutYWEOXSYCoT
EiXxpfkGT2jRRav9TJE25KyViTc2j6sdQNVh24XWCc7uM9vQAFOZGvulRoWLBRgJRAm7tpWigelE
HnsMoqTPblMcVyr2GcofDsOJKF2XCmj9qWNY8SYQxoHmhWQDdn3b7k0N4KbTPreEP9kwrZtG2l3r
/+6+q67o8WioRnFQujCoV8qDI5lOIZxYgdwqxNP0G4kaiZ7EcnddxeVmsKDEq0g12IFiVnbur3Ff
Iaw/gsaM6cHFU11WAqhB16i6u+SFLfCpM8ee0TD296wWFLhdhURDNYtVJ+ffC0p/zscf5q1LeNYo
MbNyoz11JsVERlEObXTlr+u7zQ7fn7xi1OGPiNt3m/KJl+OSPqjMtfmeIH+U3jhngRA3IU3qfW2N
/XPl4tc+HrD0XXemWp5dKI+scoWRkTZ3TUYKtVhG8UEh89WLQhp1PY6tjDzeghb0dwlYYgJoi8gD
uHr12mm/Tc6AobZFw0ptpJH7d6S0EmOjdtEKwFxz6OX+wnv0tpRJNCVYO+2B+NEdDEd36FYNjeik
kdMMJArz0bVFpKOSi4FoApAtvLN5jXslWgApqz4DYPxAL/tmQJhYkb36LD6dP7EQjBVSdZ+o/Z0C
Ta6B8gv1xYE1oLKed4zsuCApPhf3t0LLNrGwj+lm9MliVgwpm8tUjAIWZQjUqve9hgnZg4LV7mVz
SWGFMCwRbhnvePzN297ciTnQd+0opudWWAlbEMBxFEm1vInhHnVBJabefTZd75wKxAPw+yYIcz2u
nbcABNJjYZulSs3WseEJgy5UrArprZ+rR3aflU9npp0wkb4DfeWQZ5n+6uCSqPsw+wNadVdaBipR
vu35bDmxzCUWSiZCcc3xllbsH16DcGuzAsaGnsGR5ZIUpF8faccNtnf8wB/wDCcA/xVRGrZ6gCWd
dBLaHb62y3bYZGU1D/Ona9Oo55iW6FsK9rqpNtwlehkSLX4ZKkwXTy47VK7DXvIJUYnFtO4d3knR
uFz/zbiwXKiJ0UIom33KEYLj672HUJ5VvB0AFAig6VFCys/Ri9pfhu/80U3MU/FAc0EJ9bCGAQox
CllRUWNAP6G3v2FV0mHxEralF8psc2TEGxu04V5QqxAOhtUpaWND9mwQletq3WkL2rRdtpdYrwc/
WPuSvBH2RVUysuOZYTulbYMSHqPGF/e4hObuah4YWBJFin6FTKrxxtnQ6q+gPTzm8vxBjyKPc5sK
s3t/9MTtMMYKxl5teGAxyW2ohp/8+Rel2jOP9rU/T91Kcoo61PI8P7W/i7LV5BRcZqhO5ZN7mUrq
6i8L6GcRV++k8fp3sz/quxbOKTqSya9LrcezkjrVPDOBWXYyuf4IPSUW2vgbW9ibEZPtdxBnb3On
ihR67kbkkdpSOVnk0MNbvgFka82Slk0P1n2ZyYZZbmSk3ccw5dDHtJ2syJYahByHxtr+vGoxuQRh
TNVXAOGMTuRfXtrVVNKpXzIf3wMY6SDAAPjDsSFcM8yNnueKjHOv68mLyjo/sPOvEmDaCNiqfn00
SJYL2NOIC8kngIzR2l+vfZsCQUWSRgiUcMEu/wSWi/8+GJ5BsCQ4WRQAr7aJJHPOCxeZhC3LrHpu
7cizxyzEGoSdNbyemnIF5yJgZRQvMBxatffzsjBUhbZ68TxW/KiTT/SvAetzoS4di95G5EV3oTFH
A1iMBXKV6qePeXho4x3RWrrcVKZ149JdBi7zVwD56GCwLK6ZqO6xug81ipd8fbL98JPsb/3aXzM2
i8lqnj6AJIK0G8RgRG6YnLhltcseWEoG4E+RP3hHTiQNqHlQltYMs7yGcpPvBwXe7m4/99sY63S6
YdVYg+/eReI7YLlrnU07ZnPpvHUcBxOOCKE4XtvXTgMmeBijb0j33t1WGWEBg4EiEqyFeIZzwG9I
+8fDXqeg/4+DMfRZ63ezIExfJy3DZ2FYmc1cULuKJkbgrxgAsdfOmtjq+h+PgmDSOZ7YUc4/SGQH
ITxiW0yvMw8NMCI7XfX0BqILqyewIvjbcFhbPnVWSlspQU/y6gGC1mRjwdxxZMMSPPT/y6WR9GX1
F2Xt4nHwf0T/J74mcG/Oo9WJcolmC/9XKbAOKoKLLUaYFY5fsGfTO8/xlZMn6iO0ALxAkRAZuqXn
NdYHVROUpb+106LZMXpxG1fxmh3ojQ+pROPIFi2Q/PEfINp1XojPYYF9TKsEY25O9Dj30/el5fP7
vzdgYQ62mCkR8tN45t90ul7h48UrkNm1c/TL1bT9HzLQh/+MRdZHdQ1cC8RZIljDxN1S3hpdGeKI
Nigh7MuoO88Wh3UJjBJoMjXRz4QRxpACSzErdVKbv4hmUowFF3S6IHN7Rf13NewV01xQezZxhEVp
q1mNBJZtpkdKNABAa6uFlPqD0VmMgfVw5B6EZkWIBZT+lAZYGGTBxFXiPxvKVpPgsdW9wO6WgPN2
Ngg2SUGLptwxACWRvHe2k8GS438eiaN5N5OJBb5vI1WxqoUFazSNeHS74Aw8U+vuJUz8ey/refiA
XX/U4J97ZJIAgVIcXB4puoiRv3PZDW9JqQkW4I9YSzRAiPrqsWzq57U1WFHR0+VLkMpn/UTujkjh
WegnrYM/sh5RuuqMa5n2EkimPrTH2Z5DNf9GPMBadI2lZ8dg85PBy9GN2uj0LZrXjcP3PXi6Fuxd
EEkR7XVxmM736lWPaBzCcwfwXCB2VXz94Wxzo1gnqQq7cQCkiQl+iaSs70FbSWtjIOqqwJLMBLLu
XTbAAQtzoXSTrMQvsxCGVwb/24f4ezAwRf0GfOywaBMTN0BvICTZk8+rH+jiGrzfaeUX4AWo+hYO
LXSvNShcm5u8FWsfO/fbKHeDAvrPPbQZd9Os/ysq3v4+2GegFhJujV8V5RdDF8SeQoKaCzZ5Udgu
1OvqYHRFgZvQe4Hm3ribdlebRYnj0Bpb4kqfN13TQ+Une4gwcaOr82N5acCMsyBcpFMbiSfpqkNx
WyqD67NdHOoOqMNeFOjF3CFrlMbLQquulb8RCCyf9JQ4S4C2CDYj6EJYrF6IGJEp0zoZrwXoBWBD
3ifXhoje6RZoP2GsBY0WEcFcGg4J83qj8+j83An0zqcJQMMh2Ws4YAXTWjaexppLqlOSl9iQjJBb
snZsZIjwqxG8s2kRDdYkwkP0mTpuD6YiOBvtggGfC4ydpMGQZGesoeoFUbpqa7T4pE+TrM4u4Cnb
JRkgUhOVwaY1BavEqbx1uu8blSv3+UNuQPznl7napdXFrg8Xghj5VjvFWirHGbRigVi8Dnawythk
F9DCqBEr7RPkIwHa1iqWVKnaN5E66lW/XdKCkusRAeZ90pP/gfCE7fTa6sjnM9Q7dc03pS3ARAV5
ep5NYiH5hmAMStApVJMjEaFlidw7fQ+d7JhQV0esuvz/evTWDoB60nn0LtoadejkwvEi2PzwYMEX
rTgp867o1xdWU8Zx1F2jOiBW1if/MRrv7wOwIDq1fUX1Bxtqf56Vwue4fzkPiqu9XW+BABmT7yjo
/COAagM/yIrz0XQmTPdmq0HgdBfqxSF+fKIttvonRnh8N3kkGbS9KU2iYkq0H2tqokl7b8dejJ2D
vCFAibq/A0Al9eaRQMgi3Hw8p/LppOQjVGAv21/udH2Y/UG6nYv6ye2ZtVfLznPZj2B8cL7rqTmt
BEasNcSkiX18Ucnzd+lp36Ex4UTEh6GL/dQbeJqOk8zei+RjbrmxrX0bX2PhzD5EZuAnqHEOlhgE
OLfQWe3FmESrW/u+HpRlZhHw7P9oizFp2G+KsaTEuzpT2pY+AbxixKJLGm+bEASgoeAmomRnGUQT
3hcvuR3F8oyOEBVcZoSVodmkG8rJwUIyDi/yQo1D0Xw/XFZlIPRmKP0psqEH+fXELDQ8w/IaJNts
X/yOHOp4O0vPX7PH7WnEopzHdta09Ygo6v32xUbt1Fsivhsy7hEaPNVtKP1cksRLXG+VVKFd8WGX
mn9TUF7cgyksd+m9uAEQBMr5SEPGXjlg6CDEqQJ6SbFalE+hMlq7trKNzOhP/oJMkCZn/KdwFMEa
jzjruxEVa4KsotTgCG4tkFjk2GGSW0PDrJfNmfUo6VqbBMNHJ3U+a95geW6pBvNo/NQX53zsL468
VpXHJm8+wHKBkAuPaQELGSICvkU9jcFvaNRZae6eL3DfdEgzP/z4QDWklxQUU+O7MSr/IZS9y+3l
zxSW6j5E7rIiz1a8iSrmN5UnhOI3bisyhPgiejKSwkz2CgiSEx5z4+rXCdqKfXmLitvw5YWARnGf
pjw//iucanZyfH8mA60o7Xi3GClIikqgGo7JiWgxC7JWUfHhEpIS4MQaboPYC6Y2UjCn4dP5YjAR
fpTj11KE3LY/QA3mfKyi0U9DX4ub3xJdyQLgi/lciILapF8OOozNDEU7aU4zBjCv62jixwEfv5X4
Z0gWgKo9KIaRzKbzdJIjJ4zey/PYd7A6lad7KInr4AxwJGbYVhhOkGmSWX5vzv7SiAwfFnNOAvZ5
jWCAvBWZ62pwbLBoMa3hXTHgqvY7W8FhQhcJbZ1nQM+17dkWxrPbXwzVYYwOt2OuZ36TSVlx7kGJ
YUqPJII6wElrj+hrMdaWIYt5pk5Oibh00JWzNX0ZV6k82QfmdXwQjoSUWLTVdywzkeQ3JpCw+Ywi
aUD3X1Y0i3GSAewRO0IteiDEoBQreaQGT16Or9d8j6tY/KybLjEq36cmTBmq+wY0ubaq5OapP0IS
xChsxgg+o9vBZVKBxMgvIEwZlNhDJFRhm/tXatCiZLwCBhsNA5VZAM1ED7MTvPBHby1naQhVvsN0
M1w4OxLxHiE2gL4Nyg8gPbkxlKv8+W7eB94YnZ2xkDbx4QMyX6WntR3iJKwDnkrqEYQQ3MueFoaQ
7OggBpBRpxPceYuX5UQgA7qHsI88FMWWLAL9f+7ozEYfyU2PsDdT2Urf6Hu+Rr6QfxZk+MuY6imq
RTGRbOH8/FDO3hzI0z+Pa3j2YF7y5/JCdsny26LXhcoqjxBwIcz5OeGX5Bc2KBt26UPvPtQBhkfG
md1SwHbA6Ms43+O7DBEPj86/BhkCjxHaV31tFjjkavt1zaycVtG0XIN2lxcZR7U2hY0rpTv8Pgqp
/IKpksHXv5/WJlZ+sR4rqlt9ywXZSJDdGLCKLjjYqLLmibkHMl6uzF0ubfbr/MGZU26pAFQzKX22
iD5xLId8ubinqAjiPDFbPzW6hSPdqaew2ntVInG9PwhFinb8dY6nhLKH/fJ+QtcVhw7/+Blqa7yQ
ypkbaglfx9rSj+lgmdla4AkBhheXpdJowR8X0bm9mp6tv2g/AGDS/gw5Z2t3rbc1gm8ppvo5sz4q
6Y/vIFoTHZF9j5QaKCTZYlTotJn7yPt8/W5uPUha27jSxbs6eAq43cjr3nL7fP7mwehSOlH2pBL6
iNb/w06eKBCatPzxLDcHZ9nMvtzO/lDyzHchEsLvFOXtWWL8T7+PcXQGdJQoocQUWnrCcLDlmZ1V
JvuYPR9wczwmWZx2ihBzl0MBmEd+skeJ3i1n+W69yeS0HWVFe9AN8tgzF5Lq9pn8OZsjcRIvt0Pw
ifaMHMs9elreSnRHMQSyuOjz2TA3/prxZu0TdEaGlTfS6LtgRpMMJ+XkiS7ghony17Qc5K5JNHTa
QXuLrHFCVSVxMRIPQMHWikBJrVyFv1TWjNdU4N6E/qDqVLXuuR8IxSzn+IaVG7gp1LbczDTc4SKf
RGEw+eg3QfBUw08TuWOyCMYTMEkUs+2uFwE1HPGsCGrKZAdNLt22IQwdeQImIvWonrfk78HG2TVr
yeD+xg6aLUgfhAlP8OBrg1MBx/NHhWVEeB0NrffJZNMAsqsQoTBMBB9PnVN9HI1/4HkFUyq92iH7
HWZWUoLD6Y79cPMPOc2eLPYqbnczGXJAM3u8GP6N5L5bhWHky834QaSIthArHXNdc234K1Lt5/er
1yjzmdYkzxqrZxzrgoTHAlYnv97ComjW0m29jDkm9DvWGX6OsXFN4J3PaSCUcyy9CLBXlkaoLWQw
dhR0uik4kkpg1IX21gXA+0d+w9CZc0QjJ1OikT08NSBVh6WPl3PyTUjqqr7F4JPFaHKRxIDpTgZn
isvqShtfgmpNobYtljfYgWvzdZVYMfRGp+IYCKKITEHxusbK7CBkDz+C0vjTe5nzLFbMRhv6LsIN
uA3SjOHpN2oi0qcZFlXkX5q+kUPJYniY0BxYXFHfTmi4KNqzBoWKUk1cJp2J9fQ3P9z4tOrVjuRc
HyLSjLmIyWYBRm8XqeoT8aAmzq5zwcxXcmXnjiGxwLS4J07X5LeQ9OfopybzK9OwPrlikObA63i/
fcjYf9IYNMBVlfMgbeUKcCcaOKuf89U55cGMMXj8H6nTbfyz6V/hB9wzbWF/FaoUmC4eFRzAws9S
ZmWdSchu6HNs3gJrIR2PMsDa+RA909VXIMou5g5Sz/yp/QWMZGrJuojwNfvf83cvqmhu73O8ypOD
w0Aqypk8AbHYOxoZ/waqOAGEmxwCj6syGaqGqmnXEjux8+Zfzc3Zc0meAnJ1tltpTIoUU0J/3Y4R
b4e5kTnck6HObjCxzrbsxlVFQIWe8M+xfeufT1zIb4eQcqcaYX6m9eEMKASom4YN9VjdGeIT4GEf
+Dq8synPq9vO7AJcbt0NSDRKUAt0ly0bJ3/ECUKLw0HrkSU6XiycNXjNJNljN2LTq2x4r87RHT9p
g108bC1PGz52ALSRrIxRbFRik8LM10udbtknu4aYaX1D00rjn4x96NFPnVB7L+r1SuvrlldxNWuJ
yl+6wPxiZLHxF4IMe0ukd0Coy2aL4iU5FLzUWeTfpU2GZR0iyIQbCy3Mv5NOr79B6zwDPdafyHeY
EcUtYiStl+10O+sZHZylnTXuhu4djqBkcRoyRoobYSIeHdlC0fHLPGX7zHLKzNEhLnQeAt1sWteH
EKucxgykQ6K/aH+IWf65X7sUhXsBPwHOBy5RSovXuh+EmMUIyY8Zh8qtzsSvoYm+b0+IHirg4OGJ
scYcO529z36FYjTAW1bWekEGWmOj/3DVgvtCzld7yj9B1W5OsQH56TNlD8ga0yBYvoHlbWSSPLE2
QDTbVCmKVr6NN1tQ6oOmfJtIA+Qsl+RCL4xeVaRboLDoNIT+VMVsCkKyPbGbdoKFjWOT6bYo4Ts+
YglTwIojpLJHoX81xRNId5LWkTgecrvi4f1mAaBi8wkO21bh8fySCE+QhUQoYrsenKEd/y1Ib2WC
36ljaU2UR2IxdHU2mOu2qkKsBlgUeQreh4iugWVm4hrFd6iXZQoa8jmbIVSmTaSMJ+UDcOIliQZh
ZFONZiQwcQS+mcr3khzmR+nJ472eClF/U9J+lUGrSGGwANnGbPdriqRWEt1cZsM1h3BjwJm2h3KF
WFV95VwO9kN7+i66ll+xNfFZhzRpsuE4Q+V4LA2LPNG7vvQ1lT/xUO3Ik5TgntZT/OhfVFNFOX4z
yLQRAv/EOOqbmJDquni0oAAH7bmmG7VL/Cng4LZI/ZUeyDYGaS3WKxZg1jm26miNVgvi1altySq5
bAh9ZF4W1aldbL1WyQ6YG3+6AlvQvr4GxOsHlRfu6BmdJYdVLvkk8cIhFRoXsgIrR1K5og912U6f
4c2lyA2dkFEX83spzDqxNmgU6nOLOt5Xjczu8hhayX+LryAKvef+DNjRr34/LxuycBPd9dDBvZm1
NIPbiMsOrtViaFWLTPXgOaKVa0CKfy23P8mQBI4M9QPnAcUlWflxchwu9ApQObDk3/fB5SLKY1j9
f/PcLNvjDSGTGssJs4Z0OhWJJ97pHiVUWPUppzO9YK4sxGdurjSzFCmgVpGMn1QxLp0tUgMNuyza
VaBJTjB+GI2qhCAqq8UcVNvqovuITYFpXADvOOhZI/24XNWYm7ysJHWblzWI4c2OYivuQyZHQlff
khXVpw8V26hCg74na5gAOj202mJ2gOmOsnQoZes8c3EqdeVkkp8zgXRgIcae87ibl6bgGxQjmOup
vDdc82uuOWacf1PCw0pT3r0kO41IQ6xGC3vJBVuDs0f74Yg9hnkNFDWgQ+YiDuk28vNx0n0Pfx3+
ictZa0ezDbnEDyjxybyPabzgDOBW5khUSUS4uX4t4wohUgGPGuSXE49rbgOaP+B4bjFWYF1wEofj
7o40cBa38R6PFoDITYGOHKYdTpdLdUGtWJCf3LgZbaBn/7vsTkrLOvlmSdtf/9gqFdMIs6aX0ohD
eXff3UAz+966S1fTOZo7VDYonpkfdgvnP1Hyl9NszEvJGQJ6qXtF2dg6zUEbczhhfWGdc4Sdcvbh
pptMDgKQHWL+pqsrQUaMtHQjWVZAfArzwFb/ZOithW9FFodXc1rTypukU3BGQAYPhgB03F8hBM8z
i+0Dr4tBzi8DNwR2RMnsAgfvR0yt+FZgkqQN6TZHfw30PbYe485yDbqxUKAT+2ACrfL91vj7wmMB
GG73WTjCOrGepGa8CPKjvpfp6aGeqripnzapVfia++2z5XNnWiFH9Is1F1jx1igqYuCs2dA+Tbbt
Q4/Yhd9hwHnqDlCruesMHSQ+mzMwN1/knnzAzBokV8WKNPMpU7s9GcPgJlEHdz8cm/Beim/JJrey
rsvEY5e9ML1Rad0Ulq8zFZc/0tu5sHLnS2vbHeSuJKUQ9CgKUZuzRnOssl2P0uqd2/7s9uy39X55
05iaDXDltal37ZrfdhPm9TToJwpopcyeRJ4qOJ2k2uXawreNbk0wUXq+82KmJjIV8yaok2JxqAJQ
oVrZc5ncyzImGT4KrrXEC0cMKMPxI6dXUL7bCVR6YTQkug2w1x4sN/AQPdmNnvieoNkSkJeRWHc9
yxofq9w0rcPcbquiq89Txkc2tx2dmRsItTh/FcUZLZ0O/fFrELAfiYSmNqbccMCqO4Rzv/jzW01H
hx8086MPuqqKeU18ZbI89Oqa7svrV8ARb/4yA8y2VSQvLYZh8PtglW6xNzXwxYR80y+PVvoxSMLr
bs7I96+IfzP7yaeqFTo5HPrDU9VClAgclwUybEYv2sUi3zeJYJfNuc82UMR9zmHmPHQLCy2LwQaV
Tc2sj2Kankpqy4PLdH+KuDUqfb6l4+h5j0+1Zdr2GoduoG8Jyc6MM0q7Cfi6WkRR//SiuEpH1GCl
YEA7ApSE8n8fWyOHyhrbPOjv/2mkDkL6wa0oO/wkgXyro4wrOzuKBwPp1CHLveGf0BBGKe22F1bu
59obQiPPGbNTFRAmnVg4ZG0lfrUDKHUNtX24CjEbFJaJcXBWxK6jalmYwMD0Nvpr2le1QS9F7v6I
CsUdHMC2POab3XxAtRcdMGJXmlNZg4xpwZSKT2gUWQgXiu6eRTFZnmrb94glSEm2AfXrz3nxeRUr
qtX2ES6OpjU40KNOWO86BUO4W+3DmeWh7Sso9p4xkXNFao6PWiUk42JFgZFnRoGxND4CPnTkJVJ3
6v3s6M8vggYb0f0Kmz28q3YpMS6H5My7UgjK8DDiK9J9W6bJQoWJjsp/5cv4uR2jr0s+xdYySnAA
ri+S4rk81mzJsOU2+A2ZrvlelKl6cprbfFF7LRRFlnhNxo5KQWKiJ8fX7mQ2W7jdkUqrxjea3wNh
ZrtMcXkr8u5jDlBOfCJDetmDQF7vExzmV3qgO10QRKzRvGp/GA+bU/fqKc/Zor/LfluwMOBgFRIN
o486PL3WzusNE/wXhCHHmb70IdAxZbHRpAH1/0bmKi6qdUozzP/gLUa2r+clvm6tDfOiNtg/NjZ1
jCXyeYSNfJxp77TvkG9O5ZCEDazI4HlUW+r1NqRXgzG5JxgYgLGUZEy3UieEc0i5kkyitKptfRLT
5fWlnx1CuVjE6z5DBz4tgEhELI4WHyrRiIj8wYtsCu+syUQ+T+qN4BrWpJa3OnE3W92qfIlsH93W
d52PABiCdmFnH9H6KpOkKzIPhO5+8N5mYmpgaaBDXg9gvQp6hFomFQVbXdSZQQInIvcyJtXRaEms
ZfYd9/tq1bkeRqQiIUaKge18Trl+lL6v3dGEj6GE/ixSt0OdlefWvtxRNiCiWBCrzMnjObwi2Y5w
JxvZpHu5tvOI7XJsXa3+Wgw+nX8/fqwkwRE2jmsoiyQLghZ2eE++Wy1L+UfBzYXS5tOEoOrFG9QK
bWShvwRlnOeW6bgFgMu4n8+GRmQ5+KwiZMzxxnCeLHMP+pRJ4g7xN3tAc4MMM6xMtaphFKqyEjs1
bv/n/c4xgNpJ4ptywD/8kHgvJxkreWJHRY5WoT6CwPEgyfk13GTa4HsK8EmUcAfWgVwQZIVBW8a/
Uz7zLfeHWxIjv+yp+FXCPXAgjj36CiNTCOVLhnkcLeR0+3G3f6HleibFNDqODGQv6bhJVSYiK7l9
tTZyw9NjKq8K9KAmjbzqdLroc5FJuLaxShk0wWP/g8cLAwqXQSpa6mW9vtSPM1ppp5u5mnH7pqSb
kRJ9ZuaOny2g69g9QW2uTFZNfIc2npL+DDP3KW4By8ADBAxZhAJLhJtwiuW95rqz24dPebOaKEuW
RVTk1mzSiDoMBFwr8K8NU9GPVV4fARPFcCqzYVLbnOLBAY5O7P++IWbDTmZSjNxWg9sWrMeHyJbO
fChtfe28s9HHMaAC1sXTWJgLewQFcQlJvj3e4HcBF8CD0XxeFfFvinwq+2MVtaQPKwkelPdNeEZQ
a/Ea2xf8ww0B+0Rvs8FFmyYn812fhuEgEEEnq7aUHK9ww458HrPt4sHQb29LnDJlk45nxc/dsg1g
or8XdHvr7/HsA1EnHQk/s+lUH46xPFc//yL1pWTzG+CasqAd6/Kx0EuklZ1/+9XAKtwasWwWncNA
cqiev7qjPveBm9SSiDKQBhf21ZOtQPnJ6pWSaXE1pO2Aj3N0qfPT3JKrCJgM2bcKWxg6ow15TDK9
GnoN7NGDzoiNU1dwKpDYlrsTgjjnDOa9LP9v9cex+j0fEIzDSZwhsy6xQfpvepvY94TBaP5A8oLw
+dIzD9S6AC88D5KV81YdDmJiLffaU+vKa34LnJbrcrHGXtJ0Uwqn6LnUl1uwp5Im5Oz/uvmb18Xj
rewVqbsuR07zmCDcsU58eBbN9TPjou5rMxVvG8bexlTtLxKb0ZntnL3sHXq6w+kFYUOZ+zx35SiY
NnJ8EDGmroxOrOiUZECJ9lXAnHRA6V6jGIKnDY87dJbkn6h+W9+6vWb/oxW3LggkMAwnKadsr9kG
7C+cd3RSf6ATzhqv+jCXUk79uNPUyeQr4xlBNWeW75m/tGH3gPs9csYW42dffim9ks1MKJY13s2n
aYohq0YcnXBFUFAAmTLZGXPERcUj/a0/Ulqrr4waHUmsag/+Q0oCyw5e8fnHNPCn50izDrogTLqw
VLncsXeB1vHLnuV5MJ5zJiuRqhx7WFvluYHATiGdluVLyL84E8g+NC5NpTksL0N5NoA/rjyjdG4Q
tvme5w4tOHFvnuRalylWd2NxXlV/do32+yh277zVsnSGM7f8B/qnneSFsCZuaeMee6Awn08HKjrt
sgHaSaP/xk2Y76/Le8ICcz3ryqPceqqbC8iYDUpIXMQkz7/P83L6hoLSCYr4Y6L0XysERTBBwEkY
PVrENTnyqnd7bB/WmQJpJmBTNlVfl29wkVxfgMzb3vY4aWsuNT8XsGDUr9pbc2C46DT8nB7RScoi
Blxo1bNUElCSYyw0UikTBRGHdvRBm7N2BQEW7WrMSnon6PZU6dQfW4tl9MXEt9Sy//LlkaYHKupQ
VnZUixaRcRRa3tkmuIp254x+yOrpxVLJCWucmdTeTsjrZ3Wwdr42L48N5oGYq77caAkSd4adKY5S
B1vT18Mf+h3V2Rug32JlOTKpGglZVREs6pq8JIPsWkEFRdbDx1iASj82vLnz15XqO5S+kTd+8L5t
OtMpud3aU1jk5pLASKMwxfQtRPuSFKk4ucUu7RDZKargrI1aA4I8qf0e2sn+7MjWE7nGokZ7ViBQ
NH9EUg5zk1BOqZ91vtevQPof7EeAg5vs1NCzqZFK5ssBSPo6/HH3Gj8lfDWnuW8NX/hjGPKU9h7H
1n+u9qRDYL/pTt8L5Bo7iJcV3lXCo5hKGp2L7VXvx155l1M/s0JBBE6hUUObcgjIf+HyM9jOlEME
i1jSxGHaJnOi9sauZImKFpJAvm5/inM8DPlAMDvy811SJC4QzmAkvxtTfUghF/9uCjmVw/OZFSch
l6JueyKUlRXvqdgsPvZVbyt/rUnoNO5hozb0e1P9nOQHHkHC9wIltoINDd/Zrs4+Gq+pZKWkdnpg
dvwvXa+yCeq7BT+P6ja/UcLAZ7NFaU+B5I3Ux5eQu4buaiWqd7B0aloFlmBI7z4HeIKdCXjjoR9K
Hww/m9YLk/PLGmkhPOnGTax8zAWRlJ+d0+Qg85I1G5pTn0cGOJOpsT2NesbFSwJxC4HAglRr4yew
NTagGFrLDG3LKwoc1+4TAma176kKmetVTpc8ZBbaIXW+hChIvzl6DF0qNH1EErJahDj9t2XxEMwE
zKaeoNaQ8JRQZfLBBl6YDZtK6kadvgI4ndGX6y/cgHMoitmKR4G2X1AvdRtMnBMNbW9Xz+a93Ifl
8IjdrThEszlDGQus6pN3L83Uu2f4Djfz8PKi2OusIih9IQrZ2b0bBsKt7IxyuizLx4RZVhUmPSiF
bJfd+ULvmAhI4Ahnoi82P/l2+lF6u5MTZgta+Qk9iG9Pramzha5KkiS416zhcFGGwOul4MmlvCj7
LchBsKT22eLyW5RNsJ7mUAaw1ETWg2GrZ4CTqL5DTudGO44IySjNwW3vrD5YrxCURctL1RCWtR68
pHAa50lTDjLumsltunD1Mn+w/n+lNX7fRxZvGuDpukzQrbQ6uiQgJLh/KMupDT39Y32xSdQDiVqY
WeBapkSAroi50W1VpbgNlv4nsaR8eQvEzIHI1dr7vI6oIu1dQWlVUnC16J00yuHU9dHRhEn4vKie
gZgU/PG2H4Yb4kY4VeKx3u064kCwAFoyl5v/bdnAjttDI9JOznLq+FGD2Zv2vkynRnXHtGzuf6Q8
1AgzusyZ13dktMnXYjeQs5MGPcKKGGweb9S6uIyQw8oXvAVKgp86/tTVfLxIHDIGqBztVldZ7/xC
IAsHx1IaV44qkFdGd+NoNb/IcWizbBs/HwMDuLJ5SZnDaQ8+42WSfL5zjw4yU6NMgcjaEXNLakFW
FQv237VWibhbrJ87jKCWZ1b+DjBQpc8GAdx5C8aGfiH5neHhTswRk5zh0jlGpooNx6Bn+56jazXO
FaQmeuKLZpig/b1Mk/mdtAwotqwDjfIF0PPjCgoOGcpjE1Hl36pF0ccuHk40P/00KjwFNrmwNpP7
S/Db4MbSY3OnAnJXVoFbD34pMVOOSwJPIX25LD44GAs2j26mDDUw+cxfiox0If/9FxGDPNVUfE2c
EiNctqRhx6G8C+pk1z/Yx4M1wGsRmvHH5BQFyO2Wz9GMq9mYAD/aQ7Eb/vAq4oY5+cwOeHTQy5wc
08L83tV3D0WeSUZPMzzh277h/e32CurZ6oqsKeU5MzT/55kJwAActYVZfU3TCGAiQVN3wkrKxluc
/Awb9KLsCplgzCGqkHOhZuDzfPJeHP7I/ljhRnhzKS8pdF2Uw2yMVV+3YrptQI1gw+mML1w2eEcx
+98Gr5AT70hdutzZXp23euf0WkeiUEjqN7FSqYH5Vq6TaGT43jIZmIT6HC1czdEVF7HzbnhC10A8
NkDQQgeBpbaNMvVlZieT5Ue80YtGMcNmzkDOi1ESgdb1nTjd7uFuKla5BMoPdc8QrV4Lho8Corw/
g05rf0YFJw4pn9wIOGroC+m8UPSWeYvzE+yQRXRyMOPiZOuyvPQef+dhd3Hmw7ZFb8LUmMvNrh8j
C4pPsYlXyjRCRPxWpROy3sAtRFNc0JwHoD3BfGa+cx1R5QuzNNKT+cmzFILwxFPSaNWaRrNbTWvB
23KbWU+1XRT5bc/ipJtgVaf4FArrfgYMovt2yDePU4vXu32I11gTnCom7Rho5hRyKrye87YN+Pz5
xUsne6FNs+/eloDv6hx2PPGUb1MNTPQnYUHn21gozZ7MDjgdkBCEFCgeqLyVjhFVRNsbetLV5v0/
ql4G9OJlOlZY4uDhz/OBWu25zOux4RUKsPJs1+3PZtNo2rFKRDWJGrut2akO6RDX+cx2UJ3JUnXt
vxfWGjiwmSrHR+B+tQKUEqy6zffdesSfkuRj8LEgnvJfDDL0LqNKoZfzgl2ScmVSGCFEzNMoXVQU
th01iIz0Bz1Iz7cY9CgJMuEPTjiz1hot/M1e6Fr0JlQAgeynw/VuC0Mw+dpEl+1yVRZsm0NO0TT0
QxNJoRGOyYNnXjzmcW/wLamg9+Tkk6t6L5Gz+w22KncoGZaSZplas9P3AIKORfl5x8YlsGkv8aZd
7S1vIGm3O35iOpem4wDaf1Cqj3181Cl0Xn1hQI1eLa29mQb29SPCI7MBWORmwdn1jBa2xY1na4ve
RKulr9iDMtcsjbU5vOiEi+xEVYHKlM2xUbj4ewJPJYrbcwpVrWA7N+UF251aCGHoE5qWKG1d3qqU
bpzKRSkz242bc32uqNfy6wlTqvXYxaax6QPeV/FiuEv/DcDoM/clZUiDATzbzok0Qiaqw1EWBtXt
tOJCnvo4Es6v/X211Ew30DkBq2d5Bbk2pxBlNFIh7v23V2uxUfPDjNtJcZBmyctu6Wy2LkMcrbJn
9X21nOQW6sFh/XxgOQJ29oTsWB78Vwn98vEIM74SktvdaPioJmJkNmqJpurTlkl5Q20FJzG6BclR
twucIM4uSgsJvVUWUOgJWohG5MgPmrY5ep4B/1yxIsQVaIvBvQW+4dYfitUFwYmcWz4FCuUGA9M8
RzgpvDAzrz2OO/wQqrF/1EiqJlhZqBwPI0wo7HBfxkDEDoEOcy4BNsxnF6wIGCluqTYrVtahYhmr
sIKdkMFOnY+V7YczjhJg6p4YhIdRRXi4yRkiga1lffMRGbfiXtuM+vJ3vBkyS8XB4ctE533RSlVk
iFsGo91OAUzpH4fZKoa3zqoWSzYm7nYODZaNyxeEq7L43WFydAoRa6S1Uv/2wAdt/lzJ1iPZePE8
NG9dnSNdC/u74OCfqaJPkSvkgpryR+JoW0pTIM+qzCuHTucTOBfmNOPG3ThzdHL3mbsvo9X0dYqW
IDafUq+08LZoGU/B52qPJYFO45q4Mt0ZbJ1pwpgMyCgWnucnza5iUDGX8zRN5iDnPPGWRbMCNMWM
Mp18c/z962+Uc8aMjfIpXMtvUjUDr9EccQTfF3z3jPlfMe9ws3om++VETyq2/QaEcpBZ2enR0HkO
pwb/JONH9/cQZqe9h74C088lvlMR3XSUxg0otGXSSBp+aa7/+pHV6Yj0iE78DQpVMNddC+npkucz
zQCQp5EF0JFNzoi3eyqHz9b/17vtH40Utlc/ZG7pdTgli3+sibrurX5Pws2c7DpilivwtgM8Nt2q
yMr5Vz4VgJLsy7AEAhcP45VpRN0HW19eERAbzcpMm/cDU6frUXf0gTNCGDHDuULLD4fnsr+OU/lz
x4/cSS9X4tl21vLM2P01r7wELYxI7x1/73t7gn9fKVH2kyDARndndBIwAtX5wBGkbF7Nic14uJUr
v//PDji0q3oHnvpGelI36UP92LnwHJR/86cph9pnGt30aKXfyyp9IZL7QTPhCWy/erxl92vwcbi3
aaZbxkXKjaLQNFWGf2QF+IrHtoEQBnUrOqJKOx+Y5MC2SF2MtGUfDCryss8isReMQlM38FmEBtNd
YPY2wYNRsTux4IY01yBdraaeGtXCY3Neynkt/571rRcy/nh+OZPGTKMlicK5K/PDI7QcwxKFQHjd
/aF9KUhOqpRM+ZJlsLFIyq19FC5dZ0V2cjTncVvXHylT8iKpMuICVOVhmhf7km2w8ZGg5/ThNMfv
dWY9WAhz03WGfYLvyQH2JUVHsG9NN+bJ3ozap0soo4OqTLU5u4mR2oB2KFVDFq4Q+P+/Gm6vf5te
y5hrwtz3FzECOwuJ0u0HGFdV0UOv4+6DRCbXZzQlrgUlrtZ2WEd+YUzVMYO0hwwbfk2RnL1ZMYl8
DnFafS1kfiiMHVyjXWd/H5rom5vxG+H+hUz3cZblhCLUYLXvPVmcAd44YVicWEOjJAhknMEcNfu2
FbTkoJJotVmn6rIz4yYldSfOYMVvNjvjdE8xzWnVJ+btYZ2khTZCClPasWoVnEQPCxqWpL9FE6nV
91SNTWIyLh1pnsHDQY0NRM3OMPAzC2FRNqie3nVn3/vDfNaKrFXCR63MYUxJhQTk/cg3noP7B5y0
+ByskJMQanvMr7rW9Zx8MzsjtyqR2gxZObl9VOyKWPh0OdisZptuZiMlAnhY4gp4L7t5HHTg2lYV
FwRZA52K9n0+6EFztHcMUpOrpYH6f+rB6R7PLprp3OvbMpsz6of7Q+LXqWBSXdtNQ/TXwtTmSmJg
ZiBkCz85DIJhoFvh4JSwpItz5eFzka5hRh9J0gYT8ShzVgIqRwnbl2DLtYNke8mr5ubsS9WDkAwe
U9FQHD/MMBM90Y37Pg3/mbpjZHy+JfpOEWh2xEPs792y7TfgQKvqilmJNERC4j1kmMV5uDGXMOu9
73i+zoG6lHLjGmFyUx77irNtptpGu9HupU1W64BliJsq2wqEvB1cLJtMYd9YMLrCtj4Zh50tmf7m
xUl+xm2ZPer9kjzBM3jgG3XmUrhQPUCuK3wUWnr5iuRYx3/X+9A6PhHe+CUnU+i5lsAKkL2l91/n
fzjtTHXnzSFy4FWE0jif4L/b6stZ3kC819FA34z6V1pYRQxRzwMgiTNb/NmHdb6qr4ZUB2s72/pL
SL6eIF9f9G93s7LpP4ZUXGGTGt4F4bLyZaD8goQswg3rrkGcZCNwDSnbbkoGydK0oDWZ7VXCe46P
j8SkHQSRpmXZKwiSqSmQTi1aBe9pJy4VVvSjugnj98LJrhGZxsRAiajQF1JZNkpL9RFm5ktIe4ms
2y7AkzndrHIl4GPn+6rhwEYJy7k18EQjBGWTvQu5RLuM+PAM5iTNcl3xeVrLPyuX+Cb2npNRXl/Y
Bg0Fo+BOXGiWkPiqq1T/krL3ER3ZJOWqNrZ5/7NQhBeq7+diZ0H8HVCbhT4z4lOos+kspYHb34ru
xYSFj1YxZGQGjbQWDa77eQwcW5yruEmQ27m3JBUcrG3w7R4lK58+8u6xZUIJxftFAfWPcdBsuG2V
OhtrbtorsD8IcrFkDRb+1W6PTVUTxsnVZe8j5IyKjZ7hqjUXO8ePnpv9Z/IrWgF0kFaVqkUK12gn
lV2IGpXjFoP/3/IUD+jOXEc7OT4EYw7s0xeu/7r2lFjH6P/UQXL+Y6IuMtg72dlMxH+V4ZSYvAEy
A6iaVctOQRbDLU4VLolEbmDJHlL6i7vBisU8Sb94iR0l8Ahr2WZ5RvHQzZvEfd9a5Hqz7OiBTSeW
B5m3znZl5+dC1dOuFiYiDnAavt4JQbn1UMKweJUz9fPGW7zIbAv9cd3h0Pcs51wx5oc8RT09RM0y
oNGAjdrARq7zZy7NWlrHJ2DulWFH6Aiok+LwCWJ9x3kIiiQIRuvz2AaKdXSwv4h2n9TlVvXqKfm0
/WmJTMP43yd2ZffwuTxy/cnUz9bLz5hx3Ge9QzPA5EEWF4VXruKP7+hDWxGJetNGBJXuR+4/Gb27
PyL6wv4uOX8jh5J2TFxd1enq8GHekVGM6hT2bAH7kf3zH8ohq2cUhnfI7jTcCWL1ZL7ZeTY7BVIf
ejkSwNFwmK7EyjDNi49nyAtgS8eCoEHDEoiulw1xhZTLvMHjtZdgb37aF7DydI4qMw/yuZrxytx5
0FIwL9Uv4GwAK7JXR+LMxk8ap884QotMVeeq50XwoMSFPEaSzJi3vaPcJPK9AKdIVKAjpVIhFYMs
qNoe6igh1mhLUCcH96qmhd7GcWq0K31vvKdUR4Z6bftEaFR2B7r5qONqyDTTC36uHB2yjyu987eJ
xh2eFal2N0QIqJSggDuD84kh+RO0vkM0jGsKWj0itHD+snDjTTMSr1ZcsQN82eYwN7g3O6/rt7Ok
b94I4He2KfAJwGDooQlb2qdT26RB1jts0hgGCQAaf0REHJ7z+xEF8jxrxXZLyF8sBvL4ZlMHfioS
+YgDww99ftf6p4AuRqz1obRL1Z65MlNq4fIVvhWTYFSklyQpvV++tuW6yIcgrmj3JAcO1nQBrRhF
zt9nckr/8yzyFGR2ZMukaTJDYX5Y94p2VPYvJQP/X7vD+i31s01meg2FuRcfdBC+1JuL5srPgBqp
FATfOWOEP7GpPsGec2CtuLoqkJ/GwIzkjcYYHGuHxaTfVcxpOBREK0V/A09O50WUxctR/bOPjsyY
K1zDbD9120Y7OrtpXVf1lotFj1wzvoojXa+LWjOTeFoVbYRFZy0YYVreS+ZL3BzoHcBy9Z7uqdhL
hE9FPPkeZbiLJm0T2dlc3w/lhQKSKa2nzXyBt8hAF7xW6pFnq24hlP1TMj+fBLGRYdeRSttU5fvV
iJF1mD/vRiH5Wu8hTrr5eyDEJM3O9iBI1xc+RN1tfHFlJwyE/s/eNl4soDdnRqKtwVanxCPl/tof
ZcWrvgnQcoBoVNwzIn9aIlgrGIZbD72xF0Ii2cqL5sLGjAJDXoymBMu9KRe6Dtw9zG4ysM/FUUvK
crfBCuGUe1pd7f3aKJQgi8BsfI28tWDp9SohAfa1pSk64c7jGPGzhDYHkrGftqal9478kHk3ZCx4
mDjxsY/II1o5FOr7WaFGQ5j2ZAjklUwZrgf4oTd8MEJNI3I2UV/C+OTJaWo8R0xBd2mhwe5GCfLa
PJofrkeA8YoopCpJ4Uu/g9JOFgvqFRrxwaZWm4gPNq2IpmYW+WpASr5OdzYKu0ZAz4xDaZE4U9VD
RO11rE/mLemadzd91OY4gR9483SprmbIfGAeiDiRDXsEMpwfID8RRWhq45WO1DXbLSbLumB2u52i
4tlKoH68LOCr3GOxZsiV/aBohun6JnoftDHx2Tn6e4rCt+c5viE3ODADj5ZOdr4YehvihLL1cg0P
pM/AXJns+9K5rhShM00N8uzqSGp8WtHKFqynB4sHDmkJx7kp1HDEDGebvZ5rfJb5p4Y13EFBSapn
qudUbCggKzHIKPyGQjdx20ZLor9Qe5K/GuZIAPJzH9AgQ198p2BFYmQLSrpzqUA6ykgrroKkEAEh
wt0AO70Z1+3qqvxK2mKqFie1bjfEyh2HBYsO8eKSPtHldxRxQ3YuVlSDMpJw+5oWRKPrH6q6WaL9
Inx7esgSbqgMuzDUjkhJLF8VNyanNigokSA+Q22eFDdHYaw3+GDXH+1ArC4+iw71/UH/eeSeOD1x
TJ8Xyg1NnGvkWt4cF3UF/EJ7t40nL0NSeA/sHrZ6DIJj3+uVxTYD1HN+qeQ6MmAdaSu2Z4xMcV0z
pnsU2NVhNU3yz/Vy8yjf7BVORTd6JGCSHa4zpovX6Kux78sHQ/WcVDWozW+4JVnFJl7FAGTs8iGA
f8HAjbUfZZVg4Yxldh9VumyHCMXokizX15Aj1J8w66T4Qyuscn5pdA0i2p9h+qD+qRNXyYyrTyl0
/MbhQj+inhYiRfGB3F5OfTaiVjV3fw8xJSbOjMA+RbGHdcQdBs4irOF9baF4igKTUU+oQFNcJjul
WWwsGyLFLE6rbtFz5wWTVqm8ZYYugm6NOhH5lCTYfftnTKsx4L8XGQog3O7xDtAXRAdO9FwvpgyN
Ou2GC72zPmGYcHPePDcXc9ugS2ZgHGF4V8s3VpNrIntQ7Yp24IVN16uQHNM9AX4ujXQGHal2gAS4
x+TEJjNiGjW5bjgTlY59BVBsQ6U6ntO3IQcacaISnE3+UFE1C7yKH4UDfzRpZnJVwo9PsAmE64eW
J/ZUouKLTleNYMZtOZPKAW7CD+lmZzOAdLCt0XbOzuQ2mYXlWtPEZG/hIFZZBpgDBk4cjeW1Yp9S
jj3k4PaGVwTqehSQTZVaoWMYO+IY7Myzc0IbESEEalXeKrCNoxgmwpoCmUIDduZ2gjp3HnfhYlJy
wdP/VvhKuA0WRgnWJFC2JZ8juV74M5tQVs6Df71V4cnt8ZkHA5PGaR+qKSFSNr6g68zFRSiKAs8v
pbI4brM2SEptrEOEpt7/Yk8gLOeTuRNCmxyc9/8vnhTWvRkHucceuWtTtkVuGOaN1OTuRWKvSi3F
WoDeN0Nsz+5QSsbNkwkl+EtOFp7sySmxvJLMrtvfiL2jPaDenLkyP3hRKyd+JyHSLVuZpwqFhMYe
p43hHEijtlsUjgSFEU8W8J258Fdcn2+iytgq/07XHkye/n8Pzn0SZkInrPm6+LxFgAo6TTdnRrND
NlLgruC8aPdTIxa+8o1NhQRG/NR1yljcMmib4MA92/nGAQ7xAOwXK8f57Q1DNNsz58Z++Xw6EAaK
Xqg7dGhsvQ8AMwvZOvaFV0jQfWow1fwLXLCvgPCwOz2kVVSOFBPHgjpFUZ3cb+b7p2/pfzebRVLG
dR2t3tT8IguuKzbnudu+m4FxbDhV3DVMZxB9ACwKlyPrCwkxZMyYmvQSN4+GlQ/bChjhBuI6p2xR
AcOyJc7PyjcJIcn8rDkaQyzeDp37XVBPDqg6WPdTNNddnhZY/ysVrtdnyAmFKMUYBI7hkKh/ZBUb
6Y13Sh7U9JkSMJOJu09ovA0S/poBzJpTQrvvw9YQu9gNGAz+iNp+7QupehVJjHSonhWtwgzoNnwn
DXlI9SqXAwoV9q4wqFx/HKGt4ZuNPku+MxX7zXThv9kEvzDv/aA0C3eE+tTyqaIY88ngrISQ7un0
fxVGddjxZ9gVRllEOhYRS3+dQxXVHELchiexN45CNTcuhupLADEnM694xHELH7kcVMnk/36H1UIt
tiZF/ClZhi7z1Ka7BmP4URl+u/nEVFZ7/IaajLQFvdbxu1K80IJDV8FgUA64uVsoMfZDdNvOim5s
nF1730tjiK1plhCxODSd1cBvlAw8zJrmtwN6VQXFCiKOwuH8MoinGRFKLydD/KlgBBccyA4q9z1f
zY7gDjqXE//DkovyRoDT18tOIQmtQ1XNrYwZDchufKJcOPnLKcf/iHJ6PurZbctjcpFTKYcoHjwl
ue/72zSabXCMmTd7DugVnR0ke4ujeYLXKQboTCJHf/bU56FylWCX41iui/esClRZncszHEj0T9wJ
HRSGX7/+YVwm3QgRvtofTR3Bd11OSKQa0ZyETlr4fWJyxRKDFQDo5+wRC27EwR2FKLzCzzi/Wu7x
kmzwtOD6b/hzBnhDUN1EtQZkop6ogobO6OhGx+E7Eke7lc3jwkweqxNBYwAvmXqMMFCffwd8+JsP
MuEBKQQeSZPIuEPd1iUkkAsQMWAfiJZ4Q3Op+NaM8s1lOUtcwylR+r0E07bQmM5VoPhmWvW3aNaJ
Wnv2cYXM3LU4LoqC9YN4n4KteLPNYomP4DTLsaKqXlCJ7RW5arMgRWTRy9eaOFgXfsK6ydG0QUpT
BQ5wIOmxtEkb84Ai8RsFuEj0WsXKNLxwuOo3fTAWm2kBO39+FxfpjsMAjz4Aatt1MGs7yKxtp7o/
dZpfdToaYoxnh1xlD6c7ig4vA9KTId0nQRYMJX1Eb1is6JZqPoJSfdKOwq+tqsL+7pJIBygff9GP
EhW4VeymJeqKAMXvCQEEvthtDHniU2BoK+Valh2U07TPpHlvdk63FAHP8erAV2gjtNOYFnjdePo4
QwsVNzsA4TdB5HP213je7JghgiSj8RW67JWwbd5RxJDftGHj4wH/qggPP5Pt8yq/fw3FxRJ86T7g
R7AjpgqTV/CA6Zhym7cK2M5Q88NYebJfb0fJPSJdVl1UIHSTtTTC1AWYKbIvVp4GXuJnT6u/tJev
sgTCTm3SGpHsHCEfzxdAknJ/v1Upafl+T/jcW+/NESWQg+9WP0WHZlMxPgZEo1EfKAAhDvVLRIbo
9QVB8vZFuHI4OT70qquY51ny6ruLaV3H6Ibtizegww+4pOytHBnP8lVmITolnpz/RFM7uKHfJiuR
NU0vPkDL7phnjY2Y3AGSvRMhW07fGCSaWi/m6Pf7nWwJscUzEwacqSUmrDOXisuEBjmyYgr3oTYx
JMjIMFgrUMpT/DQEoBx5ahQ6YsvqKD7YQBf0GUV7HLyE7O+O0dAWUzfbJ1Fnp75HjIpLeO/weUmR
Mckh2Bvr+r94nZl+qI5bBePxg6vJfdXPls2N3Wv7/pQNAIn5eADGlWtYF/qy3mBCKNamEJcI8CkZ
YO6I88tBXWnWxNIRxH/sRiEPhCb46S0ILXEdQVwnPf0ZvLtN4e7rFIqYwEp9ih+BP/0PcT6wDcEP
wll0YfjUzi0MGcWlXXZiin0ZhWl4o4e/DMsM6+rclDmrBtIayWq1Qpd+rpCuZgAbdFlDwawqJFrE
lwIIKiTq4I3nLaTZ4YyIHpyJp8AZa6cZ2E2Uzt0o5XKYhKEei+kUnRRHLAAC0HWNq7vkFxdAAoiW
+SCuoE7GNJTro/qn150H08edzy/Iz5ULf07jpjabq6IhZniZrD4jfcRtrsP0LI7i8xWdsKcHkxf2
9DnG0tUJSd2T52YorSW4fnqY4mTgpCaQyeKIWNycRUQp9QfgLfECEOvXO7hccBmsv03bk1dD7uPZ
quE70YSI2cRPLdhz+fdMAOUALh3FJ5lO2g0wzagUqYVJjMees3tvERDA/zPM6hKaYIqW0kDqArji
PYvBtU61J7D7wRn3AZktJ5pC2/EKF8RYLfPTyGTDIpyImys3+KOEmo6gELbIjndcNupvrunWbN8H
ST4nD8e1nY/Lhl9iq8B3UlcOLIO17RyV7pJsyQfCDArfaywaHBy16vppAf4yUyC7jASDHXhvDo47
u9vm+BjPVbRcBd1e7L05hgd2i66VS7g22nzHpz+XrWpQGNlwjI5fiCUWr1wHZcBwLvvVVeuheS81
mOe+vHxBL875fUVQ8GIvSfvMWVjnP744xYVLjCmhiOpBsxgFIdZtcSnQoSSaRX6TZwM/sdjcCQBL
m33pgTKGi3Dnl0APwj0Q5ZjvX2ew6dorxBfOEMYh6+A/gsBqgOukbTIFxpqmnCRLjhf6AzVpPqFM
QL1jp0HXJ/bMlQNwezf/Q0Dm6MRppqSP9h8uGHHMrWBiPX8/mt9EB7QXEzD7xEED1SHpOqsWC3sw
iY09M61aSi/GcR286h1FdYv+QLNvbikq9qxYSeNifBRHRNzRE6KLla1kQcs+JIp0HA6/Sxo/ichL
3HbpVyqsL86p2NhdVNVoW4PTgmMUdfo5J/z6+uRiatfiJOnumUJObHcUmakmIIyTb7snLkTLpdsc
Cju4nAUuls8TDPFOvDXY8/zSErsU8XHtCE7sIogRvSd5ZnAlRFnM8awr5GrLQBlMHKEgZMcW8lmH
snPiDyqPtfIkkE9moBV/b7nGORUI17+GhhTTAd236gWPSIipdwdks0/opTC0lC10k4Z/d6tEtn79
tKAIBumwYjgwrDwotRikV7/dsNb5A8nO2Iv+K1khos5spU63TCbhHbRkQ7xbTq8wtIPzTQe6tFxk
Yj7v3E1sOYYZxTyUv5RTmIXpoR0zSVBYHb3n1/Z/9qoficXSeNaWoa6UwOTPSVb2TEEQ0Dm677jh
nH8NS+GnQSDh6d1I5hZPtmLPziVyqeE7ytTNmzi70FMf9rFm93IMDNkU2rr551asiyvyvFJ9NXWB
apkRdr75lhsCh5PAw/g7hZlKHkvYJ7Ymr5oAvD0dC5w7wL13QenZ7mL9gHY5i3BppH/RBnFledyN
5OdakJO0/ZinuDbN6WG+GvDzQhhgpwaOMksyfqlSuwE/yAhT2rAqXfGiGvAcbRfJG+5r0dcxKvMY
nVSYJtz9oDcPePOahImZcf/WKhKIfQ4hXJsQDXUVGGG3LqMK/6HOg8906iBUyl89jgAObXDSEpoi
T41hQ63JXcKJ6GCrbNLUKhkFVbIQRcWR02NAnL8/lLMAHP5vHHDMigOHmtRmhuXIdjhQdaKt5TXR
MWDefabeFbrMfKLcCy0Pb7otkgoEkTEK2Uj2gtERnpLRoGqiNJQLKr59tNAVA//ods10QQ4viZA9
kFq5TzlyNEXJJAa1UDIXMpBkK23oH1OrDE9QD6Ci+s/CcB+2ATKIEkz0H8hFIVEJekmuXictlRNZ
5/QNGyLVyGF6c+Tzrf543L6jw1Z4X4u9Fj7UHByjH9Njrf80M97okpnwzhnPPoxAPTocyS7luwIW
x0SIQyF+oTzBggdjftR485LyIdcxSTAVpfglaDcmYQKK57JQprpHUIwuNRDzVjIWcyaJ8fdAzSit
AxgJNQUCLAbvZJACI9FjTaxpVar3BIIhxgs1Dr3M4iCJD/2Uav3EWKLXFq9c4drYbeDEZJC+oTh9
deS0t1sq9TJQ8VPAx4bdtZri0thlU4jtdE9gSo3lYcc7yAUDcJnu2StM9nvUZbP1EWFrjwYuWiRv
4ogZyTtfp93pZ0nwK+N0n9DV9qwyXRRah70Dc5KSYT/ClyYC40/K3KE7ZavSknlm8mvT7ckxT/Bn
+hAAu0HyKt8iEyY1JMvrZGXWVKhibGzjIpsiqilTjL8OzgPeYZP3qhrhnoWM5NMne+xh8mm9x6OZ
r5K2pDOR7qWDK4VnEZ30OcDUDIccVHfHCunsFX8UgMSJrPn8buojxm5W+EOxNmMUEDCKehcuTFFR
2GNZZo1q3mfK8QHOD4IUtHAkfTBT5QYmB/kgPD9Erq/xOLe8sLOgfHov+BlxGmYh6LN3mMnuSsC9
xOtVwODptpnZ/T1ACDF1pIGyJpn/xG8OkiOFNbncx97xBajKCcZTzjKrbCUkK7n2UJovXmDTOfFj
sj5ZiI8UgX0BAfhM97zrnT2qkZNZXsWiZ7Xz1dxTP4OckRArxmNAFgsSUyQDVBb3/z3jhWtQEHKm
hMxoINe5z2FKdqzioNjPsKYLEdgQAyTChPNcPUOstC6CbcrS+3QanJlJd68YYXU9ogPRki2E1bpM
8N4mOnlRuIkqFGCrQIxRt29mH7YmEpOknT8+ooU67wl3E0P9eb5So7TSajzgCilZsRn/x6Do50Vc
LwKW0O1IbtnUPxriVb6ETNzEmc/JShyB1Z7ZU8A0XccIMUuwXeDGOql8UvW5xRNYMHDG5X2SMikZ
Mg+sbgBK/Sc7lywoRWr8Mutq63c0k61dVb2SxlUmWHiWlk4EmJJk8mnAlTgO5QYF9Zzvxi1m5IIu
DCa3PFhnGlgvanbw5xdPBsCt+yKHaFMgtDLSsSorBHNTCynQvv3cXoNQ2uASQuNLC3ORTadRqwpq
ivwbNftxu4i+JXQm4T6/cB548nSkJhP2tNbDOSIKqRfa9nXYej+sl4/9AuMmByCeRPNjK2Ev652T
NN3XSDRODHkHJWE3Im3hBTQ3js0GPEZKmew1v3BdWW6rbY8jopn+Rc66tIuQjm7/yRHhY8VDYhHL
ThXSMb+x+5nRPebMxZi70VV8BWOCb+58gfTUZiT9HE4BVX7FrXJhAsO3TBGi6fDZsVBNKFPD6p8z
HXz+VNTdSV7MqZO73I/1VFRQmx3hpYpK/8xOsH3GHiPSnm2Kl4O2eH7EhNx2aXWSB8hn2ePBaXYr
m164dXffs7tsMTra/d6iH2MbXaF7oMvQt2mnsyvznFn/k+hCLou7PWBSuvKmaMXt1RmwSAR17i0U
39KEls1pbFE+Zec/jBTCAV8HC0891MFLtGCbMzTKymMgAo9vqjzN2WPV/i+vx27TR6Pqv4tYe2vJ
HPdEcmIsE6BfDoJ/THQl07HpZsnvLdre47vSSEqy3dyTzUn3SkK+oGyi1261ogrbwCyW8hET6jMH
uLa+uLEpLIXeCIXj+7+1Z7Ew0ia/r1V8Qo3mn8S9oA/lLLrVwDHmcfVmjK5Xaglm4y6F4c81nOK5
xyF3to/QWFnJ8/PxHSibxD8NbC+jws3O13HvF7Kx5mNGcUqDRoaH3L8vmIk3M2h3+3ue8I4C+lJa
lgu6r0ZHbFZprCcr6ItcQ82tpwBuozvErKTgN0gJoAcJUrSyB5yMTRbtj2YSiXGcj0lgy/Hzgxsz
rsfwFX4AA4U4GZnlBI6NAN4/Yuaj40tGClNM4cg3yyOrWRayL3QKpdzViBDbUiOg8QEjUiyEns2h
3tYnoT3wL3vG5Uoua4a/6Pip/JMDrD9hEz2J9HpGwoUHL7LNYKRgX95IPPb2JzhFmXAlIbaRL5qJ
RwVa/lmatr3W6ySiPdy0yREsz1fXVS7bNL8cu2DlVmWVvTQIC2yQjhArODv9eWGog13EEkC4CaUX
d2Ei7lcaEpGkopTzp4XAy6w6NyhfUFSWlPoHCGNoGF5ZjoDOpFtiL/y/9CcAFxdP7OfEAAAdqY64
HH5T3YLkiKm/r2NkVmXDu21W4JCPDr8nq1Ij6lz3JtQRjNh9CS9dIypgWAdtSPjoiFmJ2la/IkoZ
KA6EELJqknPNB2wvDm/N/BEShR662KPb1loi1KjeJ9mHTj96xOkqS/7ImEiOjU+KH0lY9qt/i44B
asDbZo62j3GYbGd37YyNOqq2vAM0cnMK1mqFP1N2KCDfR/k5LbcZjAiWH418j/W+01BKR6G4o3qM
HXEGMjxw6nH1cb70mQPhb9ZOfLS0jrkZz3yjLjq/Edy85/CxJiPxV/DtrqamEItJ6wTEl2czOM3p
AyVviuyvmokE1Y/CF5MZD+TJEVzfLC00cU8Kz5vXQGYYr6TcHCI5G6KXSGqHMgDYwWUIbZ76HiK/
BFlWHh0D1BuHQ+AOObx593QyTr1hvrHi3EnubGvEpDU8ogAc3WOlaX4YS2d8ZDE/KEyqea/IBy2G
yI2nV9MdYZ+/fRXNT7MABsqlpU7JfPCNMKrLttFC8kbY1K4lYu8cwJ1jEvEk18dxwWovtJ++zQFN
qPI3ziSy3175561PsV3eKF4PTkvHvNop5e0yOnyAtdIVN2iasX8uGpzEVKDMY0SNveHcnCpkYW4T
YNSFHuW+j1cFNt5B8+SHlSeXEvPKLRrjwUtHb2pISTuDJOnowMIkU6BGtDa32UFtNopJXeThsMkR
SVu+hJW9ij+qeSQW/mtulG3N7n0D3yeHkPMaIQxpXY2HzDSp0PbIcdmMRyxk0pCb9GCd6GhIqZCP
78dKMsFK6FzKySw6u2+Axdc8ac3H+V4uyMe78Zmryo+H5nGAbDxvIiz/68zkJMyXCi2wYIYUZDSl
n+VfFFdtwvSHGQD0gvRrUkgQdMhIjPBxjEv4/CbdyUXS6RvqfG8HowifqAh55f5YdYN0zt/1PoYq
3FCJzBMb3/EuamQ4mMxloMC35bct3V/cqgrjA7DfbPrcB7rfQnVA8XbK+48Gi4qK/Fg3IGuPUiGy
BV79+1XoT8mJ8Dm0raLZ7u9lazmNZw8uYTioEOKKN/Vd4+OMmOlws6fsd7R7vSxF140I1nZncvfh
ZlU3gcePYusgOQqsZ3TkOJ5sN4169JuS0lSYYiDHeIipOfNz9tWkiTIHp7l+3z/cZp2nH4qEo7o/
bsBz0nWVHDLg3+jfrVZEDIj97ZlMYJyn4XCJLhhK3BxJBN/3+DtaTZ/w7mqsOhbtcBFGk9YWheZO
j9JPWLcudbQpxXQGRwDI2TCE77jO+dX++Dius6fR4C/+ORne4vD1tT/eGYYdgc8hBtqK740JIrfD
mNbKlJzxwu3/QgBVUI92KjMjph3nMnAet8nYDm8s8xHFS8hlaSzQAw8LmG0AAMiHKhvDepKbKuSc
HJSTWSyXl3lCBjbLb8q6Vx8+aeHtwaIhPnUhtb6K2Nsf66LlO8sHOdBOOVw7m0JxHKYXJOTnYWaP
KdYUvntSHFlTvaAMzGMSwhr6ONXvYaW0UvqeZ0b5PkAaJxxw2XMx55qxYdyQ7h8TepnaB+VWYkXl
oWqb2R92iiTbxJGT+d0CRmQWnxDDvh3SXZxr8u8o45hLQnXrCLNZ5fH3kI5/++tM47CmkAgJ2Utw
RDan7A99mAwtOABINkjMpgXu95i9QbeeM+0piuREOx9N/SaK0rujDCD/nciWLwt0gY+FxWt6vHe2
GX9wWcFfMs5wA8SSpEyQUIqNnJU7DkTapW4kYva3m2WLI0ur8NznzHS8jmfWhCqZqmwD5PtCkJ38
lFbn/NMO6wZMsL45VfKbE6bIuO0B5dgv84txNliJXUXXTN5tkXy72P0LgiwVlIyGdPJ0kS/c+L6N
86sW0HdKGV2XVijFxtodUGolaxA0c7/C9uYdVM0nOsl6rHoHsHNW6+e9qNGiExD6AKDTuMfcCyAG
Ckrs6pshVTQmrVK2eB0eUoNbNncuZ2WFM/m+XfifHqXzXT2FafhZkNgchz972Wgd0mlD7EG/AQo2
q9d3zqxmOTKQ7mtNKMH9vYRHK//UZ926nZ6Lvb6eVf+PpvW4yRUxVrtSSE8cwp1VPJFriApkunhN
pb9F00WlkWBoPTVfy0+KO5+urOe8WBrTHP2zmIwWj6CzgimvarUb8uy8qs70xc4tpDkbwru2aqF5
4tIejKjCHHk7wOLeSPrfKA8QZKmeJBXSCHPLyBqKXu/Y/yGcAb1wMmRfDTYp0y3Jk5JCgBEq1LLD
UU2AWbYgVq6eOvC7LYkifEVHVsX10JO5fklyjvFGLPc1wUXT7isTh+P4Ok4eSPrgf/4LXggLn0Oo
cY2LGXus7IiplCa8QOpPGIAcWV/HSzOhpMax7ZhA+ugJnaRxdO6YCzWCuvemLvcxHkiYOHUvxLer
K3nXZCgMoXLq32YkGnE0ZY7QOz/jUYhmtMiXWrASjvIZnD6AInKkzrfdTeqcpzSTG2wdhJKEYzuT
5VM/bjhEbRUl5z0KJBXFWBn0tLK0PpvcyB2eKk1J4hV0Ghylbps3ulPLUo3b63a1t4sn4hKopPKQ
pmjo3qA6Fmnwy2YjHWmPVsfWFtivy024NayRCK+F3TxqTIBsj3IfaTSpL7pE7/iVjDc6obvRvOOt
bEwIVCwvpezd7CndWEeWadH1V+B7RDRQNJUzbg3kr8nyS0MRTBYU8bCnNbIBa8bBzlsWBJQ4SRVT
sOb4/eWYLncxkOCQR5EI/xjrvVrk0fIegYCX48C/HBoTfOBw4PZB943pFUOLGpMscZsSCbeD2OzR
a83nXfr0v/eLHiBUqhGWym1OSLrzi3NLmOLiesMhN94TBZpq8FnWRUUuQenD+RLt/xh3fIFEeNiX
0BxklKzHcjAzr0Vd9WOENzZUPdFwbElEXXUay9dFaupCnJuGAEsMfCUW1WNE9R/efoZj1HLDFalu
/0JxwEcI8u95Di9AbQUhiC8dLYbTMv3QJLgFuDooeLnJpxECBDlCQ0++hjQMyz3KOMzJG22k2UiU
c1iM3MWD0h6A6Y6sUcspl3xa4X+fRdlYph8B4AvXv1hYnzyxM15WddOW/gHyE27el/KAgc4BmUdI
Slkuy/3Zya98oP4eWNiNvAqV6B6+E0O4oRoVpDhNVWfJv2duh2b06zc4fSwcY1tM9UUR853HyTw3
IwJ0ajtKKihaFw9KnBUYcI9U7ts3n96ktIkRP4ER1+XnnUvLphZ6zVUZYGgNNJAIA/O2VYUc6t9x
pVnyFxhHF/KE+kVkk7oZmIsi2HrlNpduPLmIph+6pGxyIDKyvopBqTV6O3wy3gyLTgeFn6ymU67+
D1CVTEPfkjM6d5jrIEQIJcaoyB+jTSfc5dRNDBkxfvs2dAlbPe2czTG1CrRvDk4pr1mQsCujsQ2j
4sETG3QxEh38jV1CUZp4ga6PTqHD6iV3wJr5WHisKbIKMfHwubKVrlbcUtDBTPk7UA4V5x/AhQUa
1Y2+rydh5czobrKh9OXx6J52LaO9to30efpuWtc9Es9/4aAZ71GhxbcVfo+RLi1LgOJdrjcK1We9
kOoHJ7U18hfPpXDHrGgV6hJpT7RzEx9ENoBqTekdNxzA7P8y/+D21bk+dcshU+D1b3CcDX9w944H
kv/6EyP8VVDkJYY9eDrApXSZLo3xrV9DED1QWbP+UsPbSk9w8bRx2J20QcjacpKDryO2vEa+zOHJ
/vNEu8S1Gm3cnsUOjOEFEuE1VtlmDqDpuugqtVjzcS/RCAuGofksaw6WBPwL21/oAZ0lUK/LUWHG
Gos8ssTa4us4gKVwH6/cNch1Km5pLlRJOgxonX4QhyGcDmOwN53KJJO/xYU/6h4panyxQTz4ZAbY
Uf/Eh3TNP0HWnFXcxVW3joymX7bPh1g3+O4ndBvJQ80nEO7BtQCo8+w9++AfHmTiEceKxhcDCOCn
TUNQx4iVJ6XjYP4jKhI6EM9OZshg77WiQb1TJoN5uUzi8wvh2k4QCxFnUxXkG5N2Ei3OeXmYX3Yn
1Cn3XGiA7KY4ccpNfD3IvTRr/HHqbGnyN1Lwpewvw/U98nBs10ealWKs175kUp7yECpbqxfdHurW
YCdSKGi6JxtZ1nhieGXk5DLtCnLXFUamN8Qt5kNjDylUGaiFbc6W45TkTH/pYQEg2BFtqkIKgemp
aVnFpyawQFARnx7BpvDF3YbLoLStoVgOWLfy4YF24ea7jShf5ftizpjpfvpSkROqKpFtnR9Ls9PE
vpUNTjStaCNgDl/4s5G6MK3moM0Imi4r5zSZoaO57jvYHzMK6MueW8iVGdlbYNWJrQ7HWzl1gbPT
AgnS5asw/Q13Ar9BDpEhaBgEMtwthsiOxZH1Z0c3Q0FklX8/khQQs6VFr1FmXgEXiaUa2yj1WUQq
dTkncwfDITejCwy665k0fjd2rPxDEP3wnDckHGyWVcQLDv0OkvggMEHZXSqSozDe5gUJ087gg3CB
loNtc9Fk3KjkR6GYg3IOv1Zb9LXSdExBi31gboWnx5PNGosaz+CyIYTpc4kkd1TakImOZeKxM2Jw
sNGqN9BAsRXREMRZbIUJy7jUBVFLIdZI2zG+YOUDVz6Vyc2PzJIHzS8mQHNieKZd6gXpFvm8TOTd
znEOn/jepFlmQQ6TFcHbPI3G5vDKrql67FXbV8x1QX+6GlQcBQRsDk3oiacdsXVp+1SZCskRLSmr
FENv8XVzuyeE+6jjNttVu9TYMZbEJFZqrIj4uhmj6i3iLuLDF+KdxuOBvljeMs0I+XLsSKVx519/
M8Snw16xS2t0xZx1lOnVv+seM6Xvo0XE0VrH6n80EdGTvPGzv+QXrf3ZZls2MG23KCO+PW3cRn8J
jkdq9sH5n4/UWh5LmrcsCMAeXnAhW4Ks5nE6CniLZljfc7PtVbhbH1B3j9LOTA/MUgNVU97TbOCM
sMR97XHO7M+EGn9+7t/+b+lYzUS844wpidKjF0mYvGm4M7mxdSNTxoLDMAcC0trg0Cf+mUj8jIQv
gSLTT/nd6/gUA1VHrMjmm8LjpZ7+RqnSB/8DB0cR3FJ0kkd0qTwg9GE2r24y2iZwKmh5JaDrYjXR
01QDeLx/s1VnPpsb5wSEP8N/Lxf32E3zPE8cVqSyY63J0ZLsN+RCEtARtfdfo6MNECwJRaMTCQ0r
nfUQgzaDEzsScoWQXxb9NOJh5eb/fcooVZHdEiOtKfOgb2JTel0O5IjQYjs4Qd5K6qTS35zUJQuc
0HaZfDsKaLTXbFXypUxq4SpvAkrtvjtYx2vyoFndiEnUpU2wg9cMLiG+zHPGw6xGVHAVQHk05KMh
1qqQVUHf58wwIdx8BY0jnMsPzbTzU3vJEqnEBnofPvCNgWEUAyAdQdA813mY9ZqBFFUzytccD9bw
5fTJ2Qgk+f1EysTGahF4DLLcHqwE8QtXybgcq/kdbMCDhjxvoE5OJkg6BcqvrnZS9+DxaeAFZ0Y5
qao3u/7TPsrSJoJxjkE8pO9lWk0EE2ceSjxtlnwExh4xLEwLkHDaI5qEQ8ZCjir9veTG2ALKqRSt
53NT+M2H1CZohUWnQqMu0A2yQ66R6g/uoi/PEXyCbPrF0L3gxCfMKNIdVjAwqym9MzXVmlaqHYGR
oQx9mm7eM+xbHf3sIxP9BbGELtQw2iq4/NpZF1ZFFqG8Ric9dS7SC6IVeL3Yz9YjZVFnW1S5fPk5
To1tuuCcZnK/72siV1smUj2v0UgTxkOyy2wg/TckflkP4cbFV3OZuG9ma0A3+08FrV4acLfQg8+i
2CN7xDTb9BSqDKGybD/foTrstYPisJurECXvyFoyayG4OcyNhlpHn0R3wXjwKOgVGIZmV7Qiw/gZ
OE9I7QU/PWPoFfE/ot/rXI3HpC7840d91o/32qOhYQ0LHnq428MKt1V4PmIHN7rANbzL7LRIL7Lx
udfbk9nt0sM815mf6iKUw4HeaVNVI5KBdfo4jeAkS5X43utbyQXB16NHfzrEkRmuSM7tpaHpGIZN
YKfTytcRUvPQtKaxVgDaW1gBB8MoFlKKy76CjvDiUT1cS0h9zJC3NPa8N1oIWi3Hs0yUAvRozM6U
9A8PFQnriMAxMPzmXIQGPMLVBPuh4DeiCP0ZjjNJhfn8VEHG6c5ljXn3Ag5TRaLPtwdYM5T649l2
7lvjua6oicVbfo5NIplobSO/s+6dw5vqE9hoHmB1OzudVWxRkZ4IliCC21EbbuNV4g4WWzolRtvt
INiCQWj3NQveLFXAi4nvjknCZmeWr3s7JI1g7igJyklR+k5UdikPVejGF99rIzNoD6MVXOPAeMIc
feIxy4qLlbz9at+kUeoRgtAXlj1rvzuxjQnlPnJrOIMaUh/3ZQyZUCEIGdKJvYsjIh8WOMZYSrEy
fA13PmnDGEMlPDihj7N9U4JVKxSX5/K9/A6Cd+tYTNW2+qhdqfqjgGpseTzQxByFNNHdp2iKvIev
3M1Gj02PIgH4cS9MuCSI4h/Wxocgho3iT7TCCgeVg1o7KHWLLB699CDSMxEhCvuwWITiwSEvgWeZ
DKj4xR3zbYTmJwB9GHQByh8q6+yIDU2h03YGtGnpjIzNXXgKoy+vq9j46c5gkeCFJSvLzxVbki5s
VgepBJr38hfNW/mUDhVK2jTFA8AfyG6gXPryMTYKZysHVFCDPs3dfgGvp6rZApksmVRbjclhDfcv
ki+fTy8i8bT3MPeRG4DeMH+06VA65HW/8tbUvgVF7W8DcFlANOBSYl7uqptikuMtpDau3B3W/NaO
aznwycWA+aDp0E4ar6d3HkheCNYOJqIzy5/ADDjYg2HzgDths6ryHkskHeyijPezemrn3M3kabsU
94ULE7+KFxmGc6Q4oRjSmtgk5qAFjvUV3C1NyvG/VsQAhlskchddBa8v856DBC761tac3egmN5aS
dHp0CTyHStWCbksXlO1I3uxbUFpiCaL4SMbrKN9MBnYg8CYAm/FKcjbdSkpabulOU2IGwTIMKva2
GJyZY6acNCxGOD1czgVowV06VuEVKgip2BqGYP/cvg0JCqaDms7/PDSqpeUvx6naJmcfwi76bjR7
VF+Y2Ku6apOl/ijzeGIrmvlyD7KOWeTwYH1DCzluHYt1nRv8pOMW/d/iK0lIFkUKYJ8B1BH/JQyv
0Ub8OFQ3g8rccbTiBKsPvdbTJHUPQJJWzepjWwprlS88Pblq63pHaHlYi1n32DrhgNJTnZHbV8V6
+SsUGlRvw2sCYN9uqgk0dTg8U/2YvVD2Km6V/QFxYlBffaWGF1YdD9B/XUp6aic3+qQwPJB9jN9W
42yNRDUqbpz5vcH5njMBz4a0StHnQGKVhPg6lL02jD2WbhUs+RjCr7meLCzTx84aGLUiX4aS+if6
sKmkncSD/uKSjA5KQGFdr3Tk4pqZeu3ZaZLrUWQcJyoreI9bQNKkcRVjnL2DnY1V9h+9LDWIbWxJ
W484Sn/Bh4oEMJi1X6IdmhgsiTiNzjMoOF5GwBba9C/y9EYVYCOLR+pOIiDTqn2JHCSFX+m1QS/W
XaxrijNk4IQp6ynwTHmVUSFFy8fc7djweHyLnWNmqEZ4eEYhjz9PxIhBkHr9aiyR7ZxlaBAzJQ4Q
k/SSNYsn70ySFFhqFigQ1M6Sb9WRXpvWUwqNTU2pCKQOBQ7mQH6HueO8m4dmjVeYGedWTfD7LddQ
IG7xkb6q+Dj7WKiWejU4InY0Y+RCnJ8mHyWY68aY0sLt9Ss1oWnU0LjGWBjWxYMeUFp0suqGUMOX
ZE3pKkUuyvRmUqXmLmTpps4EX5WrY/a/J06g6moLV4iNpN6xJxufI6XFDYLFq9S2LjAoN106LqpD
D5h005Hps4NaXLKUY0jm64uMxdqsAzcnyRtcPS+gcbEXh0P86XcX3NX0eua+BHwdFiWj4A+XWuxJ
ZyWsTQVpQNh7txsAXALy9s7tWX4F9bn3QpjzOHnznzcySafWi4j8gMKsDO8asDlApiUAn+4iq7Hz
4qEn6fC4IslSAKtMGDR/Yg2RTQU8VLDbEUUqlAgsUUojO9YF5/qs0twdIBKuMT0tIZlKSepkNJDw
/hW5OqZe3PE0e51bP67aftwsGMtD+ZC6UVsB2sxrgC3BMxlEDnGnCeyzgKr09URL6DtDaFBjQllx
F/t5KcnNG5TZAQ8I8EovgVXlSpuCwbk6/Ixs8mJpoYJF3NGHtkTDJUadriy8/Yt1qkepDZ612bGr
soqUN4QVgu+TaydS/K6eOFiEgz2VhEgMnMp1lQwmXCKqzu8wh/O6+35SR9R0W3lNiG6bV15WikJz
UPPfZVar+6M0Bes7QsNUoTzPJizaoFtWi3HffQQbqRLrSzlx4WSSY+rZPGo/zo7zzJacG9kXdJmC
yZ67nKjD0SF3hNrElewS7VShRq+X58bMqcp36rmePAXJF90lAPjDq7fj7a8SjU1QRWcsB+D81bdl
UllIF/NaNLUnkj3i+ZWVJun5XG6V/qRhxJYuypliqsce+Jeq3qoZ13bNBUHO66QDoOj/+WzxxG8c
Ok5l67rerhwcotqJd6wd5g3bRbdmrt0VU5hGieXb6KNvrvsNphkylmejpATsptkB3SpYV/WEw3xp
mEUfyk5V1uq5VVgcwpDNNP2K1SKy1Jt72dV5PntWUz7n4kYr8ObZUQwoke/pZ5cfea8MeUvz4GgF
/wHwWN0TWvKfbYFMgx0AzvlWA1FIM5h/qoaHR6psSR/u/a9tmteJOztFHS62HY0qaZFvyT02J/gC
Y5r1YWhUz1bq9OkU45DktqfDPgshUv7bUy80W7++3muJFFKuPqIB8Flni2lwEiT+eKDwsBJ2YNka
/qZmDPF05H68LCQX6cnxfrXrvVhLvxZMi5DS0d31rXDZZRFG0qPPFTaR6yWFLKrPnqKR7RhkBwyT
MsIK23ri8iQc2c1hMtapaapEn4qNCjj8af+XJ2LFLvZ10YVRe0yOoBDLGkf2US+W7krJrBsT7Kdj
wvEE+oviTEyWFTNMTU4yzja9+YmwjRMXqDd4JRbt9kQ7f3M3KrKMzZrPNRj7Zy2QAAq90pSG8vLP
BtUPd084Nr3QpN1uXc2qSgkwqsW+FRfOm11QlytjtjibWoHgyAUh/00cFl+qKd3fpuQjed9A3uis
IzT3Dir+stKWj/UwT+sHUolc8t3Hgd+yEswt9Q6b/4qmoNRe9pISsQy8Td/b1LsbT6dIxZe4SqFV
94KKUeR08yA/1681PddmFnsHHdcDA/AKYMd7VKDdxxrqvn0ec4adhud1/QLTBO/lXoqaUiN7ALZU
NhX60lsXIqmtmXXc4A9MUV8JlI43TQJTFGXqr5piUygVGv11ZbxyYdfqTuR/rXVDtS7wvpHMsd9G
rNCX5cxU6gVbp3vIqaNfOlNybMrkOTRm94Tt3fkqDECcJ9rckHbtaBYdWQi6zA7mOFZyPFbLqvkW
VZMpeNjR5YoAgpnYKaH3mXhizUllQbdR5J+SjopKyUGqavt45tFIec5eGCMTqXZFGMsDgsFEWYQ9
D6a8/i+6J1iyxOwk2E8ol9ONBaiFPDG4cg6bjB1FGH8gzCBVOVhLuZJYJ9Vf5OTO9VAhuHEwwcbQ
QTMnEDvV6haHL2bhl3P+yaV1kBkZvOwNaTHU3Hb/Ho9iG+h+/74V6a1GCzMqmzPYu2jjSyS4XJNk
7bMPi78x1tR22M49HKYj83X6x+QZpKi0L1AwwdxLfRNgxONqyttrcEG69v7k8t9AG59lfVRJ6DRb
CeTcrufi/Np/uWlIDW8cGcX/bfpGyBowxObAieK2Vyurn6l5EiYireKkfSXTU88at/Ci8roNN/ib
A7Cz6+s7z5vUWPMP9NgHcBw31gsRdQ80pN+4Dlf+NxW/SwM8sk6fMV/utUtwUAusGN4xCboxAepj
uxcbrU62/fSMtROPgaBfFMejXQIcTGa5cnvXVasDQZYwu+TktO8kOONMDKTCuqw7I0H2pERl29cV
qgSA/JW9idnye8JmsQQIsG6yyPXYDXzFrMP2ULZVIAqXJq1L6+/P28BNBD9RsZTXrYdIfoDhq9Dc
bpn/JpniqcFG3KZGtBxGOjwZQKBaTGA04t3LumnGckLoNmUI1HWQ57H1jMg8abtPUAwPYMDeSOHq
Eg73JH6infNqkaRij6e1WcQsl6TAw1bsrjTEdNVIX1Qmyw0VqVNtadIuzTnta+iO6hagOi892Dbv
F/tUOuTUULypd6R1yDJukRo0kpALp2dwavsrXNBXb5SIzHa+nhHZHkFEb957r7oXQOG04gnknZr8
2eVIj/MC5tLZ/pwkoksEOazoJ9d/3JYhJVzx8iOvZv8fHdSTb4dSVkMaI3B0McNbJGDx8KChu2nf
OaEXs5oTRgCV6o6GRqWmnCIveB0M2VHlZ3+fxRTxsHP0L6dbMmoIJS3uzM/txOc/zKpme7XLN5vl
/qB6KSf9zA1TjRX6wYluWjY03O08zKR87Vh42lFkRS1RG8zk5vUmF6Z7X+ITnbJmhH0lYUuULZ3G
/2JLoFnmEYrfiwik+6LFzTbRBCjUWd4lPpQhpCPkD2tXR4iKV1nyDmESM6xuwiiqUWvCxf4DO9YC
bd0Tjd9y2AitWkxniRM6BWXRQnn9qm2ORmgXWYCYwlD9ChxGkp5abEvEuW0Gow28pSiQYj+m0ju2
Tm/Hbog1lW90F2iBO1CF8DZyq5IsEl4NwhG42jM+449XCAt77GK0ChHDfpv2Boy4LL0Mds7OQYQA
l0xjx24z6dpSu4QmSAY6M5TnzlcacphFjVCozP5CH0vGoIoqPVSZq1G5J9MFRpFrbUtLn9tVfcEL
jDoCB/1L0QhkiX/vBGT95gph1pb3AQqTE/Rj/hSQKJJQxize6KasoZATTZ0lOpdwuo0LZZRRSG+0
tc9nylg4+9n6kogSAfgPV5CMzw6eqHG4Fg/S0QRVvID21VhJmi11jJUIBuenzoaAdjZIb71WA7ni
C8LayNeHOQB6Lwaf/+JKZFYMIt7+aNRZh8/vEVUD04MTtpN5IVRcjVxEtGEXwGFj07mFVt//BzGF
odGfNmRXCddsgOmHQbdCTrcEusWeoZ/Drw1zwE5UBq/qDCLLs70Xx8XYAOkjj3CTcnoDdWfhNGCw
Zd+ZTrSGug2qNg3jtkxLTLiQHyO+LqXsCEyzOlJjVIkVpt7IouMtfQG9XQ+PFE/TkI16PnYEAxOt
RTP9f1MEEVVzYDFYmCKe03fSci0tSYs+G6aemTHhjVXM8sot57HPs5xL1NTvUJnSjsmWS/aslTtm
TQJH3HU1h3T8bAMWrN0VC9eYfzBHGXx//A0WUFZm1nzVTSFIrgvirOZqAU4phnELhp8VY8LgThf2
LfPTTpSLCx4S+1iYuOWf7uYZy3I7obT6+cq5cbEuUFB+BocIEru2KLZMV18VhKXTmbA+xUn6csJ9
3mQDliTJWdMoAoS6Ayl/gSIwTzINCKqX/4SNLiqfumS7LUVdyDgO7nINDqd6fFKo2K4SIF6fB5/1
xuHw6a1vaV81apYQtz0Fl81hsbFdPmaIhshkakfwHcLi9Oqm4oSjk/idD3jt61hVQ0qo2FPy4JqI
ff50QlpO6rW6G9csCiIzFbBkRwUYMroKyKfmANSPXa/ot31eZTjId3rLSMqRqLV2NjiDPciLp0HS
ePqL9rbJDbmz2delRyy/m50LuSeLjgKpPkdMS07+TTtW0GJtsiMIbbA7lK15Snfr7WDCbSpNmvAr
dpLcf77a1FrlI4xq9EzxTT/2fjlhEBm40JVEJ7AVm8EPDBYZmp5Zfq33Od/7eJRyIQvVLmIhjuk+
jvJ2IUgRpbbOCy3738abs+AIMtyUAdSgN1q2RxL1vFM5h5kAMC0iMLcB4C33cAArTdM3Ka90tAlb
0pSjYFvH38J6sqJc5o0eqSGXD/hWXc5QPqGmQ3VOLoe4nvp/pA8yMnyB2ZRkK0rnBRqxJsLhY4Np
djPGq28uVxRujXnPRP7XZGGCVv8qZeZHPSNthZVQo5Lep3+6WlkKMMDERNkOKZymlEUkjayafR4K
lZNXREa5WITz53H+sPRB06/6g16GoYqyKGExd9xb9AbM+0VZSoeR4fHadqFRgn5x8AFQ06aoXd0e
Nikgj5qIeqmrCGMun0J7VnewLbB8kGOWtnnwnzx7T8pIqn6LzChhqQpofUWkpFafGDEGO/zaaWyr
bFsGcgko0DlJh2L/hdEy8sb4leHv3D7xdsGpr/3Sh8cvmOjuk0pgaUGZzX8nu4hUBdTwoyXo21NC
ggnairCbRGOMSj1Wwsp+adJ6Q+4f+6Q9o/zmu/VzAArVVuJBvXvCs4U8pgsgl3w2FUXlzOpT77zb
Q5xDDcjXafUCt1QbwXzRE47eCTakxm8FdXWHA+xomZ4eZX2yRCj4W4vlDKwGaekVw6Ko2UR6k+RN
1yaXv+o57XloSYa+0QeluTOpPNWzM7+tnb+RBScVvTdb+hXN/wfHUsInXNOJshBssHpA+c4ixhdu
9bC8zrebO5DdK5UvGLrWAgc7l1WThlu7EWMCdmMhmYSbWDRwGmkgLfDUMPvCkA/wN6XsYvNfVBua
be1VQv6NWfYITMfsR/1DvxtvrMYEXF29aLLUgZpNFlD/GDyttw0BkwtslusNTebTx0PxJohOAz+O
Dy8RtQSMnMdZZYmv0RYgCwOXdJImf9BrZwvXUxEGufE/tRAkbfgOpYGBvgSwET165eyLAt4Ds9Z9
nrHET6HFf9b+a6+7fGo2aCV13nX+DTBfNSYCkbkg9nRRegP+XTMngJzNSKgPphzlFcR85NUA/qx0
8JdJBBqzk/u8jC16DybymXIZaG1OjFcoTHnKTaUd3YOgLcdAqpZBdFclmzQvdOyVxJulp2+wenKs
jfoHfrP1KZkgURjTBhERR8y+BFa4tPGtAeD1W9v3owXpmDMrYhkWJhtzrwuLYKhq9R2iNfHqqYiS
xTP+QC8B8Pf3Gr0c5jHEqSfPP3eDJdIC9VVt3FlIHmhbDeOMkQXExzxCdG0rf3GhoAhCgPpDAORW
PNqgChyVwo9CLqsP+Dv87+Y5rMNONHh7jaXTtw2REQsehSFrLVsbeQ1jeWD391TTsP62L/TaNJsp
OtxCOuqW5FKCiM4swtHzekLV3hzAlQDoQsNwa3y5tqo4ZBymir7ysme/bmgbTmLgFv6AfwW4Tq69
c4sK7ziL9U62fw9dOnuy4l05HGmFHHAsU84wCx6q6yfvmpdQR5ji1fT7JOKiA7uIGQnBx3V6IcOP
vdiSyy5+HnCqn6kZ5eN/bQjwVmWcN/uyK26Jr9CTyf46gAlpkKZFUxljWHERfZ09s5UwYKB4k/Qk
+LMxS8k1C2NsjSt8BMR80IdLv+2GMLSM38fe3TDc+A8U2g57SJTsxW2s8mRvkv8jtyWSJ+QYyIRU
mjRnJBV8YpV6MxwhcUx4BfoqrsNmEOtVSJRWjBA7Wf4L1tk2iUKDUQELRsucrzvMiIfQSrNGGZoA
rvL0NcN/DfAFcdJyojZl4rVsU9BdrjfllgCt+msQgYZjxPb++7H41pN/Rsl5+7/lfs01o6+khet/
u8YZRJ9WY/FRUXgixpkNUAtxX22mxmHdNSdqx4zNRStQ6ivUSu6TLUjBTMDgnsUDqb9JH+9qYWk3
tnxEDySyDuzmrpXBvj07r7DqJFv6KV094qqRaUBvQPyrwk+KB0pjhWekMAKNNIq2M5c+vRA077Rw
MvT7GAai+ektkZaCWu3BvasxsUeL9w/ww42DdSXUhzZqeq6VukNSLobrEKcSH1Kqd+Xv7MteCokz
K5woUPjVOYDeF0/q0cplA4x4QJV4dt5pltG/gNyRIGpREItksASy7AXkR12Ez7qmAOCSAkbpK+3h
g36p+aQLajp6dqM0Ph5KLqfpuHXll0tXwv4Ss4rg2MialpZ+BNOPHUuzF8rEzLOlWbokd4LOWny3
54sVDqgFRCu7I4MDotfKjp5hsNh5pC+bAtOYGjOf4fRUcxgy8Ig4UnaiNhN3moGJAqjRByvLvtQj
iSUWwAD4v8Co3w7aboCi+V5hQTix8FZ416eE0vyIhcsdzqXfptr5kbP3LCEIgvWzw9bhbtAUYWRS
XQ5oisDyvKZwGMepG/rbH5R0Lqh7nHAEHZc8DsMZqeGUgPcyodMHf5foGpgjv59YFfKwAF8EVfVW
9ZtdSfcZ8vcEGIZlech3XGkY8gNTpN0SbMWgkGb4jbciZf0U8J+nDOokQpAJoV5QMtnn3nmls+9s
BK6+3owl0khgxC2dPp12pFdgJzz3kxaeu0aTZ6zI5QUMgv4xiDE20izsje5m1qxeIbs6R4ol7EPD
cSsHhRzxC5mzSi7QECrlUArxnUpfwXNYWFnzkP92MhM9XKOhSTKKNJWC+Fyyf08lZ47Wfr9T7rm9
l7Xfm9T/+/J5FVhXVXiSoH/jIxWtPwMTDKG/rrV/dr7TCW3d0rLuQs0M8hQfSKV/Z/esKqJwgHyq
wX/EoXwKRLp+ZqEFnkgtu0v55syE+m93k1vPAaxMItAtvVEk2Bxkz17DL7ciiv32wxZXHUHPA2ZF
RYuSC4DG28gFIboDE2izm9OJCHPBb8I4egtc3meSHHz8uALMtWXvfWiyQqsDaBDH/A6SUMscnfsa
NQoZ7jZV0z4uM9hHPklj0z3ZDaHnhDW9AjvcE6x+fhMkEh8FP84pdG+Gs0P9nAiVEiysKdb0JFiL
breVyRI73+LKCHYTPxmH8DfnJHjZ+NU3v48qB8oleiPhjEiPPw1Kes2X2mRp6vJroz9t4yLuUqzO
eQqyp5h++v7A69fSIF1RGqE6n7S1F+q7d45do1GcA2wV3ouCERW8wrYo2Bkw1VMcUqznzH3vBS+h
oj0pf+OolIiG+lhLKz5RFGZNs7KM+n4GJLAfl1DNy3jwdDrHE2ZpV23W5dje57aUdPCGZNHb7vQc
fnfewKUkP8exNVW+6vkOZln1zsRGjS8G2hogQjWEBGYw6qCKlvavvFwu3MGcrP9bNlYPu/ijQgxp
ufEHGJ3UqHq+Er92gl/74iWWX4zijISrCADkLxvu4gFRFm9XM3r4gmsZOl/sySAOBCXHMap8778l
SsCqa6Llui0Lb1y/1jiD771dOLNyGt3Q9nwcjXatKOet5AK4xi39RIlLF7A4sAXT7IrlLB+fRzM8
woKuaTWTBhuiB5EYMFBiYzI9DSChZaUcAz3czkLPpXt+HiDhDQOLEURuivO8bo56ccIvWVIn1jVp
X9FHs99hYX2w1VyCWpHGhSlU0Nc/IjJp4lSLbHwa+elBTI3e9Cw0g+40idqNLlU7zYXZi98PtyzI
FMcaNplgDayA39fBekzXxx+3daPXiLN+deWkxOlLt3eH6xV7vuIxDna43GmU/ZizMQ64Vf7Wy9cN
vZK5fFX2o4NeRfvotFAc3YJQd0vx4/qKMp5MA+njxiUEszOjyO/pVVpiTzG0G/MqKUVZuuICfBNX
ukQIocjx9iEALjEgntIYkGvyAMz6b+GkA09uzSbX/zbUvJF9qIuJUjXK9LcS8KID7HDGwCkYSpXL
VmQt6c8OfAbnbENLdW3+ar7q1fXKwpHyea9i15WGTN14crhIceHNAp0XSv/WSQMilWqzrT8T5i6Z
BDOetC+DgsPPGf8w64FjwCGp6lH0OmLoPa1ulop0yx6XoU69GYga6hjv3IcpCA7DaN9OZkVX0gBv
XA8R/bz3gT1rQHLvn7EiTiqWtss4xnTAKZ4dIPDpx/g7tFQ7OfUnabKDxchKI0Kj3F4J1Y+/PWba
3UsU1m1S/Bu+0nauSXnbSfBo05HBELFGlP6kJyg/0ovQZzR2XbeK8JPeBvyVXB7mq2jKkUUxxh84
UbOHqljqK53VC4VmDxLo9Dy41myjGPOt2JVDEvmgmTmtxanrX8d5tqaPqx7zDgRTUy/o3z31+yg4
vWVoPSUhAG2umtebIsVtKAZHogBJABh6oqo/odaIpY7FBYGQNNtzq5ktT+WihFnXWQq7mRifWUqc
xyuqi/v1m3vixcQDWl3czrbfw7YJKU8nM1ecy/0hegzCMPBF0vDUS4y/vFvy9qFQczUefaY6yONg
ZHDPJQvz/04JbbXae7Uy5zExcUEvjS2myUS0IqtDg+Gwk8qEWzhbpahkCtMHdT3pKlPsA2IbluCb
mgtNbrEpYtTL07rZEjAiXFlPhidRSGhs+Oh3qsyj07IbiDeNS0m9XpCced3acrJJVGYSxrKq+/3n
9TCimRtR8+oa+4WOqp9MoynjDADKmCPeWSX9VHsyaTn4p3cyhZb66uNYJAR9DgXVGh4q25FiB0uQ
fMcackIOLrDVTJc43zjLoIaMfDakkQFNNflGq1X7XcQzFnQIFcT5YqZsr+ZPU8vP4uqmkqNSq0UL
9ow02qzlKoZ6dn9Sx2rE2XtivI8NQEm7X5sR3TekEBfZ5aSFiw9iWfT7TT9em4Ukx1di2jmImycJ
M0XGbf2Sf8oc5D8m2qr4SCh8kNJzglR5oY12Z+zvyS8Py7U4YouVao928grT3Bt8v6CDCfEWYyMp
YqtvRDvwpgyBU9M+QTOQi2dJnDN/10wg8mSD+aMXuA6bkAHhG6Xbr1KNIbR3WRpEbJFg5btUyheL
lDIqkpUWuLgZd5WdNLBZyT7mpHJ/IrhjjOMC02khJVcJxQqgEMbTSFk39BBry/vnFbFbDorpyaKn
EnCNET73/bEiU7yMp8ucsNtAULw6UYLGwslKkASqkLv3insqxt3Qwohnaft4Pe8dVWMiZ1r8Tuau
C7priZ8mZv7mnrKKvGHfBl73oGh33LwkCmzitofuDskx2X8+RA2e7tTdYaaP6gtq44gHZfI9c3Dy
vfOb3yRDQOllQAgdVJeqj8sv6MY0aefvxT2fovfytdxE2L/U+HSPqeAFR/woBjqITDtoL6hnaUey
mK3yd0NfgJjpEjdzVLQdS60tykrqqbfP7gp+kPGbZH6Tw12wFYapFnbyed9mIn+dmD/Bu47TG0Tl
JKie3Q4Pot+rcEKSa0MNnZ9ZMS3zzSF+ALdeoLSKMq5yG4HTX0LOijHmwGuEMgVBU90uk6RMKmSV
X6Dsd1pZo/033pgJ+2NQGOJTTOC8KfvhEIb7P4W4mE1UuAPdyAeXNKzdQSgVyqzoC6G9Bp0QgJS9
NtaQBwMGpjsak4Vqt62UeKexDFTwOxtWbyODcKcVgVw/JgM4+XIj1j/s5t9PWwFNIyFLcAyeeomx
ef5flZ4c8eiJvbeZL9QSnBcKHH0/vwh/0gq+N32CcKIo8w7G2NFCIgRDViRc3r1eZC6xhAx+5IXi
/0N0nV86un8K0ufS+7IJ00pgy2YLhhaNtlRpXXdrF9A0z/YWOMcYe2S9npQPU1THlSnEJjTsAuJE
fj2yu6clpAmNnyf+bpcwKPLIk+HEd+g8OtyrsSsXN1O3RAyRFCUh9KC0SdV56ryjskLmVmo7uJsg
cs7R8ZTZ8hykeQNskJqV9G2d5KcxYfo9791h58IIjps72ZZpw1c7hFSXwFW25qhB+Qb3cyPO4oEV
L6FRId8BBSWTJlJCBHj7jpMd9n4MlpOC2wssEuGJC/xrLgta0Sbo5WJdEwwdKX2sB2noKBqYgBfw
90KxD9tyYv6TRukmeSJtTPuZYlSWMbPT6kyM8GTaOu9Tl0k4gRcXgMeyzBRCvLqIPWsxHpVvs88n
7DYZrMqqhSHp1Rz+C41Y4rClIJLyfjI+cuH2+O2v6d9qOLDf6vD+euqA+AxKXZsSS+4ISC6ObIEM
s/RugA/ACQd740MXvYzgnQOf6HKTRIagaFOcdmexMcdr4h6p/jJ+lnxsmgqTe0mv8bEBjjUMsvgO
ViSSgcZj6NLrz0SYDGAVhOzY5ynhgjusdlBA/83DniixMUtOwmsi7KlpHtcruCHk9X+4PQpjf4LQ
BY/QeckRinRvBlx7WRYGOCEx6/ka19IUs1CXCM1dqIPIV7kuSTEDsM/PIpfstbE6ZzKhYwMz4jgj
M9cGJUwk2uV1QPWByMEmfmygVT9jXfdvD7dRjIVm/9ldu3liO7Q3zByE+fjiErP+4wDpBafnlHS2
wWmaPq5JtxSe/kYwEjw66vb6IqjsaWedfDbpD5ZPg+QXs/IzelXm1b6yxEpZwJ24ixrPJag+l4Vx
FRqPwXRH6aJSFYFfReGHmgIDrXzgSNb/XylEsrWLef/RgW8N1SbhLjobNeCtIcT3peYr41x0b36K
/9fSTYCSo64HqhAD6tSE1OVHhcuTdmTAzRfY7xTKFhzGLci/V/qxMTdsiLrdolpqytC4k//S8dNC
Wf9trqzI3deS2lS30DbTUeScYnz4A5JtXX3in4eIQVTsnxTCU10LrYSdodQsdR7eYWoNP0B5l8ER
ZXfWyeJv3ELzzd7Ey9IZmpzTtSM4Ri6j89+gA/BKjUs3NESs2JfSleZg2Xz5V5caSr78tv+ZG6fo
LFb+ZupOa5E3P3gnx3V8eqDYn6X9uvYPiNh/or5m7IFZIBaZm0mm9DmOLJvNw6FzLtNganf2G/6I
AIgEN+AkTW/ZcT2KN4KES533PA924xlH6Z4eqWeCQiSrCi5ypzOKRIPK7DW5Pen7e3KOlPtIFHml
0FJ7EtXJ03Pq5ynK31+L/ReNWiydGJnO6uJXJi8Qz1JL344zKFsmOvVD4NOw0r1EwCTkbTzrzcd3
hANn+jpRkt0dbo34OG6Qsf9K7rZzpRDRHwDH/KeO+AZET6Onb5GdzivvJw6775I906YUg6k4Wyn5
lyMnEg1JGO71poC/pN5ioyHC9B8mIP1QZEdIUakWV1+2V5MBEto77xrMjGPNQFIKYcL7UkKBV1vy
ktOyn/jYId3YaEMVZnaToKODJNIqQMoHOkddkA3pBsVJYfq7Y142uo7VFa77Ps4wwV8Z2Jzu7T5B
XixB4p1mcgI2ydF2FeCbWJakdxEYDUFP+ICi0nGziGTV8dMS1AKkxIEym3Uuv7Iaq8xcxPJingBG
ZxKKhotQeiPxvZdHYI46sepNiC4kuM++GpZI/CFUH2DoUXEtAKT5X06yHCL54EGUnhPmmAIIJc2E
5CS/G05KNZjIRQX5pQrS8M4pt85iqtx9L52U66JIG5sJg8epmBSKT5K8XwTsbdANNoGqd6wPOxy0
7QeVkrJW/j3Ft6W8QYI/5jiEMnchmxASIt8f5ngzG+3USCdrt4LeITBHSmEsOdK32ghb47ZdjFDV
jpbg0OVx1tRAuWC3kQljMcWz2rdtzszBTo6jUa9tNEB3J481yUQf+NFwS48UKefnNAtKvF7yPcO4
yblMMUCs5Ek4eZC/z1KMdu36IipivvgJY+FIkJOayqB5cZFmnDNf14fTlbjq684LJYJd3hYbiaYH
0nMnvvjRsDK2VTtLyO3s5LmhbosiOoQHiMS9V8o24h/Mrz3Mp566ZuMBKc8Df+xPEKRB4AohLEci
+6xPbPBNgH6FTIh7rR1JYvJaZUkE+IVyUWSoTCERp1BKq0zdPa5QB4x3CJV5pv0xxruSroWPvVKZ
YIrOYkTuqSbHYVX4SrG7yXzMSOOGwTpNoocFNs9kI0tuGczG47HrNmadPjYKY/kcpMByQFlOiY3M
rjSWHE2DkT26HIQJnO8l4ndjKjP9DedJqOjcA2D2hWaqXNXndH8PkcrqfDIbYCTaRyKR8T9SN7ei
90V8tOOf7efTdggpfhaLu0ClcvUeH3RVVq+i/yYPX1T2JsexL9/mF4F9tAqGpW+Nmrk7kdrHtl25
QlI38xTD9BUyMlwzpw2NxjJkrf6FZI20v5k5/mtsi3CxZCF69swhESbZP8XUgRWySsDW5GiADAos
8uEIEZrgvgemhZdpUFEGYqc7opqAETBrAhl/xN9NxUPPt5NehiHq2BTKkbA/yfv+OzNbMaAb5LER
r0RqCKEoPIv1vism62Ha+3vjN1N6bC/ngdzLim3/moRAg2BLN864TU4XXw/1XNZJI5DPKDr1GEs8
Eaur+Fe8rrUUrDhcPAbExJ0kCevSaebfhMH2i+hQ3x/8QmzPz7z86JZ1jk0IzBL9kKRszOsFosiU
+R5A64dRy/RL0a+1gaUAx91UIHa2RbB5XDJ9ed/dtPsKTcbP/UebXr1zFPoBR9OMUjNAj9YFpB57
aF56PfxCqGdssdmuEpWFODM48Bgz9ciH+Zkgz6DiLcboEL5pN1SpLGivvknJUdVN1eaWzYw1Kx9M
SbD4V/YIYY8uKZmBxeSncrm85SQ2fMO5vkwbqzwiE3/G/TFFRRrG2p2lBA/0TwkywIJZAFlTAdu3
vFzv5EzDmfV9+qN9gIFxpdk/YM9RyzyhAncs7R/52DNq+WqpYDX3OmjNuiTdjSZXY1Jh387UA4S3
j39vGB3+Pa9P/IGB3m6O5hDFK9WuR4Foh1SBaHyhvXLdK6iI+GBf7Bs1aVVtYl6k+LVwVg7wQzNf
n3JOvBgXIjofvq5Teygno704LsY+d4gdWu12Hg/ePyPkP9iO3EPK57SFdWxQBlSWnN43nQscC8jL
c24chqWhrnmYvaEBqR7dYJtdfDzvFoOkFJY908wUqcZ7upYi1UQYFHcGGBrCgG1pCAzK0MCIZbfW
160SJHL9ojTnInhMfgP3QkQWk7BZTSzM9ugmUnfK3y9Hh7TnhYsWShha1xmWrfyWLYwKwVYZG7pq
UcZXExn1nJHgQn4zMuriisnJEgB0jK9FZysOwGU4MqV93EQyP5sAZvY4tYrbkrkZh0VtpDpyRA3R
yX/yc+3t2eCKSi5x1ffZGaTs1gNxyxtw/cExhgFxvGsBctQ5CSYK0XAs+BlF9JzV64QLlIqr1YE+
4tvatrsPac3xZS9AfyzdyyTAfZ5mUanovgD3goaqvvjaDZrGpXiiDOkqB1Sssy2hiePOPJCfGTFC
TK/kYRMFvqH3C++/IRCs/2bdDR0hgVs7X37vldlnkitklh1QiJi1a9saq4QcPZgdgd3LVraXuRX9
iCgTv2YaZzoIJuCr8wh2NA4mbR0iZq/yfaD/dWN2XssO2TRaiQNV5x72oQ9B03dZJPM6CmwbsN7y
bWKups1exfQ7RQlFot4b+cvuKJczrM9iNSwtcWVLY8CvQO6xe+dTAicQucZZoyTvtxXz5yRgEGRE
RJktOzAtLvsjv50wjJY3QU2SUuCwJlQ3rg4/msMEHRDes2upTQ+DVxth+FlfIr+rpjAD+1pbGUWY
2Lx/5k/Wb9Cpf5Z2EE4c7hcsIZt2+LLts69fsf0zBc9RiDArrAXfqCVok9HKeawE9xm5WTuh1Uaq
/pvH/IIDodRTmfYv99m2nGtVeBDIlh3ixBgQ96eHN/4QroXqCaYd3+0vcTAQxhPbefSvjJwA8d2E
nWy+9bb1ZzTXuhWVyXJt7lPEjmRAZr7FNOeEp+BXbg8IcsgTaWCRDSt07vgUnhRwGmGw77vDy80W
oiYZozxJ9xoq5oN39YoBlRXEaclYiRcocMvopQj1QazVYTxKfeUCTSSMVl/dO9TxicJH+I/6fSHI
YAyCaQMl9rJmogZ1+jev7VqctV49oNBy/I5w2/8qrIForW0DaCGWrOJbglTUDPkeEOnPG8/uGOwg
aEZZTSDijcsWTQzFk0FnzjG/tCBJKiV3g1WeyX78pS0mro+H2LXcYJkYqBW7OLQIF0ceJ4/ArDlx
+Vy8PHsCDWbMozf+RJZJIEQ0yxLc/Vk0VDk5jfHq9MbaCyMvsPcufHMkPoOlRF71hnYV9rEVFRFv
uysCJIaIOYqo52DeV7ggGLzY23J48hlmHGJm61XWf0DDY7+mB+3WHMZY7vaPa/UoHXhYAFOhQj3q
+T46WDqGm1CY8xweFmqLDaj8AiDbNJ+0s35dM7zQ6/hAPnLN/9AnZRWzLKn9jLiuv/uLorc7Eaf7
DQztGMcyVzMmTQUh/YmnZCq8l5dCwuZvXizayGWZvdvYbGcVKmvE/Arp9Sd0i4hHyMQ4b8ATRQiI
D853sFYz8pqB9NdA1OfyGLpY+B55xCtwNxULRq8ZwoukOjOfRXlHrNNmjKo9rTIqDKxZsgI1BAeT
XvY6UsSbE6KaIreJ3n5Md9WB3dZeQ1lAhbJA5mCPXl2Tq6csV3lTWo9Suf9byqHzLQxviibq6e4t
pP0vfZ/pvkm96WsmAMj+3pYg88OspN/m5q/c0miABsVDD9ngAzCnjriRMB/AeXVUsIvsNfZeB39J
Oi4Yp4UU5fdPwo+s7Uj/YAJZS8Bgw4oEe0A8ZeuCgybQ7Oi6hoMF0eM1wcHHBFCVvhwtKrMkpC1P
AKOkc+PyLa6r+CeoPG57T8CrDiWoIm0mbYdM2LbFmi2EPdqA4qF0u1XQiTTX0yBDCSOdiorXEFnO
A3w9EJKvDcLLfgWYDEL9FW6zvIffzUfVDc5ChKIHK1NuUYKrNqo0WxOpuTRHC1+rjmsQ27usiB7U
97YC4ibqdf3HidSi4xSrkdEgL1wTZmBXbvdW6BewKwUXKc+b+SmKuUvWOXyKKnauO/iIJNYHIsYc
slhzB4kA4RBMYnK32xBQPkDMQ4n6mbawSYYIgZ/tmuPTkc3twZZkGWT26Jf9Q//2QgR6hEiZlBaX
t3FocQvFi7b8g1TQ8DOAKarJyReWMARWdmeNkJJpH57CvyZlPWnd4Hsdm0ZiOR1pgFXtw37Ii/By
Lsd2mLVwyXwayaGyrBBaAkqIfiQn9wRQ/sNy+rUxr4HQRIPjsGAw9Vt5RXoF+xvNZ/zydJqM6Oak
O3BGphPvdjsUKudWEU0LmLtBN3oEAhbcj57rTLOoXY0lhaPeTAol6LXeQ2BDXZNkxa6hy7EvAMT5
yboFfT4YS3ms0mYDLlJRIg6bdjApm8DY5hLMHpxcZvepXf+3tIJqjw3uU9k4QzoPCH3/xGlId19n
55oXHgn3FXnsIiltZZ9lxzdZwy9p8FugnrqFzr8lmfyL4tSe2Ya8zXxfngxzJPxr3fFF3jTPZwsM
f4vi3KG83vYRCs0wRT11d0fdjmIk4IWDf2lDel5WFnScyVwYa7NsI2QfeDxkVooqjKeXPQhzHxMr
ErE64C1iK/UoVyJjAtaBSNasbWv3h0o9lu2X8k5w5MUj60FLx3InIeBs5C+wBWATsQAKORE4MEJX
M0u2eBHh+mv5CJRHIrXmAnRXlokp39v77ie0KDeIfGwZwOuU8b8K9MNDw5ZjPfitdvyR/6mX33pG
yn9DuNfZaoqFh8eTYbN8HFKY4HIK6W509k/ADXTVCm7SFzIZFS5o0hvq0uVkHLzrMAHxl43+8TJz
rJxN9NyIRHkt4H/bsLPzorQ3vopkNCp49kMNZcLRPQrayFU5csXmIrW0ReKUxn5gCmRNmeXJFsd3
RIWhefBv8AzU8jNWrSgF2JmxmeZj92lxYgsWuPjLPxB87IX1FF4U+VnCdz+86SnMEVJJHtDtnG+g
eDizwEZy8Bov6yTX/wlO11sxWi0V3NHKd/fiGes6C3lOUJDMrzQoiNaAfl1BLbPFItLjJKa6rmeC
CMWgCtydGX6DtpMFguvHAdyrcU27ldZeyDF0IR6veoDzoQETiWsEhQqSC2K2g5Ai+zHbAYzHb9F3
Tuh9uz35FxoEnylclEj/DPnZjCsTq7I/PK0/cB7hoCjwRluaGX5ek+IRlvqXjOipnyOzoaKhip+x
BdeR2vuE7m0OZE7L3UoqeeTvDV7wK2dXsvwPnZV1SwIJN2ZeLgzLQvu3k2cjJUbrtYTBX5/DkB0o
e8A42AEplWPlUt3CslDDRDY3RnP0e8qu46RS0fgQGFb4sknZG1q5GUAJGJ1shb/OcifWujYAR+CL
TR2HGKet4gvZLA9HJPBNongGGLiCYsJpNV569LRy4auQmcoa9viEvXMmtHrigNx/0NzT9TvNkfVh
874IarcLzHv6AXx/n9CqQJHnp0axEI2Hmi+Xt9FEvc8SwOyZR0XTVsnwoxl4uOsipGa8LkOC4Lhy
jtaZtKkqDnvQLpJD2AecSQUpXNCP2R71rAOtcoaGzp3bidRTmgSmGGEaccpW8Vx0RzQ9u4R74bfX
KcCbFXYeHxt2P5DqF5dnq4JpKSRrnvuovHEeTrEoXWzQaj+7qG8lUVlM/cvPz0skE/2sFt5JToVL
pNtx2YD2yMApfCWgcER53v+IxD+Qa1Ql+/bPYQdf08sZb65wPmoKbCkQCLznZ9yExRjNyVSoQLH5
ZIbhJ7O+0Bor6PVxsKlEwLvGI3dQVm8EONT4Zi6wD+WKoYFda0T9P4GVRwPCVGWnh4HHhtM/zPcc
miUiXxGSC32RNv2W/p2R7AY6Bbd7hQRP2UKylej/Jvqq1/uBrEQbOqhuR7zU9Rd0DFsyJun1uH38
Qr+lidC4nMIsdHO54tV2FAAPxRnCcR5IugUxAgb7LYFt9WVNgPlFocOMlEEi9S41KpO0rt4CthMv
BmYVbXM6fO7Tvf8Su+SxVhJkRpFW1CRzkQDO3nL9UoXlCUtDh7iQIsqKBq3reunUPk2PqHdkrEtV
2j4Kcb9ilye+QP5pDAnWmdPEHpozKkIQyJI7k3yoHLhz6NYPkMVlDafaQ8merltDvC5MvAuwRoVi
PCvwXVM/niESeaUoDnHxmAn1Ysxj22tIAV9rKA6iXQC/Xffv81rr+F1ZfyLWvdxeh41sqdwiaP4B
wu5GDvRiCDNkJqAfBFDGMX3eo6uVGCeeUhGXmUk00lOENQOG1xT3ABIHo1XlXR3+5x5dX7FTGxQY
QqMAa5/W+OT5c79LOksMF2NO0ciKa8bqs2sQx3zTfELSH9OTZCrig/A6SeNKBXbylh5Yl591Is5C
+Qs/+9aHm6kN/3jO5OWau4tJaGdEnIy5O1PXzfxy+dnABfQSe7fh3SXAXXcYdV4eVPCPgKuSfUkG
a1yCuKbeUz18m8kekkGOEI3jh4KddCDpZm4jHy7YluY+UIA2dBfFU5v3YmoeSvTU24Wz8SIC4lwS
KH+rUladJKUAjACr4RXsnhITmKGAezP1SAEuDQcb0vCQF+lLmbXQizN69mEGPlGISlTGaZmAT4ax
93fSNbl+T3D/2ZG1fieGZOtwx903c83TRKh9M9Zc/MYHAtoA5+Qh8IeCSFOkLfap0BMqY5mIVESr
MJcXrMJxJioqQNmYk102xguuo3KJGgTMetQlEEL7I590RGreAn9icm2mguM28Oqwp63ypetCdqkP
Pb8bZcUzG+K3s6equYWfE4uslqi8jwODLpsRAUiy2/0RfsjvI1+0lQVlkWiGnwuhXsueQbOCpXAv
SeRxI2Y7FI8YPnY4YEPFkrFOfZDkWUnEC7C8LO3OWsoTZENAn8jrW+dIEOIHFhdGf7WsaMOPYdao
eR6HozjUALR/QurAsHccJeXgoWj6YmS+yGFv1iOc7pDgyrN/vGCYDnQ9Et/pzGZ0/62EZ2yr8cg5
gCzqBv997Yiu68qZ4oIS3y8rDclK4Ckwmf/bibREXyCE+E0GqZ59XPDJ4pgQJdHnWOxScvYl6mYn
y7/3/csEY4ew3SJNVewp+ZEtwRIcuBjZ23g0uYJ2sDKJGsdk7mLWkw0F46TsvEFPCchPLUJ6z3Rj
U+50qpQtvrT4Dxn5hhPsbDOLzwO5rNxIInYTJlBsQOuzYQUVnp2l+ZXr/Orr30EYBJREpoXYYmO2
v1Rh0+2mKkQ3TxRKEKnNcOqavreCN4SGFQSs+d8lqshQKWtp8oxLDgd6NBTJD9GK7HM3SjORMToz
VssdnV+7LjgRCbw1SIKzkGrZZ3ZI2ZhzeotJZaugA02vpEzkjwDC//hHvPFTVTO6gnmytKn5sblG
MnTPs0GosF3cgbW0igukQwsaJqsX47oUCJjCXp8o6XhN+MaGf6gGpXL/v2hLxJoRbPUhTRmILppY
Dsiqi/5+aDOl50uGyvzD2CJPLLV4hO/o9sBm82xWqeekiWNaPWQbvESXcQOSFx0CX5fpBzu+tKiQ
ouSjEOij7v7dgeU95mZydkbIMY8RVM0A5sb8uxXyAqVic7I5xjPaxDGzZby+ltnWSoYTj6XdeDUR
cDlN3i6UI3C9aW5zqQ4eV+YjPv6zU3EiEgVDH44+0NmqGtUh4+fhpLchMzB06hc4KfzLsVL/qtVs
mmH/OONTX6msgb5SuCdCTnVys1Mo6SeR0gE9RPlH+E8aA2reApApVQpKKMLn01u2Vq1w1S6Qhua0
eD27Ez/qeqwU1P6XzzkEOU3We75FmCRVyruSbS44JAkAbcE4C2yPZkxSMao3XMXlCw2v86cHLux0
MKcgpiGaAjUc7CO7ES1vbJUHbjnbN4C5TsaQJH8cCBqCMAn5k6V5I3z7pPxxaOs2jcomy9X7YRWy
9r/8etVre8o2ZKOdJasUmf8pYpik6v8i2bhVjygJ0hZAv1I/dKamvk/yVTNG4fdvfLVO3eXvk9ZG
iVIqbTxvRYpWNzoh4az2ZbkCn9mkfrcg5UhWltCg8dhY6oQ5n94uovEXkLG8D/rw8l6akZ/+yLPF
RM2aGXf3I74iMYtqe6+o5TnSe1g8ByCBihsMs+nV5OS/x3pk1YfLXDV8cOkPB8ejrEoSEEBZ2UyA
xhQoJSxfmFc1YlS3JZN8mTq3MbxUV91DeemBmtp5+VFm/5LUuMqNsEx9hAChNocMb5Ixi09W+iyT
xENhZ/1LokgTmzcW4iecW5gKJ3UG0lt6rOO/ihfYvzcdFztbs3DbpATq+rrOzd3I78aFscCOPjk+
mXGTKBgnzdCxPIpoCt7/rzgAjNvUBdE1zCeKdr5sDQBD/HqHBMK/t6DRJ1eO9kgK+xB2faOuuKxg
k6WZvUDjvKLUgF3B3pMjSqfYaQ0LrXFxtPDRj8lgtj/j7+jDU8tfdoE5PeV0AVV9yslkSNTXzf6R
UqytXN1Jvod0Ye60cVVMJ6xEHAp52IJ+HArAz+ghUeQ65D1zBVEJk1VVdMI6v72VjycZjgXP2lDc
WNsoE+FfpEiryLT2nWckLAWGDZA2AywoRe6EtW6xASsHWXavnGNbbJLimTdtpFwH5Ok71o8NBKFF
g5dPKBuL/fqqS37m/5l9AQoEuq5j5UljSEojiNTreUgLjBuu4G7USt5Qel1dIDvRm9PxlxyO/nVP
A95WX6+orSnuKRLp4fot6cJWeF2NOf/k8Z8rFR+E4TIYeNhRJtYT1DaFmdryZ3J005obnN0++RZH
Zv9ddua+dS20hXae4OkWP90IONp6Z6XZsvkaVA4FFseAelLmv/aoiSfCuX07LqqBO1Bs6eZerI91
burUd/zSh7CLF6JoACDLzxPqZ6IRT0CS5NScKHXQkpu81KlbqwvSc5WTOuFGuAn2EPiLmbB4SkUo
rN4dyviv9trnM6o1vt66y6NAwQ/nGS4vjlyxatFeWdvJiPL9PGV2WyOIacJeQIrs2hN4YSMioM9O
8xXNkyx/eDGGmXVD6qs2vl505c1OZEgeEDHGn+sJkTM4OaJ8sti1HK/Yrz1lUfzFTBGYpyGHj+0A
8XW36HVv5nqAF4Xv/yQvL3mkPMbmwiQRLUjzagrWC+6ukQpOVUxVmPJBAW4uIk9QDB+G4PGeMx1Z
LFOyM85xNmpd3DwKltzsNfho21YNn7pD9PZZKivi3y2h3R8YwuVSStQ9xk35HEXTfK7pUBrVucVs
Pp9KKNeUuHN6STHVHrXbvPBJOdKPNhxmeHaWjBf5mRD5mqD7m0rCdv/oUQ//Z0UTdJ0+/1xSk/b4
E1UsGf83rW+/KTmHTjnWQrNQ9GwUAiGBHKlfCMyot+ui37TbJFFDye3vmkOaVNZ/SrBT+oXtXybB
4BehPL5u5/VlRDCb2P/sXH7Kw7NHuN4I1g9wozJ06TmY+wYiTLlH5QP+zELR9heZn5Ar83m0qGnw
hjcrc6BRxmU9B/imS+MrDTflTedqY80LcxiPDNVk+A5XBvG+9Ejb6T0tR/4MA8i0GXNvaKxjNe9L
JSYNCOAvGvRZvpVWjWuhjVFYdC+vjhzPk1FXg66bwnVu/NhbjyEfUzMxvBpBZSOtX2869ublRg8b
j7f3K98PgUZgStRfU9xa9/ZxDKpQR/KNPCLQog7LAmv1qEn2/Wmj+Nl0wn+DM78o45LidkU6iwkh
Bt4qUIY+GDLwAW7ukF87Xw2lkwsUggRAOIUhaA78FMHIDWL4MrEeoN+p3WH0zj9iTiOrdoVpEpHS
98Ee033FYmudX4KsA5d99vwAYT/4BoEvCCceFlyKdbDeJWsleRtHskSq6o4iToCSOLRMpf/EpqvO
g8bun+egV4oLfRmUbEbRzfKd8x7SvF31JzUGXyJDKU8AYg+G2/ULimKXXwGDS6uLT7OQOZDu6GH5
zPn982K8Mpournj5FHT/M1NJ//66O5CM6i/jIbwvnudkLWyxQW0fwTqERXdjWRVWH9Tj9DuV8n0r
01m6rUgUQrwVp1UhSDvYmFsqP/aZhKQsRtvEGepRk07xRfPLGg8wl1+5GgRji+7pOBm8fY7eUnKl
Ils+ppYMfdlxd/Xguuiaou3YbsLrwz/URgwoSvbzBH+/An1ccsM7K9L7KkWdKTeNTveI6x9zDY4q
AyVcZ/eP1KvSZEmqxg5+/goZ9oUYatZ6ltmCtF0Vj7S6GaJrFo9tmWqIG4/+2SbfUIi2dpwpnnT+
rKzFZlqnh+CNgV0djVu37gbQapDSTp0o2mcaH8OhXakgCvrCyu/sq9CJ3qj3o/C6tbYb3jFGohD3
XClf31P+FqEXIDYwT1mUmqq9mF9pw9Se7jzexD+fpOZxOgffidpWSwnFBLhXgfBl5oHW8xshPvGO
zA3CamSSqtTgwD+ZQ2XspboMnpP7SjdyXEXTLAo8YuvZ432XFiaZqsDHsAxYmZkU9Fub3pggxBek
Pcxvw6GmxQ3N8E0/RmNbaLFMtPHiaz3jgw8Y5GwYxzWcdsNaL1qsApGdzFyqOgabWKIy5+N8dGhJ
EuI2CQ7ntrDbfZZpK3wVj5rPr1gNzx4juaLMsH4yOp1svliOw69eP2IESdr16n9KohZB8h3PnhUV
P4fyGP+nd1P8ey7hNjrApPCm9ADafP8g8KW6BR/LYG4kDW7mkWCTVkGQalt/SxTJwNbn4TZpQGj4
tN9TOC/vkMxWQ0WBV7qQfCsJZln+XDj7yX2wVKbPvzdaAvDsWamt9WnvfSNCZaXbS6vcl2qivo+2
QL7LZ87xrqGB+64aOs/niFlz0YgUb3CfgQ95f7g8LjL8roy+aLSG/15qRRb0cIIO+q3R8PRC3QPq
ULjhkY5+EFAEskZP7rfg9PcKvbwm0CllStoeloDktfA4p+NHTI0cieQkkWHe9Z2eU2ubqelOCrZE
pvde4MFNJ+ECxiDyOVNKCgc/QUDrElZbsLuouJYrfAjSnZNlQO4cjZ4YF3hVEW966mlb8SbF4iRi
v5sXOHl0wmuvepJQ8HLjnvEqYH/S0ezW9kwgK7g22of81c/QVUPmNucYaXjuG/n5gC737I8JtUsS
7w7m6CT/wps5XjQDe9mkZqVVjIBBR/MMTZ6mDQ3HgOMDJKPkjDX8bfRiL2/gJuk9lt0CS+Q72do2
zWddyTT5gqpWZGtn2Frr/NTdgJGxvUSbrZb3nM3r8KyKKcixLBdMBjfJE2p5pDMMYlHtCARsmcZZ
y+RtK9e04lZYE6IGEHmODxt768AipmIJt75b6al6U9+xSTjcfOgJrIIV+GZd4faxB2i2pSGZl8Xa
LOjQfBJ2USlUkD29w4ILJOKRj2EFMINx+Eco0KnbSbFICuv9n6x0IGcyMAjd4q5ohEvPWftwJmHQ
Lr1QL6oTJM4w5XEXEMItLrvEfIqdIIgE3vSJPKaVLsdscyVxuEJTXL0KE7ly4bvM3NZ5xUaxUWKK
xqEnM8lgy3+IGm1WXIVNkY7hDYSa9/Nl/yhtDh6TGtyOslCbgkasLBCdnp+KboBFmhtkFEPlAmrX
9pjj+jqe0M7Sy3Plt1+8V8DwZdW1ldJHn/iyGbE2IpvuglD5MNlohizOTkjqQUb/G53ap9gr9aaK
TgRqZ91KK1F1pkDMDMbEv6A5wzbVwsckYZfLVYSTvEhvEYANagMEMirzLmhy2T/gtgRkS0AcrvDL
ENJ+8JZzddjgJ0ty3WGEZvJstu7hVP2xGwzVx9bDQMkxrMyB8+DwUJ7dRPcFk3pUNs884nQ4q1Rn
9h/MLO0DxXQh4zOW8tzE6Tm9DcZdP9APxYTEiDjCHwpXZ1Bvtg6c1du7kYxmF54kRVdVejlX0U9H
g9asGRPmHHbIglN4PNaYflTpOSc+kBfrxlpd+GpPAOyVR84ucjIB9RDJ5GWit3LRkGu4SrPQAi2s
kDZ0pApTCKpAeYkVY0vbxGWaAzHT2dGXqP5kuqKkqAJqnjZEQl79JNyHYoze7ulk5yldUvXDOAiE
f7iyvwvTenZf0GTMDMmCNcJDi6pqLa6ClA/atGP5pWfbG/ET6/xSg+aLrPbeF8K5ZLudcTxkI5+o
Yh3coM7h41DjD0233G3doJxGAHOprMsHE3kZ/TIPqNKf//mCOs77J8Bi2GCc/QXjbJYy1dBZih5+
O3c1H5TK1n8knAoNScrSzb5Ri4Z/TMMnm1uRALYjhmHjJdXOD553j3PDsD06kdAHtpvz9P57F9i9
EP9C+CMCpwFEt6zvm36JfYP9EyedW9BxME6p5VORKVJuadHDq7CCzFSNTEIxC3g0GP70OSKnWiyB
r8G/Ml7z62MoaN9tCKhIdiWzD+Jff041BOQ9INtrXnOj2cuBiw09KxLK/nYmwULZjY2ee+YT4hC8
yfrd1Kh2V4gybU61B4Gg5Sxyq5mLIOliaVrYa9YiiPXQdisBnzBvjSreRvk8KTupkrTdTHtaaDbZ
ngneqNy/D20L18e4JvKG8Ri8gEQg/NHfdC1ZF6Q6Fy/fvDcQpq/TDbFNqUTxlVD0bjWmEkU/G/gB
izBDLU/3aBU3qMY+G/Qed5I87MXUSu4R2Jeb9clixrjpcYy2HrMZMEqebhu47iVjmfoVNDPkY0K6
TijMNJEX+hhAWPxM1SDEgaZZGD+dwaE+fsbzWqEjJA+cAkW7W527HQCJ/26OvTqCjrz50I9/6Dd/
BLcGrFFhMnGvRHjRlUoIV/o8cKFOfAXYswW9B3huGAZW0/g3S3KxxVuLaB7Twkyy4QP5Uz/+CYv1
pGZJe+1sQlSfi+vF3XxlUejGwGGqk/56zLPes2xDMR7kXv6DlrVE3KXYjktfG65mj40wYQ9g4AGX
HufIsgLU8BbINRaqfbRrUsg4gZk+fbGfKf198PnppzrPv5PrjQ1jE4WdlXlYJs5Q3YVSVCnB8mad
wFN7D3nOYW4IcXthuxjkx81CuJ3oqxKMG5/SO3BWLZotT1K4BDfLzXe5Q54s++Wot95utQr4eq1R
X3aaqiOvnnPoPvvIB1lyQfDjub2EMRxxpfPNFBAHrrFSMcHdvwNyu4INDpfSKUIksmamnPbhdZMJ
pCacZ8nQOzjtZN6gCVJZHPMX8ySJIOUd0DL9TR8myahE2SedBMhjyxStR3YbSVVkSKbUTEeYxHg5
kYfjfRTJsEowF8A8+Byvpqx3SX+x7azmVCXNKq00tac+pLsGEoJD5nv9LGFJ7tUqA0rPTAjXzWMg
gx0CscgS0iGfoV0HSaeK0CT/gQZHHFKQKo5LZo8gFSrlrDN5GwIIa1qrdSHLqWUmDz9pYgaJLz/y
vvWpLGXoBVmBLZ97/mud+nvxn33M89q2E8cxEfhRnjUSSf4FSxEX86XvINB8r1wZHjxNoFwdojuP
tBd17Xa52RFSZstIz+/NvQqkO4hpIaMEXjGKfyD5B/RAp9rmD7sTQZZDRBuWquZOt91oumvbu6LK
d9KrArZNzLvYCjFhuTPRvDaSjQ4EKQGnXSXrRdIPf8PrFPk9SnjgrZ/dLVhiH1oHaci8uYv0H2ff
UGUch9S5lla0/cpHWbGblbVviwOSqtj5gD44bLuLnvgdKLmAnmcmq1CrIDRCMfSrj8dpRyw8BMpK
Q7mRO1PI2GP1r0xSGnMTjQgzQd4/GVCgKchBopKcJ8kf9EJO1MgkZdJUNe58EqNc9YO79jOBC3K3
YTUVrEfAsQvzoPQoWmqDeK355d2E/oMyuaCDscivWt5tLLyirie0oIQveiIJrs7hxlCvx0GEsxu9
otdBqn64Gin2z0zdhLEViXgL68w8UHTDW5RrRMz6G5kijmBvWt75r0yp/JKHiHLBxtifOb/g6aA4
Ds3u09sUODbItb5UJMimJQbeuHexug6UtwHDYDpN70FJiM3ne9LqEwEVE59Yw/4Caxk6IPkm6Crt
lfpbJPdHXqobNZJhq12NZeWnGzh5+aYjYoQWdzl5BvqV5lGeNs3r77Jxr0VSZow7z9o8mtfEiHlQ
cdxDe5qGhM0H0SbsxjwK+UZhHW1MZetl0K7gSJhtdH+dm03vBP+io6eEusVEaHa8HKrJAhwK16cB
b/T15kLFNRI8Vxp7y0zaRzcPND9EZv6xa18fN8p5IXnV6JGqSqJkM0mS5qgmsAuOgls7hX/Eve2l
p5DU++JZS9UrXLrmMg1stF/6NIihTgjKThkMJAMtlFtbxDc4tWtOtjf0Mx7BosS1yvv1/ThZ3kiz
21SmGiZiIeXUOMV6zOTZDZEt4wSc/qE3Ro+bS+lFuNNnhsmGL1G35wwsfVSJ5ySEXLCYMjRHhbXG
kecN9E6W6KaMjq/gtU2sCysx6rBC2ZW7adOxXIgKEKqFFQxzaePkdPAMZWDrUOui407HJjNXt0/z
YFDP/MEU5/ErErYg2SOxU8D39JZMVcUB+Hcorsq7pbMEWpfqcwXTbFwXjZWXHhdByXz2L1ET9QP4
QcAFV1MX4guGJU6XKuL1WNdFrjW0/uZN4mda8uXrHPgJ4QlkFprxHwrxMyutlTmV+dMOGMhSVUVp
/Ch/i75P6li8gQPGgGpoNJV6NOq4C5DPOsrsCP3b9/fXdo6dpxG4qNQWNissD7S8sjYV7z1ggLTg
/s8IG0RRMA9VGjSUFJjHiQdapVL+wGOIUE8yEaWnJQUxYh7F6JQ3QUlxNZmjIIkR6Aau4yFrIKA9
/f1PH9FR97iuf3xijjUIX7Y57BytAxGt83uCqP+i9RLqecHI0OuRogxuPLv9qBNuikWAgb3cUt5E
czUAcSIyPPa4ZBGNE+UXZQP+3YibLTisjtZeHkB4wXH/sgva5hRiWVIN6PYSc8Rewo7BPxM2u2fg
peZTLDoxhqzDh2+gZ3yChzDoTp2v7yi+/x9PEgs8CDlTpdeGhSIa0a6gEbfeY7dEyMIvrDSnhf/j
nr8VoLITWD+UTvNKpk/mggyy9iRxuSj6lIPiMWJbUJwWobLt7MAr3+1wh0e2PV8x1KT9/kHWPH4v
Gyzw+sFz1ENOf/ag5UK7dM8NFil4q4Pp5MTmZKKmbg4qlXGLNCCVL8lOG6/wwJzhOYearFECJID+
wvFyI/qKK8p1LawRLMQyxX/uFT8KKGswnDH9ffAgHt63EpngDh+Be+F2NW/+FMFgqk9Lse/vkBmN
8Cd4XaJ3H/PznwFt92R0tVpHHNxLPsObRHGoPh75WqCqT5oJngtyeFynWW+/JzpBJsYTlFvDyNXq
UAh0MEm4zevPuW6dV+0yFNr+opV2QKHZW34KjpiYEeWb7MFiscW1UbhW06vokHzkdBIFtP7bgrcN
6FQDpIyeHP8tzElEhSon9qCgMeSEf+G1IDdUumb6hDlQ8Zx0YsONLuF2kjsPMKoCzw9LxqucHXCe
oyt4qyE286NOESzqNPs5mL7A4hlc5dih2DoLGz261pUMlPu7on9pkVXL+tKPC18TMWVuLWWEl+JA
e2HFy018cvbH8uPcO7coQvdNsGMfKRznp0H1Tr9ZVd3z8BXhNwWLJnkaVFYcPT1ix+28V0v0OCOX
n9d31Kb+MmxIGWCKpt7myV/HXc+xArdPO+TVFFplfbU2b3MC/F81kYgnT2PNEwk+IlMg4IBWf/l9
o5Aj9pr8l5U7aHUj7CkIoCQOa/wboE7EvQc51Zb3fRsVpODkNyAgu6Oc/HuROMfzmUM3gvQz9XD8
FRazJNG0veUJj89yzOyiCEbvx08rK+pK0MnPfINyhhaTzi3jYTzyo5C4S/A2iv0nYAjVlyWsvyYj
VIE2NkUb8kL36V85TnVY40nhUzbJ//nFclO3OHT5JeQIPI4JmMDPbLHImpf/WFhOONOSRjbccGj2
rZO+M4LUwxHdYoL7rpqZIldCDKdZ7vZXo9BaV50e/ZDxWr6dmTvnos3YnrxMrKCt6PS9nrRrD1cs
byFCr7s/48z8+66sIZOI0esaeOIvRfsIZoJx224a2BgdKMgd5so/HTYnEyakCCSl4P5vqyCM1txb
4MVNdQjz1yGhebEJvbsCbHtus9qN2rq3UHs7owuIAQ11zZffag7IJk7Bp5fNoFU7PJcHR+N8inE9
nz2f2qdlfmWSj3eto8WIRDA4bOdPLpFIJgRw/6Vt3dh2E3vakMVFhZhRYJQ6ghS6Wv24Jkkqgm+D
Laj1ymI6leXXi9GVbOTz2pQnrWPebCkVU9seccG+q+KFUWVgWMAcrKGfFbv3ulBrua0GYjXAt4m1
mJ5PFMPsU2ss4gd8OGUaWrCKoiH+7GYffh4adis6swctjammEaNCaNrdfuwJnjWMrLc+Fd/shRNo
PR+Fkl474opBJE5ao4pXnbSGELTXwCuG6sQInPrBrcLGc56btddzOAc7BeURba8jfAbfujyBa4cV
mkpPNG7jnN5/B8n1vWlsCDfSBnMzqemiNdXFfWIuRGnszsYxL7eB5T1w+Y805q6zq9O7H+jErMSJ
3jxHnT17XjJOh4/ScHu26Fgiccdhzho5kV0wHsWnlBfrspPbGzWKQoRXwYtIQK9j0ws/EZbqWGEQ
V3NHVqwx2rFxEz99uMcaKtSmV6ZMqc6Eq/0KsODBu5+HBdGI0+5xJkvBKQO6pf3saCK0sPXGYhc8
AK7C9FJeT9CIJJfMFhJ23aCdutuh9qsF5lfebS85EkYT671Y9HSAEqFTsDqeEI4eT2iugkGGC5ZJ
XXxoNVQj8XJA+ET5/yx/fn90BrUcSGkvRzg6i3njoHwspodsxpLbfxNRSnjDFA6md6nWjv2Q2U/A
3uDeWfL6WAvSG1RAmZMqgBH/yaGbI/4CmShGwAPEYHr4iTja3reltsZldsH69NVN4d2+Ub7t07cT
QIfSdgXrD+5trMDK7UM1hkiJVtJ4tT+reWn3zsbqmG6vK6a9RACFe2v2t/VpAKQtKtDkN9xcy1kY
2xlZzITj0Vm1r2copmI97+Sy0a4QlHT/LN+ptcJhV1KdNLyL18z4AOfByFoMv5NpCBEc4C1ssmS/
T3TMi1vHpTAPmbD088pMEk71kYkcsRCB0q70UKrlJpBbuPEhQl5ax9ekm+Uel/4jhSqHrcAhqVym
VmA3m7+Kvn3ZBYj0A5bHocVfr5I357Bct6feKeO2md4OCkx0dmdsiCSYWJITuGdestdSoHEfGKJu
tP9Sbood/y/S4Gl2obTZ9YkMo94oddu44BIZxPLsBBLpoC9oM9m9l+SsWlm5fUH0e77qpvrJB0QY
7QiIfjcPWNiajBwipSNwWd1gr25DeNR5PrOwrKAfIVFK27IDTDDfge0K9cZVjQAQLBIXTLTATraQ
IJ4YB+w7h+mHloeUT3URQpG/ZUgZQGH1Fmyi/0qOkfr9vSLRfmQGGVqGO1VWISafm1ho+rwjhZIv
HeAJ8J8LZiJsAZx4w+w0iTwUe6yTkII9PKWXAoFlCp7iKRxOiye09T40k6zmO5vrPvf03mXoLFie
9Mk3PgiLKdh94D35wL9LWuZkOT1zU7sGMJAktGAAQVlfv29nCFZ03jFqJMf8jnhPK1lh7U/8gayk
mtPsNGct8yG29sFbC2TQOIiuWy5zkOCES4klnsR2BUjf3LnhL5r8varuUjI42Yxbi1KNMv1E2aVC
XDomZSnFxPiHErZUt/OHBKcNLgkAwrSgH0QA0IiqOlur/0sOX7FCJuInOddsDNshOQqh7AbbRhc5
hbIoUdTBPEqz6dKpOlOWVKJiNyT66u2mahmgwAr1U2froW5t9pk+4pIKzbIp3o+kW35GPHxeshvh
yZMl1VJ0G6cH5eZQrrMYI3jZ/yYxKXOkpPjC6dOkk9+p9oG9uT+GoykpYWwc/D027EIiX1cJMiOa
xXKW2P4YUo8zmvYqkOQF6i9G6HXZzJInmfdZxpUFR/3b5zp6RHLsT9WibrNsp9j/wcX5Mu7ysQ8a
kJxSwB57Mi2ZCz9a0T/jNr6ZESwTCtmR722z2im7f7TWew5HfW5q2mMWeV98YafRHsyUieJBYrhm
nBws1cWKfPx5VRn4WkcvS4WzR272S40M38n0VZ+69r19xIeGz+/GdbWrgAVGTQKQWR4RS4eNBgtI
SPVvEJJMbzw4r/qecR1CDXBugMqk5JDB67vc7dAi4WukBDiF1pCx+X0nE8xyFb4L9BEYjLC5zCHI
5bcHF2PSprfxn9hXuICbCB8/7pKUwFcaUsK9rsUjA4DWaGfQrxQXqKpV7FQNMvFQ7WLTKC4fsO87
60/Fvcq+3Q3tpvVQUxHre1xb5CE+U6AL+wY3c6lkP4aO71tiy6aVFZNhGKSWbc1Q1N1cqUh3ygTZ
mYj24pdUk7rEOpBOn5QxbMQ4Bfln9Xukz/POR7QROs8ZdqfBEocpVLwVBhNlBRFJelc34yM4aY3d
yb/l462t0A9425mL7USFEPIVIhTaQuGbdz9JiOVxu+dwxU5mdOT1f+ehcIRSHwi541hotHDDErxK
/etFBXPgPwzRnwQiWaRWTjNTgw7nzSiDN+NHn2EOuw6jJhNs6akaewrsN+OAVcaK/6ssd/VpnXgN
NVPQsWEUxhVVzxB1OYsXWX6UC08/zg6sCF0UhBxICb5zd7ouD9hkc0pjucPPiEaAyLVDuFSMrT/W
nN6NYR5oOVmC54wIzfQhwRKtnHbvUDwYe9K1mg+QTlDj561sOSMtQNlC0GuYjS8ZjE8rw/Slchol
T3ykG0P594BiAlLWeywO3aS6EOaBNYTfudqFWMHvycJCJb/7aoJw+QjEyzS4lJcsR121CMBpSExB
1NWDJRlcn5l5sJrhUurDI94a/s37iTJZjS4jzwuVLL971FptObh7UNnxfzyyWqMDmgaQ+FUgMuBY
Pqp1PBRzDEJWCSKjdYmcWuHRv1Mzk80ptRcrzNwx3AitZpkjaNvTj+dwrB2mKFM5tMfymym7uHdA
rg43rSWORffL0IDQSwg7EtivwQ+SikndL3gcViU46MXckPaXu+aDbC6jvdP6tBumBKhR6ob7xX2b
4sDANwv6uJ2UrFfBis/us9cvMp2CnvMwgkls+Oy1BBQGBxYyetUfr2P+gsRVQWx2A9dG3EqxtQt+
LHETjpDnopcG8qj21Xsqjbgwr/OS4SWC6k4p+eaD/CTpLLcVWNxi5/SG94RNIl7ZXjXOXk60xzx/
gKsPrtYm8zsk/S3T+SJV2cIQ9pdxvCM4wBVJ0NdUDoz+gNZz3n2RqKPXxo7t8kBAiO54xgi32dsm
c/hgf2vnua9M4FuT5wzNOJ8K1+fs8p3ww1C0i+f2k2KpewSmqTazQN66trSkeSY+kAFq9/w9wZzw
AN84SmCw3/71udtLBXqIU7hTC0+HvkJwh6+26MkVf5b45YhwDHj2fPnTPYMjavk27RtqF0teko98
cwwVgC3/kdjALFmA5W3vDgnzXtWphFXlXyQJqAV0tSMH7e2i/+JgZpAA9h2wmqee33xvu7Ktlwjz
bXi6HFDHPFFqZMNWHPFe5JNfn6L2AtVygADrR8L0K8Dx9VbAYjkolxAppSZgCcivgxdDoMoEDP7R
vCzI1AihXVoAQluYP+fBIYwLYi7ZxtRh2h8e/ns17NCik8yBvPXV6ZE/GdxhlW2PT61chVIgab6T
HIWZni6rIs5lQKQ0wJ58L37GLAn/EuL3cIHoS9lm1bbjkDtYFfdNm0KSVUYwYsDJSgfj0z17ykuE
iPo81q4ThEqz7jn1lR1QkWm33HXPg4toWo9ZBbM1OzWUJtolB/nw9R98pXHO1vSsHTx+iq95EIZL
pzKdjS6aWfUCZb1n0L/8N61TuxogQadT1Vvz+pe4pyKzDmiLf3Ci4YGExgERENZvF+X2mVLivFW9
n1pjtaVuXRqWsEBEYtP+9soNY3SnTJ+XxcCtMWUuWHTIiUkrgbnhwPCnBLRASgAqcJm0I2KgSY3v
1y5n+Mqw5m3nuzuy/VbJr0TgRHrmEuGofYGifjJ3tnO0VJAoJH0tIobNX3gS64cNpFJE7oq93M9B
maIaS4z25WE9GZcvLfOuRG8l+AWi5RURRJWcIY0gGVA9TDBRhLOvI8rB2nuetupVPTfuv83plwCd
eooToEiqDOecE3KgcLdcdBKOfDTHKq6vdDlBkeP8o7ae2IVQ/gVPNOedYHOE5+mG+3Sl+yPByvvK
kTADWWWdRx4Hx2v6MmTFQkQFzxWNSWW5NfCTgmRPFhGvCkHSDxtZJDNXjbFBWBy5ZohVTTL1HAT2
jQtq1MOezIolr6NS7PieTizgtwOoOuoPgL2GOaJ48LFCL9Se22AbEeybNSb/WjJTAcCwc/X2n3pl
iZd5rQRWBkWw7btii2MBTLwz4tUngpiGgUvyRjUNB0Jk6hXc/vmwOqf+97B4+V3EmtlPAYYB7A+4
tsjcpZxFR0WAcTSrE7O46oF3v2S9zqltFm8MkRP5srNgCWl7Ph1op4zjj3/5UfuSUdfxb/AS72TD
NMUZakXr2jhX6o9vRjkUSJAgxC0+va9LMbqZTYrcExjXFGV/7AUs1PX54F3ps6EmGQCedUvodmh2
jYj8gxG0hbex2gVdMn1xWC1m9hy/L6K/zc6MDYMzhdb343AKs/OMGCV0YJ/eTec0spt6/GihuAoG
oMf2Bw1mWie8HZxBx0zSvaXPWCgZ7gL8hO1hEPZkKl8jurD8AQAA1JuZXdP+j4H8HPm8dlbrRlag
4hgD47BvH60tcP09m7UTO2Z3seVgeKe4VaOzJ0+cB2PG5QvpHVht1m4AQNj3RgvSSmmQguEr5Lw2
37O+Z+B+eFeaaS+h6o4qm1nGvvCcu/7US9sXfXxSrBRunDmtUgJr8PZ6OtHTX8Hq+Y8dPfdQdEVg
zdT/iDOr/LMfa0vS5AqtWAhH40HzN1QIvQq0CwgNslh7GTui02sjdLoFyjYQmQNOVAXHe2pamERp
Ivox+285tDJewdmq7W49ImgDX40JgTu+b5RTp5//mNnheSQlixQgKD7mEcyXZGM2pov+AMfWVagf
/73VQTvMU8YmQsNlChCZ0J4w0AM91/Ch6Nzv9iFNsn8pYphLw67XUV9VfiCWZcUG53WyuVuQnG5r
GTVn18yAWuDzquTEDE6Jc9+gQ1NEYTL+U35piglHUB4awvrUZIaTd5hEERQ+V07XWhjde/xT9xp4
5CdmHz7NTmuP6gKsQpG4ROZp6vHPrb3hl8nXQSfOV/yIB94a8pelL8xLd1Z8a9YPwTcO2hF2+DBR
GPGEFuccLqCJ0/yJRHSJpNcXPCxEYSCzpKrXIjEQTjImmHPQk4LcVrc64chsxbxDkMJLzQo+XSTL
DtSURgTFrVbhRdrFXTUx8YHGN3swQI2pd/oEeQ9ZNbnMrWZGTAXORd+Kv41I7xAzyg5UMkHVPdXt
zCccUtrzl5cp9g4z95dTC2DvFueuGlphcIbzkPWOSfo8hIXtsU6Y1JwUyp+B8w2s/fiJnH3Z7VOY
7Q1RABgWLE7lmU3hBWV92aNLHWR9Q4zaKFa144FSpsxminfrIQKqCTg59AAmHoA5+Xs471x4HxgV
LhBuEZ+NjIqvwTHLKtm2lqshuuvkVZVD3TELXk5kMiE1bPj1wZc4wVk0j4cY/i4L0tJP3WfkWdgD
GfPQGQD+4aIti8AzfCfIbJSCmDyuzOMUH420shhTGf47JVUQY2vIAA6HBW2iZ+MJY7IRUjy1Nl9Y
IG6UdAVi4CBbHXlbv2Pesm591kxQ/5JPDVzi4vkT5VOuCEijlXvWw/iBkM4vAafMQ/4PDDctOTVa
Nf3wp+8bvXTh+jNicCcj+ljsHKrzi9ntgM7H1v7grd1WE8LeJOkzh0nuAhTtnlx+JfxvYprBPsz0
ctrt7NsxppR/7mQwnC3V1Bt0NKxwU+rlTpsMC7dsJgcAP6/heEdJd8I3HYOK3CTWXulkeshSuEtk
UeINt81/vHlrXZfCfCxwgUv3CJft8QV8qyh7OReXYQnt2LkFsybrRbuh6/Fg767NAsIUCMsJwEGW
Kw+RCykTBGZesskQUoSXwxxNiHIx2uFHTQl5oFjsyWH+Ebm3YtQgQG4SkEaBJoCoGUUqI614tnDt
jenAcOqC3mNOKi8g9blVn0l+nhibSZwuahp9912JVlq8yRKMJ5vVENccHW0yL993RgR8VtnGzJv1
yztKSE+CMOnICvsHzkoNtfaPUhPs+th3mRO7OPy9S8iN1PmjQf9I0iKlcsoa+pH1thng7sb8+BTJ
hiZ3L5vUFYMEBN+5oWUaiLJNN6hoHKmxJA7S8JBwsBeJ7Pix6LwSdSMHDWcsFmmuKNj3bLianKOL
mqKGAehoT3Z8UHOVkXKBOLeHvRxncBg6Vi3Rh7Ie1OviyXh58EA83ABdYe1ofYYLYVsubQky6/B3
PdTHBE1h6Bo/WiEe6qWOP4ec4KvNXUKW5v2pt74C39AErurMruAXKrIco0IcoA3lZ3daLYo0a55b
9Os9PinZIKd4GQTayWbQhIHZ0bFXmwcrhaGaeZXKhvqNm1yEefZe/1z9BKGfKUAXs1Mj5GP1NUVG
PKJxfpBd35x+/bzVCoQPQTbexNd4jNfyz0jfmz7wpaUT8YuomVZeCumBYlh0aHyi5/vge7rMMkRV
EzzC2W9+9FjnVKvUFZjWPJFGgmSICsUuBJFw2XcusK9KEA7tOCgF3h8UhRqqd3tHYyFW4fPTOvXG
NnjQNgY9akX85gA01AI5WMvjDcCkdPc8C9nlcfae9g5G3b/WJ+Zf5Pvgg+9daOJfMC4e111vVVHf
MIEUsP8zHE4CkFEh50/2/97gQpVdMFjPYg1QKsQFol7UswvmF++PbbNwX1PzSuez7phZE8mTjcst
6BVBhcbU3oQrKLdh02VFr7LiAsbfsPZf+zahctqfb1GFaSojEaTVEdCuIJ7SSY4ofIVvKAIr6k40
MLTU0lJcivvLweemAJKStAsi/JNH2cU17xuXIFTwn5pyBUNbGcZSXvIuSALOkDNDMIgbe62MDK8e
efYg1cTKP3pSzQH7+88gsy0zjQFPQJq4SGwvSy/wD9ALK0mYLQ6kTyb9v5NhZLqMZ88q4mBTKKuf
ZTyiq5RYan6f0PSs2nlexTG+59IBNt2DSEFMNctExRyTsTaPsJjM9uqFyqOJFOKR91aO/MTAVSLI
6QbMSZo3aPb7jVmYhzMxhya6C6pBGVh6cALlimDoZ+TFCkGft1RGyrFCpQ0kRRAwOssAglSFTzPY
3m65PtAtaRczls0U8UWB1BI6OJm6oJCA7ucDet7ZES9dtCcqJuzJlrbchVu9hBlLTnzYJInVJmaM
nk6lggi114hHf8J5ht/OcHV7oG2APqi4kaacEGPuaevAwO5QdngoT4ZVLlb/oenQ2bqtahFUw6+z
20UG7UUQtOAJBqOPXw5k9LQOXD2cVQZB/mtqm5NXrLMlWi0cuWjgMYOfQaSphmMnnlbQTByXC+UO
YaQeQroTDVahklglfHCXLfuNLNxugNDibHVK2DwfwNR0G0SoVYQwiq1oQrrx0kXEurZDm8NHgoyF
TZswVzDk8uedCkT5AJtldx6eBvJzkLkGex0M9pgniaQcjOaeFy7BFIfjko7r9wnaxQfvlYKIRwJC
F9Ut94NDSngAM7rUPJ5ov1mH20NdLSrbr7FDvWaxEier4VkprkTG8RxEZuK1N8YpMm2YVSSgJJz0
pljllIJC1DHegaX4iF+LbrTYZTG9lV7B1qakIL85NkIyEUUTFG4elwjmxTeqKi/gmz0HJ7kD8jVa
uyRTZzuQDNABsmk+y/fVElY0iid5O2jTC0MvrXmNiX3yrV6v2A7rfLgnJKHZwAcrisyA7mbFyA4z
E2mdre20JauqF25HHn2zYjOUiMA7bO9Q22SYRyeUUwiFcnVvMHxtH/kVmbpFCNaMDEVrlIFq58k0
v2D1MtYpSlNzVgwM9g+j2Xn1HSAN5bFjn40s4As+HHxvNqcr18pX87jHQdSUPynswepIAh8eQoGg
RmSmowDHI+ZNygOdjKkgq+Zx6+Dbb0lI0D75lPOCgSK4cDom3V3NKxBRg0xr/6QgX305CKT+Sn9h
1D06tIyFlgTc0yPM6zKw9yQj03UjKoMPrC3JcfwdPhSEV01HlwuBgqi3ybODjwQvNhg6bQXj9b4P
ZEOz9lUc51x9MYTKeL6/k+vulWDgfI7Dbq436K1AvHtcdEd4JRBmLhklWnIunpCmutNNw/XtB9zC
3CWjWurnyukcG/OtqqHu6T8GhVI2rsxEa+QpNnJcpaI/12/4dTMl/SFDG5w45FNuiEER58XN/Ytb
ougJK4Sk0ELfxR5Sw/5UOOETRsSXPDvKP65c0FCZurXymOzkhj9fTmazK0/8I2JXIU4hbSpdhKwB
I+0qL47Lx58qzRNKkOXEuanI0m9r6g0LLDimHunJuBXywvXZy2uSuzqcvblxRDDtP9IHIwbLbPqT
hydh6kkxw4qRzKNzK2rpo+3gWX4IxOsulgwNLCAF0lMKwFa+t1YBvDTYhZtJE3QZg/v9e6+8Pc9C
5FElIkTO6/zpB9A7RDT0E0OJ9NRM90uRr30NFhmZ/jqM/mWUPKxYpDH4XDmH5E2/Cnal75hINVin
mA3PxYxfv+ANk6R+Qa078AAtLQ42SoubPD8q6QA866e9OFUFbZBugTUZ49+YpFJlHjuRkQa8fP+h
HTqMbF7bSgp/wUit07URW31C3fwYLee8vWW/W7ZdHl7peCIu+w3IBX8gN900IgAvT1pjc66iTqkn
wpwTB4szQvqHqmzkyFZDUb6g+XvwYi2bMi7kMpi3W54f1+UZuBS2/qgMlJGfkA4N4TquCdevr0zl
ywhRe2FGn9/pqWmJE0Es0K8n0nP8gUnEyA/tTkDgGObYnLn/iVSJ5abF2QJ0nDDRWNbdLW5zzb29
j+2bM60x6Bc4ZpOZdQrVmEL8VnteAJjluL7hhwEM8X73b+XzTHZkbfdg6OIDW7IhFRPaNpjbhH44
J8vzO9tZyZAyIgbi7Qo7VWp/ACkvcfTGlfv9rLi8Pn/n49RpiDbIvKJBujZASKht7eMZGJbpIhHI
PyDu+7tUwCgGG/HlPi7wMQkzvBuuXOPmfKRG6QY7i2ir0pWk1W7Y/u0KEp6k7V1pSTj41LFvPH5r
ApVPVsIkaz8c5Z0FH3UXavTnWCUKb+yO65Wqem1AeIw2yHJXNyRfTQ1SMrDfCy12C8U6A+HpXkg/
MdaHroqLoKSMDP8JzKaam8p0n1QYwTRo9z8yofHL65ik8O7dBzagzcRp+BdX97apdSLbWzFrqa4g
Mize2vbCd6FT2WJfqcVIAvBi7KtNRP7QzKJfkn9HJNaMyZx5nK0gukKogLkw0WwQOysq300iUmuD
4OX6O01jSW0+J5LIJeg3pVXB0xq88Do8c/rWQsILZvwp8XoDA2s8sAWwrQIuxMYNKhJW5ixcpTJ/
3KPkobUDNEnSO+NF2dCVW8UU5V6koW9sefLB8vd23m3mLkjp3F5KrXds3N8eD8PaswOHWLkRWU7y
3TdE13mixPYacMWhI1UwkShkkP2lNRUF17/x6PVEGSM3Bn1sCtm0oCejZVEJys9titIjTXmvHJWi
DAOo4/x/TfSbC7LcCZ6dtazeg3SCkc0GYACuDLzdVb95p3P5ema5eDup61a7hn8XoOc/TbwciCXe
ZU43etpxINdr7WdNL/pBQOFZO08oFYiuQF+2WVx75tUn6RI/l4FRVf7ps6CpmFskXCYhqko0QhRH
KZz7PzXEwQq1I3WPeiWylYeGu4FRNxLmaAh4zLCo3IPfib9tY1jWCeQJVUEuuwfhHxVXsWGI1J3B
nVoQ9Amj7cxZ/fMYxmgZptXw42kGv+Snm7TYuEM0no+nmoZ+nXOLsNMYkwibwE5ir0HfbPl/NOxt
4Bb1ydQFPmyxUi7rgQUn2ZtubakimH8pT204nvSYjf4EvwY96YPMKGnf30QRs1ZRGkHNLVDVwB6W
sOLPMQGowFlmmOKpy5ym8IiMQQvB7gmPfIND+9yCgqpbS2HSKjIo1AmMUNipzxifBOpnDEGMNwHq
XU2EpzyFKuxLYX73hDyEe0j/T7To3A0MoyFxcE7K2R0eFJmOVS5jQFH/BJWr7tsxjQeG0fEn9wnS
nonEnL77FQML1LdNalapALXFiwSCD3NG/SCSq2eMzodrqMh61OO2MpMTdrt5Cf1fK8kRjt+9mSH8
E2dAJE1ZUex8vsiD/wK/6XcRnMPsk6cUQPSIbSTRJOwIslaTVWTJZOHEtYC/48iYwsLjitsunPlc
eeFGPAaVEPjV+9FU/JxfQKV1ar806TQ/+tozIdribgz07/IBMJWvWmId0sMc4f+DwmtbKT/NsMsB
0FqUU2wYRxwTQlwianteD4UHmJiwTttQ5wUV7DKzsTRtbVkvM2N6oRuYr9cspKA1Qnw3aGzXmibB
No/pjlHE3u8e7cXdwn8SDUfQj630dRlzwGdLc+Spjz5rtzFUTYj9oWIm+g2jk1aQB7aGZMr//Z63
kwQoIv0R8K3p7lakOF99KMM9BVyUesmsWBJgXcfumkzjgcfaeCoQ7mK9Li2R+VrH8S/gn3KtBZP3
vH8OYmwKpDjhRGQyjPze4lOnoWmlglxFc/8n7tcvcPvkqaVlHHoz26NCEk5klxo5/eaIcVHKReLA
lQ/dzEPCSeYmYujnvXzLmbVwkmWTbEXs1EUGUm04aktRiq02ZH/yfWHHuO4by0O98594uWwfAbi5
ScGxEy/x91/jrDaJYA7ouNMtvju3pGFXPxp3LDIUopJgzrwasASyL3LNfmx+YQ9ZL3UC1nmSwQNf
sE8uTaI2aVr1/VljkjpDgup+ksBolSfARxBVah3B8uF5R4hyN83a8EO5GIbXYfkR7YC4/M6EptIW
fzfSl+gE+E48Z+NJ6COuvtLX6G3SjPvmyJiKQZuAH0p4/nH9kVBZWgHP1RCAgP3fSZ+C+EXVhVxu
30i+xY/J1LGw4UucHgXi1TWKGsaLgOEul1Je1R0ZEPY+6Q0rcVEc1ojv0TsjClCxX5b4xmdEMTlN
pXKxZ6N0vcnRWyg0JvH5f9Kgx0ZJ3nOgq6Up6ElHoPnzSO5Bww4Btrrj6U1fBvtsOfu2ojC0+kkY
Xhb+HgB7s2lx442JJmrdc6hCsN7kCBvVJ5044ovFReo2uaecRC2eQExe6Zk2vLgwRJcYbwHkPcTE
PgbdSZ922GaMEoEF40N4kaglJEfQ0zK/dztY8rP6C3TQi5vEOqG/CNmi4Xsiv9S85ox7mJS5s4dV
FMrT9L8spEba0haT6tlRvsEdEoRnJZGeLsr1Xb7CPvwADim+vDE2t3MjhH/xPyEMNNX+sLUkcCHk
zTuBlJtW+LKmh33dimEPgzAKzZP+6qdVTPTiRVIfA6Jl2rNoyJp9b9YVU288/hNb9PFfZMUyY50O
na4CU49CwR2Z5/shjTCGgILUXRcLwCkKbYUKbY+jpmJZyJCwirWcAernWeAfEyH93b+P2gNbCZUb
IXnnIdOnX6nYntK82S5NS0hyBQpN+0W+OTUwoIlETYxRie3TR6WqyCP5IeH5bGR2vMFUQfwhM1hM
HaueNZAiZ0RsebisMbvl12Xb8RpENZFPPqAadXUNTUWmRdixHNJLR5jzDJ6EjMCeSNKC/Kt221YY
f5WiDfJQqSA9a5RQ5ftCY9gS8bMBie273C7zDecYf4+QSc/Ga72xZw5PHOCWkJp2feSoc61M4E1G
k7MGSWgOnvxuLJt339BGTytLXDsj70GwjR9DHZKau9tFPMyBw0I9vmrtNd8oHFHChymFOAQQBdlc
r03uVcRjwXAjHE77B8v7hXxxXbdDbx/C40P6YG2i5h37PckXmQQ4exfX+yg7xx292UD34zjnhBD8
Gpz/f3tUIFvLRUyhTRzHIg5eZ/gpaGHCofWjpezkxv/PSyEftE5GZW0yN8d+9//HbQhAfD5yte/H
tQ0QNQqThD14YJUIjpO/0lVA8Cjb9HbZDmsVEQoinCjJWblvMNeoQAuB0PHBwizSOLDWB/E91zSp
xCS564Kq0kGcs7Nu2XpQGJuQXe4qm23kTDi/Aky4GTf9ss7SxrxdHwj+2iBRKQJ6Kmoelz/fs46f
I9cTrbADxCpr5d20pWCtDrQl4SOeBGviiaO+kJbQzN7kmcZcI5jtm/N7t1Kr5+ib3BjElGd1i6Vd
vqXow1r6Un8xy8Q/jQQGKUOMSeyUEFz1FN15FAbpWPUWiI3SKL6fm1+PM9aqsXYbGA/+KA0HrWf8
/mgiI03xAhqBsVncG7uYzNsV7f5XmcJZYAtfdFUUAX2heoFN+V31mPDy/yVg/kk0TfOE5P5uGv91
7uXkyCJSdbv40irSzS5wiyURQBbRufkIgUd3b5nuZiccJ1CVaQ1/iUhFiNJhWtUkqSTz+OhG6+bc
WpaCfCNlctYj0RX/bQeMhpa7qxzhfZefBDNKzYw7mVmTbzfxzoCw9TuSXzGKOQlk2DHEjA5Aqy2d
aoWgj16VE68o1YT8aThd6bph3uEOzJ0HkN2tdh40+3fZNrvioZXbVQmrLFGhbjSwcw8PST4ldDAb
6XNAvgXubCswb/4LUusUnl2sm/eH/HxiI5KsT2wDVUHRBvQRclu6vSaxhs8xKc+gfQqo+l3kSw4D
UQrdFyF/JfyHOm1efruoEQz1wvaMfImqSE7NFTBXVWsvxorTBAXpMElHj9rRirQgKaU3kPO3q1Bp
mfBVL5J+R1G3OvSVqQ7PYP08FUSqECQbAKFHC9K4ZpMNvFQ6uFdFYyXREEFZ01bNawLOiXEf7rLe
Szb4Vv5V0iAK4xdfqQzQcDpknoy5z5MOloupZNt7t6arn4gg3I697Pyp31n1IUrg9ETmyVwA2buw
4jmzxAYkXYF/lsfUJdK+d05i1YDb0zVciyEsg4sbbAEOz/V+TWYpUA5n9mhzt9g24Y3HLkeeZyvQ
9Ll16gK3Biew/kCPThP+1TIAff2Krz00gNbdS3XX/T4W0BYMN2c1sz2cU7WPTroWsWYYLQzcEPLZ
d50oejCq9Aw2WNofVqeCMwdRvxjSOTUq7LKR6M1pVT6lSXfJkehMaQOrKfsnueEJxM9NjQh8fM3Y
OL++WF0i1NBpGsPspRXxkBKLaADzRQSz9EBQUcjJMo64roeNBUSo4zyf6eYBUnfbJi/vZwAcTbvP
fOaQcgpZ71+ntR0y9vBWfQXGL3RqBZ1rKtjCRdZXccUc4TdzdI+79abT2Mr6PhJKS4eeSCgvcb2f
ZF8Iwy98P76gF/MvwB1VaMcCaSHp7mCP+sIgwE6Igllhzxfm52qnBEKYoOadPq/FF/SA583Y38HB
zeOvDWYH8YM2LdTwg4AwKCGcpT6TBJWhaXftxW7OOojHVEeiUm5es7kyFI8A1k7XLaR6ladl+9WZ
XkHp3c2VnBo0skKDll9Y3D7R+Gp2ThrTXwNkOhKIR6m3aJT4ycDIr2gNSxIQ5MSk7+jQUmN8c3YV
5HYQyV4F902mo12uXDCNavxeij8pZUYLge0q5Q/dch01Ym77cKek1TdoLBUQmhW+ks44uJZbFC/H
qNJGfqr+7XKIJh7jguDC9xNumDzrJfBaO6/BtHPimzeRwPO2vu0TImXSFy/QPT84J3JYvqpxA+t4
uvLLKsZ4SxQAHua2Qy3eGy3ea5sJEtVgJT+6yFT/tUdxsxVcC7FhBkDNaQonnf5IbOF3/pFlqk+K
gcvvQXrD3Ub7HZQcwu8GcIY6AO+NxfQVpVVeSInpCG0Fd0baq5eZcvBWSgIIwrePFtu8pxdIG3zc
O+lFXm0IaFMlWMla6QJr6RyyUxHZJUlwb9VaU5OBJYxUVconlmKCS0HvfIwMce0Mir53Xd5FvHN0
zA/zGV6jbVkQSpeBc+hhlSQDZ7ADyphtlcVoSd1JSvtJ2yVE4mt+MCCRVseACj3YWlKSaDs1AKsq
QpsQdMexgja0KnBQm4EqwTk6GU8AsmEbNJC9g0xUE6gNqG3fFlLuCxVYTiagI61bcxWE4knd9DcR
7dTo/APgYxlCHgqaSoFMCEyk1mJxZ1sLqkHfUtx87ITcK1RX1Zs/o4bLwzop6y1g+v9apl3Xsset
NuUYvA6285dwauZVnmtoz5sgBw3w8lS56ixSPnSNLxnOx2Ra/mMWchZY8YPRzI82ZdiyEfFRWO7/
uvusdgR6qournVfnB/LXUHn7BqI2X07BgV5ab5KezYBPet4Q4ZMIYI9lvxJQhAtMCcTBSEodhm4y
Ilh8fHyQdmsMvmu3uvkSnZr8qoPXA45Np7cU3SA9G1sdPfvqkgdirAAKxsilrJqtnmWbQj+dALSl
VjtFbdP4EqB2xuqmmoorACvcXqoHB22os3lir8bOBJYsz6Ke1OY6Khk0b2Laz9TERDh7v4zmrvc1
P8Ul6BXvhgFGtlGn0BVs2oCL+FjxtR1NGmMmQUJ7Hs/vHjK6lscJr7F53b8G8o0KXK+3MDpJeU1y
Zss6OZ17qJuoj5nsXAWbLHmb6aQkwbKCVMFFCHyMLk9w3qvgu70d7G4XZZPnDkTOEww8CdvP/gnN
Nr/qtmmL5ASLZMCR9DZ5qC3cmviVHW5xK2H9onjFpiCbLx0XLLnT0iy44Kmg11d8qmNbkEntQuxz
HiBl19Rs8eeVutLu5s1GgTAnvEDzjoS3WJ/EO8sFdybyXaY8r1MC+qCOgX/1IRoCJC8xlrt2MRax
asjM6fi5QCrhfW9V65Y45DwQuoKfhq4TDj+b8U4rf1e9yrkC7GoEolqAm7Hu9VM3P02LMOBj13Mr
o8o0DJBFGjDpoM3IZgB18RXnhXL1S5DlkvLj0/DqrMA4pj1cDV//OJktRx+dSrXSBpnJHaQom1ph
9vIK9Kkobs+rf/QqsShEmxYTZt5R8HTVQf5untGCjpzD3U3yDB5GkdLTrMQRj02H/nhkFFtjRfEB
j9xBxLJqrLWpj+84Sx3FTZCK2HnOP0DcRbvKiYpBoMxl0krk/nbYJT9FggpKaYuU2YO7ZwbUB++m
D90ygMJHv+TAt7DlzKaN/4YmjNFehGUcFFXlyRGQMLQQYfu6ApsbRjmHvIlz+up75XQ4aQx9TkIB
l7B8RKZMFpLvVys/Rq4zSwFvRTgZu0zNJP+Mjs1PTDiiLzI6bUCYAjH1p+Zre3lzEC0zjtPpyV3B
zSl6hFaPOBNQ4GlFGJ8ThfLcLt7EjdqAZ173lSH8VDY+p+SJscHNx+mOINZ8ydBamB733SvHeRbf
EPUgi/V/VsUxXGpcnpRNTa4K+hge96Jm2/7N/GOuQ9LrqdiUddhbRV/Fufqsnv02phIriDgSZ/i1
YESg79jPdeW5GL0C7h4tpLkIF7EGb+8l6Ys+bq6UumFoWa5dEStIurQPIiLpin3LkfFidYlIIrHo
b7QBvQIjdvexsPxcPA/BAcnDRDYJ6canvGeRRkWCPLDMc/f3iGth85uuwwreqYBNgUf3PWbBH/p4
QONEMmYwWfDqdRpNXvrXQ8bdOxyApatPqs7tckPCogftjTIZVd0UXfIPbEHpQULHklckg07sAzTx
qXPkoxpeoXxd0CFBy7VBK8hddsKEU+s0JwcB/ZEjY8WT1gOaUGnYa0yar0Msq7RJmhLB66lNz/wE
Uw7LOBMShUXHQxz4kU9/sWiICpOrksskmyUQx/KA4BvBeWkehHWNsTvv7mH36ZA8MpGOY10zma0m
aMM9SpmXiLch9Ch7bzOH7Po79XkU3vNvYEV/BeCXl5VXH5TSWVqzelN8WqfupyMC6nI/fR+OqLK7
QGX3NP55j8jtImA0VrIC1cXlr4cLkSlhhWDR50qKcqEst2lLZKQkpo3hecs0bDFKyi8dJm2IyFCp
bQMj7xCaXKIgq4fRE7N6DNK6wjCqTM96ui/cXGKPnq45hbrfgnH/KJnt9m+KMVhW3yYxqkGLZE/q
DnYFu2xtwKIJQ14tNuf6D45FbNAqT6y+ILaEvyPY8VvE1oGYdK46sYJcCuS5mNxpxPa35UEyDzwk
sraczWxdIdgjFDthG5EOmiG7G/hMfKCue64lK52eZeDpEnhS4EQZYH21K4Cr51FeQhDns92K5TqB
oxxEtXfwbd9Fhz7dsVlemx9E4MSKrBLClh4hDpHyGvO3SWpLYjfkX0R/1cIOonlzYUjKF5X6Sxeb
TWMBhOQW2R9XsHvaGwlXx9km3LkAILe9JOQpf0DRgAUzhQY/18td2AsFKvp1/Xi5NbAZa+fsGnOp
faDAEmhahIlKLyqSuQT3lRPXkw3qXZHA6pzr6KfH1TYhtFjnDspiNAhnuYuRE3otlbbLUVaqKNQ7
PVkJ8+3bTn58ysRF+fgArsa8K+JSGtQ7rtQh0Zq2P0YpyY68vdJwTck+y9EqZNB07uRz39m4Owj1
uGXoRNYPXJ9QJLyWDoAEJDgGNfRLUJejbEDZYOcqV1JRIot8RIqi3Hkdo3EEGfALpWZzN11VBTMn
YGRs4Ps/FxKqhBo+gg47/YI2HQY0OvALL0H9tT9KAaruhYFVnlb2zd4ogxQYr+Thn0A8iZTpxZwG
CNES1DzhDXWiFWm3jTd1OgQgxl1uQXtUo7qpoV09LD9dYqKa7XocDDz6EnSGAKz2PXRU54zd0YdG
GQxE3UCrwXe8WVB+T7Mh4XNo1x8tbWFofyfgG+xQ/3CLSiLgM8gn5/2oF+9NAzQf4WRzZGLGUFQa
3rS7MZDH/ZfUNioLMfj3ln22ZXveRo3K3z4XxPeflFbUpp1P1yMQzKlQn4TOwVF8ENr/2E2q0yx9
75v6g4doFCwjYQ/dWbxwZoAdGOijFkAEvv4JH11ojUdQQ8IXsAraXPKWWMFRo/8xAwc0ambvIY6s
/QvUPB5MdYqaivP/ZxMlIjaA2WsYf9z4WG+8N+sNCx+hzw3hicGOUXj2jCKKqXH57S1TAzSusvlb
7OBRtHYErZjvgw5id1wRboUE+nB1w3TvUZEVzq5deLVtWMDJDO/DINc/n8/oKWLQbtbmK9iJU8sX
XFUNgiFrWLtdbipWeCfFVPslTLEN0tmM702mReepuNLh1UutkPqq0N7HTvLzSj7sZkahC/MwUzCk
a0/e75/BSe1eZiX8UR0OWldHMytzvAKAQCgeoJ7STzfr5QAz2vecSoJf0B2+Cput5K2lwnGaxEhD
vRkSPAgaQrHxBtL5XaDfnOu/keSZaHJbX3r3CnEUj1xw2Qb07XIpUxlcqy7T/XjWWDwzsR7nI3Ep
xlpX8Ztlb1b6Tr7jofuNOBRE2PXWEb6KJw+Cs4otAXVM47YVWBUvMfvW/R/IXpCnrFO0/cTicaI0
OPge12qmlM1Z0Gg1jzI701yA5xrQ/u+YrFhhWJAU6TQDBul6rJA9NQYGsg7Z02dw8SWLfwIXMHLa
GQKSqN+HktcFCSZ9+hTQz3AGRPHmd7pC4dcSk6PnVFO0opc/3VPnN528ZypL+VI5EHlEULpNvebc
YNzbaA9vPFldsTDPMMXw84TMCxyxn2TRCPcbjUfDSyCjj0aS5OuhTPfTj+H1wHjvdmzZSEOmTb89
pq5sBtEcorm1Uzi6PxFOufIVM2IlfOZHXaNtynM76fkREBHTjo2wHPx9MNRiqIF2OgeuT2s6bxlQ
6FK9gpXn1ObSrRKdAMpzGWjcCfKKrwesjN6t6moPehjE7wRAWuT89/AtJ9Tg8FjdpEZhBiSbZ5Rk
kf7MJ2uPiVErt+SZoNMX7k2oAExdi3sVKAka3JqZiPtXgLx+8l/ThvQHKXU1TNiFwUKzoj76Aby5
76AxiOG1jrZjeeYtC1ag+SXEyIIwBNPuLvW0v22xbNoccE6tasMWqdjMnHxoLvqTkB2cbZW1vj4j
J58EpoDmNpdC+8rT4SnkggGVR7GuoGInBgXDYW1Swu5/XMjmwGHjo4tCbdXzloLfSfmGybiNkrVr
Nx6uDXYh9NCbbq2jUVgIcqhV4FPf2uQCqSpGjDmK0/oIkS7zqiGOtnESqWviPeC0Ryq2ShDsGHSw
AhLFV+4dB6u51QO+WhSl9BP1iHMDuAxhQxKWaydzQQCjbCzjiZbocedvtVScmlMDU4e+jx6FFPwP
ISAleb6O5eFWzeLaR3v94l09/v51KAuyzkC3wWjvuY1KQx70aSLFfZce8EluOd8eWpbAiNSbYUt7
TY4Xj2ay+/6WN1PNdN8r4W3SNcwnGqOY4r4qNTyBaO22Sp9GRMvGmEaGs4VdvDyDfbUDfiYHQ+1Y
aJfMGc8BQRrTKjphZrHTXC8brLGI/j1HSfSfB/oQaFMBiub7mLGQZTQKjBKXGG7d0jLTvxSnIotJ
oZ9pMSCnLwUKrizl/kVAoq1pWWb2xRqvovqvAo83MOBRqulXIPPA+nZuTb5mCG37/cccdAIHDNwS
D7PAXsgsl5UDE13Fy4m5mgITmVdHgOpwMeZS3xERVYOLHjnIB+/hx1RCDyK93XCrMCWvAQCmOKw4
bt+UWttbIvgOgzvfGPltH5Hog1mtYdod2X0HCXpwaub3IJfeIVfTWVgh6Z/cEmECpFcg2mGVkC84
BAjyoOdGReEHr9UTPAZXSrKWeJy4Lyn+oEEs18OYkMr3RcZfFPtQ4d6fP88etDBzBpEtQUvHGfs8
2RT8gRn2Hu9itMfhOqMh8QWbtXHpPiNkT5N5u6u8hrs5bgqwOJe+l7QLxsuLuVPFNBpNI7AG5V7l
ZegmfCra7L2s8lhmnpHZjnohzUx7BnUQJ/akoDSJ97L/L/NTnrYHQxE0ybxcSBd/wsyE6goTOTaS
HUuxT7dHPaskfF0PaPs850fc/rCrOyEn3XY1kD5DxiHkR07cZFiyMDDcsqv81v5wJRapwIG+ZvkP
mvHE0KVoZUGexO5YKUNHF5TXGHCRO1t5ALoieQlXljfYIMJhr+2WiuWy459cE+0WiNXROc+HYSNH
NK/9oc3eavheAbr8bDAYwnYwswTvcTjDC+sOYUjHHZAjVoVszJwiBPh1EWYulj7+sylcScbeNWK0
MDu1z34XElYr6nqLYS4EXGBu8tYR4bnCnn3UvGFO21R9ds+UMXUpMQagZEo5K3dUCJQhCY02UC+u
7ueFyHDriz9U7S5apLmn9cwAiH9MpG75llNOJUmAY1O5W7oO4N1T/hLW3ojCYTP2zMNWcnPNyw6h
rYEL1SLcwCLR0UOc7b31Myak9/YEWNzyoW4eOwqZbWAZFG/gL9wZ7nMIdVK/0TYEhQRTkteC6a/v
6SEHhPMJEdBevCZXsCgXX7cEyw0zKo1P/WpDHTcdoMb64qY5O2899vaOmIQpyjzWR/yAzpsSH72f
89eSifns+CPsMArBVkTuwBRCMDDFRbxmKUwTkwHJ4JvuNvP5NJRkk2hTdy2tT14U0vtLFQZD17IJ
ce/EiMQFoqtDW/+7xAj44arn2naTO/MKh9G6DHchB95q2ezgh+E0B9It7g903JUkwfHPcL3YJxwR
5FJ+h8B/A++ne+xPWGEeUdrBx6daOFYxwYLvnsinDj18FFsPho3FFIYXaN/V6IjoCyJEf8SbxY5a
fMeYb4lhiEBH+9yMBEuI9Paig2rNO+ePzpbDkECqgUJjF15bI6TnAr7Fxxh/kno+fPKS8lVLrpOp
YasJxVi4DpB/m/NgKcNupOyl2NP1GGdFNPyMgUcQ5dCU4QrReu/poVM6gK+qfUQLQ1hyHjpUtJ2V
azJC3wVPoT78oukCO476QSEfNjxPo2nZeMXMHx2mySOHCpOzYX53AYNQWVEKeaIHfrWFf7iwHnqt
xLwn9GI6P6BuWI3ribRAMaGcwgSi/jy/Y3uxOv9sJj8DOI4xNd9kfVa+z4jT8mTHuS6VRQNWcR/d
iqAVLjT8alnSZtN4mLKzTM9gnr07WwMzRtkBoj/84Btb1LBqaWdwWRCzs3dFZggLvBwraL3C0SoD
Bq5CdaWbptvj7E21BoEPatlkL6clX/0upnl3XlC5yPWKXsMYyh9NekEMLEUrpRZB0nIgvxYjYlja
tbGq0wYG1rmKqjjN+955QBTQIGMC8/xxWD1Yi3l6QmuL3g7sCZ8vDN2W/lflGQ/nZHrbC9ZTLaND
snpnIhY3kggI5ggibN0eWQu03w4vZTKpgT3RUcaRJYvgdsrfSZ8JtfSHgkggCLKUTBNBSTV05LWm
ktmENqVb/VwVSw8oSN6reG9u56gR+VkHXmoIegsOYj1s8wjWAfDMxMXpPMYCO0joQdt78jEW6IpX
iWNh+oNDdYWnB9hcBXUVrlgQG9PfX7hhayUfLW71aB2c3kuu9CDu9h2KSBNKSytbOa18trnqCs4+
xIQN+xUF6PPOZbtGvqPVlbeQTtfaM0CwC7HaP+jH943ll71tjRz7hBdbkWuPBzOGQ4ut6ISLqI3W
S0QqudwCb7vYlxpcNC2MXY3kupbyqq4LIgqkxmK5qKWSHOrFCFsFcv63n6llWd4dGXA0r90DqZDA
rnlx+S0Mqiw6zRlOR72a8820ZCfqgGUgA77xRmlV4U6SaH+6StUrCNn/CkjvDAbyh2H/fxAUVO4B
QcKWhP5qhZLT4HLdhpc4qELb7R5GDrclvGZwwvAn2lCZrGqjBwGPflKwg26ShexjtIDgnd64FfVb
mbTH6Lif69RyICYEz6dE9nXxTRYQ0cCO+UvhSO9OVGPphIArfuhv+CT/rFv+MxTUkqPdOCeFYErJ
Fi5OFWGyQCPh1eXpIs7qJ73jdxBLepxROdMWn7BRbWd62GsXUSjJaeAkUiPHh0RlKUEzGLfkY6Zb
rYVBn3o1eXWgTR86+d+gZFPQCtZKPmarP0xKpOKINLYtbtdgbQE9bzsoKO1EG/OBQ1OQ6Iqv/fHz
K2crzZXe01ZJMH7xT5Ghv3r0gRX3mSbHvrTHmIfAbVu2Agh/26E5Hw8XYUCPB/q1psL9HzfdWO8k
cIug9bIMvPuM2YvNau5AMamz76foHajdd8wyIIePLQGWuq58lxgVgXALlYI8Y5g2NEu6TceyvgRe
HMsBb2zjJoKtdy9wZAMI96ShMwMuP73Tu4Ovt0b6GVF4+JvaHC9/P+HQxLwfJppg98OZEiEtQPGf
5Mp4a97XRe81XjCwrElppMKxV50d48gnYrvMfRjI5pqs7+T7uaAl4VWjwWsNWhcdh07hIC7gsKKA
QVxSR0j3ThkltEksO7vZDCzyKNFsTVZqLou+RtsGwMHIL2kJQxZLvWwL6gxHeuS5X++BYxndQsm0
qQ3fZq7VzLpjZxLDS9AyiEicmQ9wbrox5+a7r8WbpiA/Xv68cjruzq+Nk1g6i1nBfJ/woBb5ie+c
sYn/4riTHgDSXvSGfSZxtkDqAXoToC9OXu6o3gz6Rhvab3Cwr2aSQginaQMjkVgDQFri4R6o0xQz
ORWdv+m7DEgTpuGbmzhNflC7MrX7qpdDF6AHA+AFGgOKUOfqupvH3PE4F9JqXzZFTh3E1G03z8cb
t+K43GRzf1ALO7ijDtU5jtzgzfyEQ/ei4TGJkagWe7KrD/cyIqVzlE3EGIEguVZzHUSCodZf4+1P
TasqfSlSRLT5fkhOlZGutZzcfzKIfw5O5wL1qnnDtSJ2Z9xjpUxcvM93WqLM34jG5dVZzaiZl5df
Z+Bfrp2KIiMvYhZvAzDBYoM2ZRaAFi8pXgSwmpcmrzYw1gJMhOgyla8kMwyKC1mhieSwwS0rsQss
Ib0/YinnLoA5wkKtePxsoBVvbdNHsSh5PTymgLqunp0RdOeUaeFrdatc3WOeTBVxoP0j3z3njoTu
+4Ky4HdAhwqWNCOv6QMdarKIC4lhDPKvLPLVzf+lXrf0oRQ21A9/1/bSxXMPJJKSiA9BBXQQD7yk
f1X7grQl6gfdcczaoXXIyDt4s3CgU1M13inTuupE1KOEJnwCRWvzWYuhO8DKhl6nAHoh2oSdPK5W
h/aAKAU76omIObZsN3J1LKYrRZYCY0TNQ6oV4nF2karK5gIqDW8Q3PeUr2Ul75nfAGf36ZSfNxAR
54heVXGemU1xqeU2OTcrfoq+97UXtoypUnEf6hv9FBZlZQXe7fPy3pJIojNVVpSolwmQbV6OkgI8
G6YCxbhDuEc22ih6HuyqeEXgowhE/r/DYQ7BYBw9ujQuSoaziR6Xj0DDpP+HwmuNZVa9qlL/tU1J
+pdo+3CDSp2n/NkZfWlHLazW3gwBxg8bQJ8sYzl6LRmUP3wV0iZNoJb8Fexur/CtBTfeMf6igwKr
jy/rA5PJdgAcQHAWtpgIcqfQqhML6admqHOsOPFapLN25d4XCCvg+ChIbQbQG3jpbiwr+FtCqPRB
vUpLtt5rdfY0U2fHulgTYp1Z5kngddQ/kHGL14/nzTIabOqaTPMjesF327xFA9JsXLZgKyf9DKEH
25mhv/jJCRd/b5s5z+7gIXKVpjWfsrvsmM452jO6/ZXsqk6937ObZ/yYpE6dg75OtxKLm6T0wFYu
byHpFFHx/00w4hW2R5wKEpzF8Pvz86PhcDsFZn7lret3YfS9wv8Z1BRoUX4zGRg6/lBKV+6u764i
TBeJi7U+aZLsjPR0XLg5orQSQF4TCspKOpjkYjLI1sB7rdoTjYmpYEO2hlHIo0s+9mYjetuvKnvL
oGi/raPmay/Y4JC1vrR5eZml89X4pKwH8XTMn6npHzhKxuheEikfc2lpziypwLtBOKH/Sdd66izA
pDpoBFLMAEUiiP5z8SVmrJb/PH6O+Khzieq3lRBiptm+D8q2/qeAluS5s/+jG8PhPRkGSHwiJ06T
YyPLNOmLcmPjuGY0jHSRjqM+m9ydIZt/o+VSivzt/Qv5fF//MXWGJTsP0k00/Lh9HOHAC0f3Rys9
CQ41Zp9pguIsTB1qfNuxHnfGjWifHZDQl3jTkOJWggq9oSEQTfoQUcQPZSSDYfp/4Uo48MzOHCfv
yYgim6YNBeTTcY/nB8HiKyp0Q9RY1o48DuPHU7FY3dlv82tEvkUClSJ5as457atDC+algoCS2+xf
B8AhGNqTLE7bXRMOJItIHzUokON5nhk5EJV8pqyxn3R6TfdJDUSwqRqkiUFwb2TF97gLAKFoh+9H
VJviP4538VRYf2WuLVi22rE5Cu8UrNDOsybq8Fl9VBMNGSsZ1KYS9RCAuCON0S6RKjxf9SPDp509
7oSJOePCv7Cjft0G1B9LHGbI8B+cLrgK5rr3c/oQ6cY53Tudgq0H4MyyzpUwXgG3YN40HfNU41FR
J0iD9VBTvp0ZHp2C1Vx7OiiXVy8kAq0ECdsJg3x7CNSkr2Us+Xh11s9QyA1k0e3I6tVWgLORVRG7
9FiSjfhCWoWnuvuk+Wm53gp4+BXvYOqJ0hG+qS82QmbTszHdbVIEmvWOY6oGAO7G+Q2ZaxZ9BMvX
nuuXSwMJe9UPFV7TIePDcakodPq/JK/dYDZDe8kXB0hMVRD5Upija/xmh3XufWGVtQmUN2Xh2K1c
wjP1HkUFZ7kJzlz1P8/Do/m7VZxsb3qe/Fqgazh30D7zPG9kkmEuQbBa0ZDnZJIsqvuHcLjhCvOz
eeMdT1G8pjxpu09sDyGt5ivIv9iTYw7sNYlhRLf9Cw8sI8/WIlNLB0UggjMJmR4agq+9QV+5IDVy
VYR89CqHRpE7vzj7uW7n2K+Lbo5IcbKhwFEFBXjTMp4clXoPjMQtHPzgnqkw6kioigYqdm4SAnJU
rbvqbELMudYemNXtbE2PJ0K+8kJscRM2mshRz6c3GpqAB9v+6DxY8NckluvSCa/EdCiRQhA6P9nR
ACdhRGZfZ+SQTw8uuSPuJlhE5GIf1QqN5YjKs2VR6xuW8HFGnNx2Tyr5HkJ7mqYhoJH5y0HmGUUS
IAuh6A0s6kFGhD7xMxcO5conPetCTjq6Z1BuQERhL5k/fClt5icdDOrkTKozVDIlRJrwEODlwOWG
22TTou0YykzbT37Aa7D6hVkaGsQXLzfZ8TQfN9k6M8uSzf3B/2zBPzAmkvPS3SQ8GxUUPSIGDOXl
anEFtHAdKtOIn9xa4kC+v2p0tEf0qRYX/MBqgkNHzqoYeZwE+0oaykj8NfFivnA0GxLv7EvbB+uc
EijFMZ6U2Kn14QvS6xZsA1Yuyox51OulHcmsMY73XhsMO5uwaPCZAF+crjvzTg8zQLFCzneUAovP
pIvgM1su6n1oJERwh5xr7Fyy2INISy5jmhRgsb8kFahNqh4jibLnGW+Lx3ufX6rjK+Jzr1ujj+YA
GTDcwArkfSGox1TbpRzS6aiOwM6E8ZbPKO3TF0JHaR4eJSbTTpGYU8OpoxKwwrB5e77sydM6da3B
oU4Xu8QJ9lm1l20H92LTpJTsxafX0Zp8e0Pucb88O5Sdo65iBoDACh57gCS+FnE8ur15+936xs86
23wrwEhDcLj9MKfBl6TlfLCSozLCsq2f5zKpVggSWVFmtm60zA2kKSskv1okMPfpm3+FBkqseLAq
WDFJ3qeZtfDV387tFlSVm9cL6ubyP2Qyb1yKsq2quJKrns23vVXzUjcf6FrTPyS4R5mAZF4fGl2M
k5UiogtyobePs1g+O95lf9RgC93tzGWI3lzu2fTVQSsDr0hko7Kg0qisiDOS3D+XjJgy69pTRHwl
8CC2G0R+XvGfkrPEyq+tSCJz/Ec/dbZVq9y6iXIaY7+JWdoV9+Kw0/QbZ3EtBymZCcHxFJkTpoV/
/tpausCV0qTjii9yW0zwADx7Ph7Ur8nPe6CpKT0/pZ3W56DbwwZEU7WyjkAyh6EJSuUmWGhdZ2qA
6iN3viF5gb7RQ2IZhj5eyB6w5vo7+F4jv1SmQE7And6RGdorgA1O+uLt1x96QHgz5gTIGZb/QXdx
7NQzHo2+sY5s+1vviA5XN5p8wbPoBLo/2kIDp+PfGVPQBosBKN9htdF9OOoJ2J3P6F535KFm1GHh
PnWXUADtqMz85f0Jf26sANohS/Ey0ETf2O+cPIlem+7Xe3MITN3QsxVBMnDvv7bKrlc2OC/rttcR
DxVXjAOFVqwK75VrHFYMTi1hL8psg/8O8Uk+yS1xcW1IqoA5sAdfwkYEQUHyin7jU2kYX5P3y8VH
Iep55JjHKs93UhVJbQnpdqJqQ7t1xs9HqfC7zjhQaH9KnIF3L1DjMyMlbbGnsDu+qelOqF0/OQZt
e9t6SimkGMmINDYExYsPITw63qNAtKvlOB840KLqEqDeuRnpdAZrUA6CNCkDcVCAv/97QnXvniUC
/oPNROaq19U3csG51Z2Q4oan/96AFWy5BEL08w3w8OxDwpHPZSM0smVesxszWKaVgPJB+zGEmBND
95fIwV8XNE9wjKkq+TB5LW/jOdAj0XDAIMyVvduIrr+FP0Hv3kjKWRHHTDBRkwsyclX0Brix3VLV
BZlWJocCHAomE4b9kxND0rh4V7QylhPvYaJf9sBIAFDmMq1YudbLKJpThuMWQh9RnREPFX9Ffqy3
QpCqWh/zTHISPYiBaNil/8bNZVbWMIXqh6DcE3w10xEwa4ajzb3NeITYj83JS/nm77ifkDLxEf63
JUMSzm8YA3hHCQIgVrl7AFb16XKAJm8dfyRS4+071zsfR3EdC3tY/CyTaFxK0vscKXvZa6gRdpQk
lRieRm2D+QqFAzRLYJMo/EtAeiwya5NW0ce/cQVb+WzJz1bsHWuHSj+HTvJ14EfipjwOtF9HMpFz
y8RJj4OK1t3aVprkm+c5J5fvhLtDvnLpxESRs7g6k///oOmLg8eaCDyCnArcrJsE9q3DZOGkX3kx
QgTCF5EYdaxQTTxqJYs3oEUWmNXOq8CyNVigiHubAjwI2iDp7XgBniOv8aIwmY0PQNzlJsPUzn+5
zAeXV7GULHe0TWvGtDcfU9tw7xbMJOJBOGviFF6V8riObrwp2Sq9j/p/XPFbyLI1gUu6p7zHO2Ad
Pj9q0HcRqQVNXOa3iBC3qXmoS63MApBSWW7ivvYMzv2jN+c2+RA1mK3JiOE+IuYWLPrP6vlarmXz
l4ZTdQBTO6Y9mb6wTIpnc6MCrf7ob9uAjT7oOm+qqJ+uZUc7fCrzl+RlXxcmyz4P/SGAXpEF+1EY
X3wL+HxbkMWgDwDEaKva3xzb/65lvs1NkN5KUTy/AIP+tNume0w7T/h02eCCp0jHDRJvdG5K1Fbm
mlgDaLgJP7YbjvRsy2ANTQDavciyPj3fy3zKgsfq0QDMr9uV2kWa8vrdP1YOOCdvAlfuzhFqd5Wz
nCZP5981pt0jBPcmQ2YFIzMOCY0rB2Xn3+RUl+CRU27K7UpUB96WqLv5/RDXpeX1coiTlwLIu/AK
WSRwahHQi/KXoga5NfClc/jmQOOCA1ypiPzeSH612Hz4Pv17WXWVQwrYj1ZDjkl+wIEM2d0VMfO9
3Igi6DUnIQGPcMw5HdU0IoNpiVbF3ON1wfDsxUvDUszqaoupf7v60AeKaul/pJsJDTjfiIP5UrDZ
mHcpZJIZF7Q3NHJkoNpxvi23Y7eWCaHk4aYYVtO15sU8gJ8Uyf3gh+Sbh/ymJuDRRjNCz85G6w6H
m1fd4aeuvJgXo2HVtApH/pSSGCntbOGrdTieZ7p6CWeSCQUWTkopNcJvanH+66E2tnonx/avfvZX
mOWxxGxXSBOSXb3hp4WRS7Ramets9ubGviXMYGuTkqn2c1fYSGUtZEiwDIJd5IWKgW7xgjecPbXU
10mDoaqUPgV24EutIQAVvE9H7cxHU227T5OOn3r5nKa50tz1A3zep8d2CJT4iKfXC+KP4IozQdvp
YMAVdtV7KmQv1gcFFeqFxXab0DGGbLs5iZRvjt5hP19Nvdv0lG2Ouu91maCK7WajaNMUK8Y8YEA8
ApsdtG8n7EUFK0Gr014hOvEKR7GRfk3/l3QAQa0W8JuHkkxqNrACnhDtHV9St1cptlpk/cRYK+DO
1/CmyDy4noHOAkNECMOSH/7BgfaDXGxVUTTe+brrj+o/zODoeVhikDAhHxEDIWoHcZHg5fGP/sAS
irnBlyFA9XVqVTvHzpyhrWljUCNAXO7gGCs6YxwoHFb4QwJ2wsxyRZ4/n1x/KVHmHg06jUn91LbH
1/pCvhsuvuItaOutcesfRUVP4Yir+rDrznRmBmIg3HoULFBJkVCOwvkDwRF/qZCUTIMhnlXMvdRA
2uWYhQIsgkKNOdD1NBtLIoImfooJiuaQtsqwHjAwrDe9baOmaD++wp+SCXN1cH08m/UhOX/arAfw
uYJP+erWUE968nkPBGe19T5zOv/cBVwL267ZhFOYJjMYTbN9ckIhZbu/7+UuSrhoGbOlrk3n3N+P
WwZGhTe3Bk1+pUNkpUfz1vWClpD/uJsqvJLBy3V2G8F0gYB7zn+mDIz8dToycZYSrqNFR/HWaFlW
TAywHcRD/5N8gY1EatOYEi3FYR43fFSp7uG2abh2DPkG/L+fFW0ODOzUc6nguRoPS/oFfWKSf8L3
4IYcyc8BKBK4/sTDkjZkxc/3u3WBCEw39HR8B7LDZGhKxWDjT4a3j78j5fI1HIwQF/aG55EBYrhg
N0d/Vdzuak9lHwpbQwEYBCee2aVk/W35R4yDcON9/rfgAj8OGs0GspDwqdsOkrwOEEmJv4LPUDhR
+IFYLO0Cbf/iihPmC+YlHyoDfIOulKGsNXCycf9rO/OjKapoU6cio6t3DMfR7+0SeiG6MzFVGr32
jooFdnEP3S5UqFjlCXIRzfEiVonMrP5ZH0JtpKCeOPdemgav1m6bWpFcl8GXEJppEx+H+PHhF0gK
FKjORgkz4ac6DAnlqsSTIfkz76vJS4UcXee7akAdJWIoeCXtKHzVrrJQ2hUbIO92VJYToZPdBMzp
nKJn3FwAzyVSA7uoq/0TONLnsof8UVqmC4gt6fhn4PfWdcJtWQrsQ6bhqZ67qKNb0qgmd6KbpYhH
jmWhtXHelfrGgF/wrAok685PSfwAVfpeK4W1X5lyEH2qAf0qG6pnOfIUEsRM9tQKj7+sSs/Rn6LW
MlzameDmA2/AeQpD88/mLGjtoNcPBnD1QPXx4wtuZFPLMDYnsKHT6k3G4X0zKWkvNAf+8AuQmu2Z
cL2UAj04B+J9FlYeZ4SEdXg3X4AkA0NtNJ5QStXDWVtfisK4yBaET9D9VCJWDR6bFHpqZokxikim
VWf5UATWA3UNrkz27KfAIt79XsGGr1gtJny8wQfOLF/3qAyr9hrnLK3urC5VbHp4I/K1UVaf1syg
dTrQ/HuIFjX7WXblHVvJXqihLu3R4muSqHNFhAyn+q90h0Xe0YmZoEfG5xBcm5RiaiVovrBF/3Cu
5pcoSuyDHCiLxWi6+Gz+hlHShuIEekCZRLtVNk2jHL3K/98lqGwToFscGgbYLTN693O1k6Zg2xJy
kKIzpXy4pkqAxg/SjyXngKZ5kKZq30DgaZQBe+qP3gZPOX42zNg3HcCjZ8NNklmPQjTzKZdTmtwU
F5Cj4QNIOwMvYvLUEC1ilUCozhD0wKfAYo3BOy8jB17Hi/CUnl2huN0Klfnv3v3NUyKk0moWUMOL
31PrV8hSKn0iOK6QjMunwbuOOoXCH2AnuFlSlc9gyevLXzAdc0evv37feWRRCH/f0P5iHtxOAzkB
LaHNnJunbBWz76PA5aavfnHkOybVZOEhOExQmBEzjQa9ZQy0WitQaEy3mC1m9vm6pIddeP+McbAr
J8/q4wOa7qilj1h8SKuZ/i0ccZr7PtRpf6+c3e6nh2257ZTsfBE5PI7CYdMiyGAEhUHW+9K98ptK
dkMFFyZ7N3CAZmHcL/6cnXCU2x2civRFEZJcl6omXhApj/IMVy3qGzVSYdsH/MROuE0Fn4/TU3SI
yeZk4eLnbr3NUROk0zyBTHgjy5ul2y5t7s0IY+SFwzT5AVdKaVqI0QaY5YkoZBBMhbVr7C+e3pwp
SXeLYrcbtsxpSSdo/QWAlnDTKAQ/Kzn48bo1yZtnW2/pWwg7/oJRVJ5O2d5LK1MhZD45RqIfkEHV
S9kU4JSplHUOEKYc+jaLdeYqcbqIuw3nbRszndNuyE9niUskXtwdaKMgrVsoJO/mLoLYFpkeobZ5
81KBBfsZd5wdpS1FmoOrpjcNJiYIPxdv9y/npf6F3dYOHnaLy1WZcTQfLdUPqyjz4YsOqtq0Szkd
lrmIf9fNR9ogiRyF38TASsfK3Oy02r9psLscaJXfM1AQ8fiAy+QTxSX/9AQE6Q/7dR9BjTBa+XGL
mikVGBbmC4Kv3wPTafh9DcUihPKk1izzUijPCFE0u2K0EATfB2teZDvdXaCKv50awKH2xmkb2bOt
D8iGWiwhdF/3F2Q8kXbwEIF5Tkq/kioWRlUdQa6qFvr27lw+lDOCinnc5lnRiuZ8oFy2ZD1rABBC
1djOTL3SwhXOznjENZ8eSxCGHQ6ycZESBtSBem211+ZQalf8ORXcSzJZh4gd0DYv3AXw2alCZtYV
2jYQJe062WBRAJPTm/7wOS4A/RBT/dITXyfFb+m97dX9iWA9s+OSrAPwIIR8az4HCnhpWo/tAvOR
CtbtOffaigJ0gSYgedAQytbODN98bVDNcx2w3Jnd5RUq9+IqCxRPLTH/Q2Bus2BMkb1X2hQni9q8
w63cp9QefCUk8cpKpt5+8P4aPFE+bHgvU7ljt2qmRLgQ0pDxixcRJ0c+fMj13n8Dna4QH0JoewZn
7+YQGRh4Knm7ut5wlQbjUbFlpJOa17f87vHNiJYNqfoMCE3zll7O61zoR1AvaXDOnpOipJc8YZI7
h3z/A/j3w6DGnkRjZmW/i8LWH8jVQhVfHFozWaYsHuRA0VmzlNJf7d+8p/+z+w6E35oST/Jwe2VJ
wFFCY22ojv7JtOZdO5D31AlSWAhI5sbEwsDNmfws1sBhCt1azNWu6AZafAU37mwSiZ6ek7UX1ZN0
lkODbnXNjMqUZ0h4mbXCQApjIFXmMTbhWDiJlnse3/WdyHdkCGwklYlP7cw3KR88taa1tEXNmjUN
uei1/lb2jY31k1MeavoEd2ARiu/e7RGYOa/4OqXb76ypBfMKrfne/t3HJvxkQgm5Kt3fMxl/mwFh
jpiY64w9+xRrZSTsb9nzy+/3b20IhOzp1414cgj3Jp/Qz2BtX3w3DSi33rSu5X+mxLMxtv/4EfBF
WJZj9yXapT3747MTVdbFwqwbJslvakRChgu1+bFECxADrhSOrUsIUgW56r+Dob56qWVj5IYAvd9w
itKh6HK7yQ+yMxDVKaq/Bp84N9jhfuB7N3EOjCpri/8zKpZbpjK+/je0uCyq5uDpWwZAVfIasEeg
TUIM6l5SVYrtN9y7zwYzMkHpBLq97CSrNGTj61AqrTnwzJHoCovxZtqD4U0QiNXzHRAlFBqEneiw
vEhKBCnPKwOl98tIFxK9mWtbcyOUCJFJCyyxVGhSgM/uHxA48iHI2NMZkhPrY42tt5A7CX2beLMY
5jZY4cUn5zc8Mc/ZIMutBGyb+sJm+Ffr9FDi1IDEdH935TJ6vxp1ozryWaAvFvr993N3gwdMRNNw
OEAJO57N6sDL3sxU9lM5M7bTjYLkvU4avWNHPNZ3rkz1WC3p7JPF49eyg+KE118KPA27Uo8KOIjG
Mz8oXbQrEIsLOoUUm0U4YAZdns7DlCngAW+0MzihZHwBqWgEe8AVlyZwFYy7G/kB964euSeODy8D
J+TznSVOlae3cOtjwvjTbfVXE85jtvHHS1TpFnnxb8EbECrODEDmU91cgVrWgff+gc1ib+q4HGEY
YjlXcOL+83LKfBmWmISDIAEU6eS+kYvw7q3v9VaMn29u9AhnYglqnu0ujFLrHyGNLr0tKmuEjXJg
MbLIGkDoKKzKcIJwHQS6n7Qx4D1raBEYTkZixvALUNa8W/+p0OfHXy/aukSpcXi6jvKk9z5iKV0c
FmaMvBmnP1GyS6pzr1WDjbBlJQpiOt1M33+H3X2f35CpTMM+L6wlMtPdCrGrEd9MwLzLSa6BH8oA
cHbOK5Vt4kzMADvlhm8qRQwWEPzYYt0Ujw4DBwH2ykHBRFSKbqVJ8ExanW1/xz8n7EI+dTFDY5JP
zEl0Xq8T/5kQW791K9OCPLL2khfKaeMRFbWe1EfJWQ2pCHoag48sqv68ilgkz9b6eJOKUfEhk4z6
/Ao8HXQtgXMZx9P21HeZ+LpoCz0ZCf2ZLchQr/biItov0cthwen1CdllwLFzxP984z0LK0yU1S+p
SC4J9HhOHk2mLrl/b8uHg6paRk0hgsRtr8iIFtecZ10X4GKJcpnoTcv3HYLdvNm4pqne+2nw4Wug
XmuV04wC51WE2fP4VbPqni+O033YxALYo9QMhLPZYJW3PZqbcM4mLIWEzT3tB72I3RQQGoOM2yoA
BqlvcfpxKPORUT0yb82eBC1mcCFZy//SeY5ZdPD86CiNgQJJCrjhfJ8ZAXU9qxrVCP178zBpkdsK
xLs67lFOB4B8IFh0n87nfVTdN12V5+CFCNdnPwh9K2rdi6jERgbeXPnuAri9RTnC1ue4ANFYEg5k
cW36vBvcc92kqqt3vJxB9LTIcimJpXFKFGvtAOdTiG7f5BjXsho3VmBAs8aOdyPOT+MFMNMmb+CX
LsR01yIiJVy6J2B9kcmN0cWQpaH7Jg/v7EPFJ926aEftsFbHLG8eOMZftusVeKtg51oOA7HIHYZN
Fh1h2baWz4W6IqdCv6PcVf25p8HSOcbTKqjtdN8AIgO5ofhGcelny1I9gL8rpW0RcMUVOvYWJDTL
6Fmi2TFtuldKX3/n6ryl8ee6QXAULWfJHFMUlOJeU8DpJ3UN1AeW+sB7a1P64L+FtcM21euakS2o
qjcWKGy2TZIKjb6ohETYvyNVlqpBgcbyD8F2FMsxsbQyZVx1b5fGb51CfvG7WrP0WIz9CF3AxNRl
Tu8DxBd8W07EtxOZCKtQzwnWuMInhahNDQe8m8K5dmeah5Xx7kHcZdCftYXMcOsfAI1Uumq3uX9g
VWIvOWUN53fkBqrWDIml1Pw7Duqzc1Sd8CfpUpz8zVmZHCQ//ZBUkvTdbOZELGO0pAyXRMrJ0gja
l+cYELgZCmdhXaSsJVyxPp3oluOp/hj7qNVyjRvDVQfB2+2Mtlsd2PtsxapkheRrGkgGIdLM7r3c
o42t7Z+Da40PH5Xn2Ewbg7U9N6EL5d+TnAgXUEH+H4EJfjJ5BedwxTcrEUSptRdV7R7sE3nuZn5T
u4XzgUoK/DiURBb82RT4MLAgsgEUZZ9Ylt87HStZ2/BDEO3EoOBbsAh4EsWZ0IxEyLAg3fSEMa8x
RuENdb6I6ukqivutQMpXRDL2Dxco92HwE1ZjG4xa+L8D9Vg0Swf/uPCf+DzHtIL3tmkt4fzarHsz
E7JW5ogGQGTxO/p+Rv99tAJidfn97xRFaYqJzO4yHZIj2ENchJ/AtvGWXP1cSjIcunF8PhOdcEIx
4cDlMaZIZulYcDlPIxc89pylgpdFcL4Curcd+yRpxYDyhD9rJwE94yWhY7oiaRs0ssf3MB4tp7QR
ApFZA8/2wPAWGNkkESkBEd6O0wz9PmIiAZhMmALxYtPmPW1P1OjqIR8ofet5YtlA54/vcFBN5Xyk
XIPHtcY17IwK9aIhTG9cV1/Mk62F+KTAbe3mkmhEfFp6+vEwkNTk0oBoVpkKGXQ5rX4p/r7vjNYn
tXwDRWXWBMgVx4bVZhIq9P9qFOioy7k2rOYs41HfFUpeeKOMRuriy+xzA3bGBHNBWJz6JNiDSHpm
zHsYd8GOqfNo3hNcNgdOLJeuY2NWbQX6owCOt1IoBuFjQkJeFYNM04TE3BuwRtiZcaqArJqsjPmi
NeV2kq44COhXutU5P16F95yw3AQhZBG53wByKK0BcZ4qb/Q5neARWBB+jxuG4cukHqa5FnXXEYCt
zH0K80nmKrVk+0gpBnIlDuVw3Tv634tVWYhTJox5kHhV3tp9pR5xJ5zugsG5b7uwNkx6FYQh1NjQ
4QeRRr6ylKs8Kv7gr7RWHSvbE3aOds3OCW2fvAQtXIRVYMHejmLcybOxQi+c01J2OtXokKLFYKvd
ksfGv3zBneK3O+yl3sENyTl056dNTHB5KRLyUNG6ObDhTgg9G0IMWrqL10HUj/IPHchFKwJXJwAV
viF/95Y2Mh9Fmlkt3jNT4r7oLqZMStE0Hm2n5/xX4jtO8U05uk4m8v2DSQ5xRXZNFHH1vMlZw74/
rLfhSW+RJJW4USsQu+ftxt6ZWkq977N0/haiFhSQx6IaEkS6Dg/FZd/ShoRg1JsXB/TzQrbDRsVG
Fs+anwlaNVg7QOBmhp3wBckcgjpxBOv0qbJ04NS2SCpyoqjDlW95O7QCr5jjxhdIShq/jFHnzv7S
ahHSI/goIj400lWv4YKXHdyrgm34kYiozr2Mxy4c90zJu1exUwf3fwdU8LU2EYj9hKyEqpv3PAUN
Mo3fz+wJBTGfwH1Il0OxmKclTeXn7ZCkqTX9EGJAg+OVFFpCAedJIZVNa82R2aHi2h6O5CiHl2rH
aWeNKfJ9vz/EX4rNtA5HwwzQN2f9bNqiKR5BMzDHmaNvb0ms6Fcwo3kSFxqFH5SmLFt/DjmajC4I
6iaDoFdsPheK1aBW0cWvwuy3lF1yYlBYDjP4t46aLze5FhQCDh4USUaXnm/xdlNb/JM4shZttzcm
Gu+ZU3Kv/uZSRCD0BuSgSHBGGGGcfUc8HRIyzO23axMp75GVlUOygMTY2l/Q2YuWluaI0Itxsg78
CMSR4gcDWzNWWKzP/VjG63iW1ONRh+8i8kiydE94t6YoQ4wB0J7nN7FWzO3y0aLWEc+US/NK8s5d
CSlmdiSXADOlFPSBXdPM/UoKqXO1lCrUa7o09cQh9jjOVP4gB0ortbT3AuNGk1JzLoS/BNgRS7e/
cC75cFp1PJwwxwkTaLxC8iJxBNhP3knO/EaY6weMsKA6FBh5pjNF1bdcwdxes7FomaxB9abYUAqf
iZrJen5xRmgWjENU2ybsJjj/AsBm2L/Zr/Lkj/UtawP+u84c6zRRU70t/t6uGJ2UWsT9eXVFRGhM
mC2qDB+V2o918eH2NmsqkIB/k/jHktfuJPFNMoNbgp79IhHkgz0VOhU2SUPF8gxfOz6MmNSWc+gt
UE/d1V+qWpGujM8/ANp27HCSHgMJtyjD+Os/6TqlKK4Aff5n7ydeMBEMzDjaR5mROF3AFECiYFh3
IlJCzYu9+WDDfsENihlagmUkDeP5LmW0WnrRUgiRdDURp+J910QacDdrcaV6PJUF3ciI9G6Mqmny
C8ImWWUP7a68qsaIwkx16D5GUXdEPMLFATHo8YSiFocXZs2TIgg7IP3FB0vQhFSQh/i/p7Wmv3O6
/8Vem0Wj3oFI/Iz48sm+MFxxxgJuT0amXpWTSKEmwRTJG/sokhYmdo7/R3A8eGFDcssxh7/MnRdv
006yssG/vM7SZKwSfZk8U9Z8tCDB4/mgByuLs2xskIVE9QqeNZqfp9UXpt6adBkUyZMtDNgXylZA
zGUfVsHeFOclInyQl3rKbtpXPWdZr216C3LW9oxHPoeTbtnCetXxC2HRt83h+yfaDO01LX4fWUX/
XA3/809OoNGE/vqNYmIFMqmNRRk4la5xhx8qfQMVZfT68wpxmFX3sRL2o4koW4csg6BEVZhWPLOQ
U0YhoZVS7RMNBupUvEXXyuTqB/QrcnS8cezhHToIAbC1XkORvLhQ3PQSCXhUU0uwejD2REllj7TT
lCYpn0oxZ0letQTtXffP2Gn4wDRQGBcuvVNg++hX9lRDsm4oHg4eyBWka0s3fUXqagGEr4ttwm5t
3kz/FH1t8RD7K42fwUwBQXt+fFDTuk71FoYUU1E756Sj3/2DTjvre70utoYRN86NZirjDAvmTXdJ
eXpfDTW81lI+Q6gwO5OQaiekHf5fNqAv225x1TxzNPJXrlKT1sn48QqoqNsl0CiPOspEDy+v7mwJ
+PipWw9Ffb7MTcZuZD8EnlBRCCZXXAn9U8j38y8hUOBPkLxB2Rr3p9zw1AwQOYaoxAzKdFvOFwj3
AcAWqYMqyOvh2HUtIJk6tEzUZ55+yWlzjFQgR3RXIT6QJryEM+NlpVRKhtkKrmVyt5LYSmox1mSv
v1sgpy8kFoTUeZNZTutQDYhYpK41OecCHJvifvOYGBgJvOuh7u4q76wCO6VKbxsGuSN6I3kbI4vD
VaZPcItDWUJ8FfYpKVrkR4TJQaz13Aq+aoQoj2S4PqX1sTht0IuoKXT1ZVeVSEYoxAWqcG/efmCN
atYiDNsqAQdvb9/AkqQ9G2AiUPz/9gKvMP8Fm12bw11RVptTdVyI/JAvZITe40GNWA+nmKW+qL/P
cqkqRZ0HV1b4F8AAsKG6KBt3wh/kjr83+ru0TdXYRDGnyZ/xLkb67s8kHohs7pY3YrJZEYNVezoG
QQV82T8jyN2dTJ7Xu0JnVOIfTcvMvlmbmxKOqVtWxsuAhHRFuYBJLFBUahWYDBVMXmJ4+YWp7JTU
aRk0Geb5zx8i4sq8PZxFGKSh87aTpq1bDqg5rwxOiz6TlI4WRfi+INUnWhc7yT4UYpjh1htsoSpt
7KJAlfBZxVvh33gNrKSJG+A46UI50WdOyqwYoRtjEhCDzgv7cCjaCwg+qtERZ1GedF0GChG5IFCx
8pg/Gb/GpzXP+ITqT9KfxI3z2v9edpcfiTsgSjkEkvbaowwdzxTbZt+aDBCjq3dKxaCz0N0ehFct
lRdQHpVEaJpgJrd7QRSOX3JrBS97/QBad65nIUnM87jcAyXgqBPlG2cqv487ZdpzzPteBTFD5XuZ
u1Q2480bZQp0IgptA0LcgJ+GGchUbw6i1tSR0WGjmajbrHOzS4PY08hbi9n9l4eVEJh0aMBsjzKA
8P3LsneroUxaEuBArk0PY6OyLqCLSX3/22ZNoEY0ugG0rqQiz+eMdUFTnb6+4ktNG+q6o4kKOQRU
IvomnsRvP5lUzR3hGZ9kg8f5kV5XgujpVCZ4sEk7BdMnS6dgs676eToJQojfng1ygs8sJggZL+os
KyjpvPD35YOVl4btnnN1SZS0EugbL+8FdP9YCSafxkGXvxODqRc9vQrdvre60Jpwod96Yk/pDXf6
CYzS5jgbwqk2XGvMsxRhYLgHaXSHtVR2WhRJmnY6qmSKkdfZIqYOHtmPGmTL+UN/A1azSk+BQcO2
4qBWDJefVJF0/SiOJej7C7TVx9vZylzKwIgvaoBabOiIUiy2sZ7D+yPJ0ouMXetO3g4Hr2/Jtcw/
xqiCz/ISFx55J5hW+23VIE3cfjuwAoUDrIjfC5sFmS0ItAOZ+Qxkf7fCmg2ruMEegLcAtPDeiUkD
CNXApdZl6beXDFPe6vYXaW5ftu475RRneAstwKsZHZKvZOoRLEpHwWix821d4wASS8TyLILKKkcJ
yPHdw3KZqo5NFFR0LzAUlnvFNM+cODi5iJSe69DJnQp9A2BOzIxZZ7/+xY/3NDmcgKrdR8xwVpl8
bFlLwK1Gxd9Ea9K03uZa+CHCdtPBfv3KH+2zopSUqeAYzsQ99J6CqE7OjzmPRxmoLhn+tCWmKWpv
TEc5Swo/AxENtZQ0R3J9EnNEzA/RxswV1v+N3yjhbDMG6lS1KhYN1o20n4Q4KPsyPXMZxIUiaPfS
MllFCsXk2dIVG7I4rox3dKtu8AzlVWboUUFLHs9OFEfGUBHipOB0gBPOJUVXBfdAewt8MIGLSop2
KOsk9+4DSaItOtO9Rf0FK7S2wSOygluQ/MDRApSF3fjYfKmVelx9Df5xluw5BlUnjIIzq4C+jTBM
IMv3x+byZCphoLmkgidy8qR7nGO5vBlqP8a3b1l90gn45vxHOAo7+vGRjs+K8YGYQ7NUlytzuwxl
+7+TIfhkbWb4+pi5APm9p05+j4hJPYymXsDYEKhFvRgXRY9GqWtisY1M4kPAhkLA7ok3py59DcnC
dxs1vaGZFlllVWqWXRo66TCQg9jSFHZf3jJ20HF6FIeJYswWGahx2uRxbFTuf94D0aHYFYizDKQp
9fgKFx0i2Rcwb3CwEXw++axZ1WmI+dAidd5hOkNFZGbWTfXvcUYPdzngDOCGhCjS18QX8j8l6uHw
cWP15G35NQlsXFCcA+RgmVvYBCiDF7JKebSu6DGkAdT4b315EfMNSGH7l/HvHDZ+nC8frZ6K6O2e
HTNxNPDM8G20OGL1V4nFEJq92p9bDYgkzRWnkqIPYYX1ppBI1K2t8XNd88zMhPdQAjMT19bejAty
ujOjUz4JtaffD54kDQPy5OIIWktppwwFHMN2+iWjIMdgvGk3FJY6VAGpC+ISESoL3ePmCZaoH5tj
1XilsM/Hln1KkmVs/DKbMCLIso9WBYeyGOjtta0YrZo3J53JRBm3ILQxFHVy3IzVxtvIXVxPBqJN
pygFt11xQ2Fyn1KbG+1FsIGdVvrhAAFgfMq9y31a1ssjtYjk5Cqdm3W32vU01JRrPVdTq1aTOYFJ
uhfrthmOln9f+cPM+/7fhtBC3+GTSYnwCmCh/vxyPaKrIFdRIfO+AeTjcaizfwGu59BBrexJ9GvH
f2UK170QhM4TBuJa6QBLmUDtPAKw4R6ZRdpHeFYXK8/ECgEyYVjDLGuxatT5n/6ewK8eCTrFHqmN
1l6RSLR+JuakjZ4sH/D51etKcEjByjuJFG/pSXVSBhIeJcCIQtUTVAZqk/BmgXsbKDyIBwUeO/yl
E6pHWYXPnKlTcqH3tycJxxLJHMQACp/yk+UTG6cz/8HMt66RS0Xpq9CaMPH13AmMl7ml82XvXDUZ
OTjmLvNnZ90jCIF5c6wUTpOYlBanLDT+MQr7Cmt5RoF3lObuwdWYYgXZZakStlAOP3SaOUyNLfgb
ItXan3MtR8Y1aosjWgLbgA/vhYmwXgUh2JBT4Ev+1hhRoYi3mM+uTu8HbBI=
`protect end_protected

