module return_conf(
   // clk
   input clk,
   input reset,
   // Configuration via UART
   input    wire [9:0]    conf_addr_r,      // host: pc, core: esn
   input    wire          conf_c2h_en_r,
   output   reg  [15:0]   conf_c2h_d,       // core-to-host data
   // Registers
   input wire [15:0] w_in [0:7][0:39],       // input weights for 16 neurons x 4 inputs
   input wire [15:0] w_x [0:7][0:7],       // reservoir weights rn0~rn15
   input wire [15:0] w_out [0:3][0:47]       // output weights 2 output nodes x 20 (rstate + input)
);
   
   always@ (posedge clk) begin
      if (reset) begin
         conf_c2h_d <= 16'd0;
      end
      else if (conf_c2h_en_r) begin
         case (conf_addr_r)
            10'd0: begin conf_c2h_d <= w_in[0][0]; end
            10'd1: begin conf_c2h_d <= w_in[0][1]; end
            10'd2: begin conf_c2h_d <= w_in[0][2]; end
            10'd3: begin conf_c2h_d <= w_in[0][3]; end
            10'd4: begin conf_c2h_d <= w_in[0][4]; end
            10'd5: begin conf_c2h_d <= w_in[0][5]; end
            10'd6: begin conf_c2h_d <= w_in[0][6]; end
            10'd7: begin conf_c2h_d <= w_in[0][7]; end
            10'd8: begin conf_c2h_d <= w_in[0][8]; end
            10'd9: begin conf_c2h_d <= w_in[0][9]; end
            10'd10: begin conf_c2h_d <= w_in[0][10]; end
            10'd11: begin conf_c2h_d <= w_in[0][11]; end
            10'd12: begin conf_c2h_d <= w_in[0][12]; end
            10'd13: begin conf_c2h_d <= w_in[0][13]; end
            10'd14: begin conf_c2h_d <= w_in[0][14]; end
            10'd15: begin conf_c2h_d <= w_in[0][15]; end
            10'd16: begin conf_c2h_d <= w_in[0][16]; end
            10'd17: begin conf_c2h_d <= w_in[0][17]; end
            10'd18: begin conf_c2h_d <= w_in[0][18]; end
            10'd19: begin conf_c2h_d <= w_in[0][19]; end
            10'd20: begin conf_c2h_d <= w_in[0][20]; end
            10'd21: begin conf_c2h_d <= w_in[0][21]; end
            10'd22: begin conf_c2h_d <= w_in[0][22]; end
            10'd23: begin conf_c2h_d <= w_in[0][23]; end
            10'd24: begin conf_c2h_d <= w_in[0][24]; end
            10'd25: begin conf_c2h_d <= w_in[0][25]; end
            10'd26: begin conf_c2h_d <= w_in[0][26]; end
            10'd27: begin conf_c2h_d <= w_in[0][27]; end
            10'd28: begin conf_c2h_d <= w_in[0][28]; end
            10'd29: begin conf_c2h_d <= w_in[0][29]; end
            10'd30: begin conf_c2h_d <= w_in[0][30]; end
            10'd31: begin conf_c2h_d <= w_in[0][31]; end
            10'd32: begin conf_c2h_d <= w_in[0][32]; end
            10'd33: begin conf_c2h_d <= w_in[0][33]; end
            10'd34: begin conf_c2h_d <= w_in[0][34]; end
            10'd35: begin conf_c2h_d <= w_in[0][35]; end
            10'd36: begin conf_c2h_d <= w_in[0][36]; end
            10'd37: begin conf_c2h_d <= w_in[0][37]; end
            10'd38: begin conf_c2h_d <= w_in[0][38]; end
            10'd39: begin conf_c2h_d <= w_in[0][39]; end
            10'd40: begin conf_c2h_d <= w_in[1][0]; end
            10'd41: begin conf_c2h_d <= w_in[1][1]; end
            10'd42: begin conf_c2h_d <= w_in[1][2]; end
            10'd43: begin conf_c2h_d <= w_in[1][3]; end
            10'd44: begin conf_c2h_d <= w_in[1][4]; end
            10'd45: begin conf_c2h_d <= w_in[1][5]; end
            10'd46: begin conf_c2h_d <= w_in[1][6]; end
            10'd47: begin conf_c2h_d <= w_in[1][7]; end
            10'd48: begin conf_c2h_d <= w_in[1][8]; end
            10'd49: begin conf_c2h_d <= w_in[1][9]; end
            10'd50: begin conf_c2h_d <= w_in[1][10]; end
            10'd51: begin conf_c2h_d <= w_in[1][11]; end
            10'd52: begin conf_c2h_d <= w_in[1][12]; end
            10'd53: begin conf_c2h_d <= w_in[1][13]; end
            10'd54: begin conf_c2h_d <= w_in[1][14]; end
            10'd55: begin conf_c2h_d <= w_in[1][15]; end
            10'd56: begin conf_c2h_d <= w_in[1][16]; end
            10'd57: begin conf_c2h_d <= w_in[1][17]; end
            10'd58: begin conf_c2h_d <= w_in[1][18]; end
            10'd59: begin conf_c2h_d <= w_in[1][19]; end
            10'd60: begin conf_c2h_d <= w_in[1][20]; end
            10'd61: begin conf_c2h_d <= w_in[1][21]; end
            10'd62: begin conf_c2h_d <= w_in[1][22]; end
            10'd63: begin conf_c2h_d <= w_in[1][23]; end
            10'd64: begin conf_c2h_d <= w_in[1][24]; end
            10'd65: begin conf_c2h_d <= w_in[1][25]; end
            10'd66: begin conf_c2h_d <= w_in[1][26]; end
            10'd67: begin conf_c2h_d <= w_in[1][27]; end
            10'd68: begin conf_c2h_d <= w_in[1][28]; end
            10'd69: begin conf_c2h_d <= w_in[1][29]; end
            10'd70: begin conf_c2h_d <= w_in[1][30]; end
            10'd71: begin conf_c2h_d <= w_in[1][31]; end
            10'd72: begin conf_c2h_d <= w_in[1][32]; end
            10'd73: begin conf_c2h_d <= w_in[1][33]; end
            10'd74: begin conf_c2h_d <= w_in[1][34]; end
            10'd75: begin conf_c2h_d <= w_in[1][35]; end
            10'd76: begin conf_c2h_d <= w_in[1][36]; end
            10'd77: begin conf_c2h_d <= w_in[1][37]; end
            10'd78: begin conf_c2h_d <= w_in[1][38]; end
            10'd79: begin conf_c2h_d <= w_in[1][39]; end
            10'd80: begin conf_c2h_d <= w_in[2][0]; end
            10'd81: begin conf_c2h_d <= w_in[2][1]; end
            10'd82: begin conf_c2h_d <= w_in[2][2]; end
            10'd83: begin conf_c2h_d <= w_in[2][3]; end
            10'd84: begin conf_c2h_d <= w_in[2][4]; end
            10'd85: begin conf_c2h_d <= w_in[2][5]; end
            10'd86: begin conf_c2h_d <= w_in[2][6]; end
            10'd87: begin conf_c2h_d <= w_in[2][7]; end
            10'd88: begin conf_c2h_d <= w_in[2][8]; end
            10'd89: begin conf_c2h_d <= w_in[2][9]; end
            10'd90: begin conf_c2h_d <= w_in[2][10]; end
            10'd91: begin conf_c2h_d <= w_in[2][11]; end
            10'd92: begin conf_c2h_d <= w_in[2][12]; end
            10'd93: begin conf_c2h_d <= w_in[2][13]; end
            10'd94: begin conf_c2h_d <= w_in[2][14]; end
            10'd95: begin conf_c2h_d <= w_in[2][15]; end
            10'd96: begin conf_c2h_d <= w_in[2][16]; end
            10'd97: begin conf_c2h_d <= w_in[2][17]; end
            10'd98: begin conf_c2h_d <= w_in[2][18]; end
            10'd99: begin conf_c2h_d <= w_in[2][19]; end
            10'd100: begin conf_c2h_d <= w_in[2][20]; end
            10'd101: begin conf_c2h_d <= w_in[2][21]; end
            10'd102: begin conf_c2h_d <= w_in[2][22]; end
            10'd103: begin conf_c2h_d <= w_in[2][23]; end
            10'd104: begin conf_c2h_d <= w_in[2][24]; end
            10'd105: begin conf_c2h_d <= w_in[2][25]; end
            10'd106: begin conf_c2h_d <= w_in[2][26]; end
            10'd107: begin conf_c2h_d <= w_in[2][27]; end
            10'd108: begin conf_c2h_d <= w_in[2][28]; end
            10'd109: begin conf_c2h_d <= w_in[2][29]; end
            10'd110: begin conf_c2h_d <= w_in[2][30]; end
            10'd111: begin conf_c2h_d <= w_in[2][31]; end
            10'd112: begin conf_c2h_d <= w_in[2][32]; end
            10'd113: begin conf_c2h_d <= w_in[2][33]; end
            10'd114: begin conf_c2h_d <= w_in[2][34]; end
            10'd115: begin conf_c2h_d <= w_in[2][35]; end
            10'd116: begin conf_c2h_d <= w_in[2][36]; end
            10'd117: begin conf_c2h_d <= w_in[2][37]; end
            10'd118: begin conf_c2h_d <= w_in[2][38]; end
            10'd119: begin conf_c2h_d <= w_in[2][39]; end
            10'd120: begin conf_c2h_d <= w_in[3][0]; end
            10'd121: begin conf_c2h_d <= w_in[3][1]; end
            10'd122: begin conf_c2h_d <= w_in[3][2]; end
            10'd123: begin conf_c2h_d <= w_in[3][3]; end
            10'd124: begin conf_c2h_d <= w_in[3][4]; end
            10'd125: begin conf_c2h_d <= w_in[3][5]; end
            10'd126: begin conf_c2h_d <= w_in[3][6]; end
            10'd127: begin conf_c2h_d <= w_in[3][7]; end
            10'd128: begin conf_c2h_d <= w_in[3][8]; end
            10'd129: begin conf_c2h_d <= w_in[3][9]; end
            10'd130: begin conf_c2h_d <= w_in[3][10]; end
            10'd131: begin conf_c2h_d <= w_in[3][11]; end
            10'd132: begin conf_c2h_d <= w_in[3][12]; end
            10'd133: begin conf_c2h_d <= w_in[3][13]; end
            10'd134: begin conf_c2h_d <= w_in[3][14]; end
            10'd135: begin conf_c2h_d <= w_in[3][15]; end
            10'd136: begin conf_c2h_d <= w_in[3][16]; end
            10'd137: begin conf_c2h_d <= w_in[3][17]; end
            10'd138: begin conf_c2h_d <= w_in[3][18]; end
            10'd139: begin conf_c2h_d <= w_in[3][19]; end
            10'd140: begin conf_c2h_d <= w_in[3][20]; end
            10'd141: begin conf_c2h_d <= w_in[3][21]; end
            10'd142: begin conf_c2h_d <= w_in[3][22]; end
            10'd143: begin conf_c2h_d <= w_in[3][23]; end
            10'd144: begin conf_c2h_d <= w_in[3][24]; end
            10'd145: begin conf_c2h_d <= w_in[3][25]; end
            10'd146: begin conf_c2h_d <= w_in[3][26]; end
            10'd147: begin conf_c2h_d <= w_in[3][27]; end
            10'd148: begin conf_c2h_d <= w_in[3][28]; end
            10'd149: begin conf_c2h_d <= w_in[3][29]; end
            10'd150: begin conf_c2h_d <= w_in[3][30]; end
            10'd151: begin conf_c2h_d <= w_in[3][31]; end
            10'd152: begin conf_c2h_d <= w_in[3][32]; end
            10'd153: begin conf_c2h_d <= w_in[3][33]; end
            10'd154: begin conf_c2h_d <= w_in[3][34]; end
            10'd155: begin conf_c2h_d <= w_in[3][35]; end
            10'd156: begin conf_c2h_d <= w_in[3][36]; end
            10'd157: begin conf_c2h_d <= w_in[3][37]; end
            10'd158: begin conf_c2h_d <= w_in[3][38]; end
            10'd159: begin conf_c2h_d <= w_in[3][39]; end
            10'd160: begin conf_c2h_d <= w_in[4][0]; end
            10'd161: begin conf_c2h_d <= w_in[4][1]; end
            10'd162: begin conf_c2h_d <= w_in[4][2]; end
            10'd163: begin conf_c2h_d <= w_in[4][3]; end
            10'd164: begin conf_c2h_d <= w_in[4][4]; end
            10'd165: begin conf_c2h_d <= w_in[4][5]; end
            10'd166: begin conf_c2h_d <= w_in[4][6]; end
            10'd167: begin conf_c2h_d <= w_in[4][7]; end
            10'd168: begin conf_c2h_d <= w_in[4][8]; end
            10'd169: begin conf_c2h_d <= w_in[4][9]; end
            10'd170: begin conf_c2h_d <= w_in[4][10]; end
            10'd171: begin conf_c2h_d <= w_in[4][11]; end
            10'd172: begin conf_c2h_d <= w_in[4][12]; end
            10'd173: begin conf_c2h_d <= w_in[4][13]; end
            10'd174: begin conf_c2h_d <= w_in[4][14]; end
            10'd175: begin conf_c2h_d <= w_in[4][15]; end
            10'd176: begin conf_c2h_d <= w_in[4][16]; end
            10'd177: begin conf_c2h_d <= w_in[4][17]; end
            10'd178: begin conf_c2h_d <= w_in[4][18]; end
            10'd179: begin conf_c2h_d <= w_in[4][19]; end
            10'd180: begin conf_c2h_d <= w_in[4][20]; end
            10'd181: begin conf_c2h_d <= w_in[4][21]; end
            10'd182: begin conf_c2h_d <= w_in[4][22]; end
            10'd183: begin conf_c2h_d <= w_in[4][23]; end
            10'd184: begin conf_c2h_d <= w_in[4][24]; end
            10'd185: begin conf_c2h_d <= w_in[4][25]; end
            10'd186: begin conf_c2h_d <= w_in[4][26]; end
            10'd187: begin conf_c2h_d <= w_in[4][27]; end
            10'd188: begin conf_c2h_d <= w_in[4][28]; end
            10'd189: begin conf_c2h_d <= w_in[4][29]; end
            10'd190: begin conf_c2h_d <= w_in[4][30]; end
            10'd191: begin conf_c2h_d <= w_in[4][31]; end
            10'd192: begin conf_c2h_d <= w_in[4][32]; end
            10'd193: begin conf_c2h_d <= w_in[4][33]; end
            10'd194: begin conf_c2h_d <= w_in[4][34]; end
            10'd195: begin conf_c2h_d <= w_in[4][35]; end
            10'd196: begin conf_c2h_d <= w_in[4][36]; end
            10'd197: begin conf_c2h_d <= w_in[4][37]; end
            10'd198: begin conf_c2h_d <= w_in[4][38]; end
            10'd199: begin conf_c2h_d <= w_in[4][39]; end
            10'd200: begin conf_c2h_d <= w_in[5][0]; end
            10'd201: begin conf_c2h_d <= w_in[5][1]; end
            10'd202: begin conf_c2h_d <= w_in[5][2]; end
            10'd203: begin conf_c2h_d <= w_in[5][3]; end
            10'd204: begin conf_c2h_d <= w_in[5][4]; end
            10'd205: begin conf_c2h_d <= w_in[5][5]; end
            10'd206: begin conf_c2h_d <= w_in[5][6]; end
            10'd207: begin conf_c2h_d <= w_in[5][7]; end
            10'd208: begin conf_c2h_d <= w_in[5][8]; end
            10'd209: begin conf_c2h_d <= w_in[5][9]; end
            10'd210: begin conf_c2h_d <= w_in[5][10]; end
            10'd211: begin conf_c2h_d <= w_in[5][11]; end
            10'd212: begin conf_c2h_d <= w_in[5][12]; end
            10'd213: begin conf_c2h_d <= w_in[5][13]; end
            10'd214: begin conf_c2h_d <= w_in[5][14]; end
            10'd215: begin conf_c2h_d <= w_in[5][15]; end
            10'd216: begin conf_c2h_d <= w_in[5][16]; end
            10'd217: begin conf_c2h_d <= w_in[5][17]; end
            10'd218: begin conf_c2h_d <= w_in[5][18]; end
            10'd219: begin conf_c2h_d <= w_in[5][19]; end
            10'd220: begin conf_c2h_d <= w_in[5][20]; end
            10'd221: begin conf_c2h_d <= w_in[5][21]; end
            10'd222: begin conf_c2h_d <= w_in[5][22]; end
            10'd223: begin conf_c2h_d <= w_in[5][23]; end
            10'd224: begin conf_c2h_d <= w_in[5][24]; end
            10'd225: begin conf_c2h_d <= w_in[5][25]; end
            10'd226: begin conf_c2h_d <= w_in[5][26]; end
            10'd227: begin conf_c2h_d <= w_in[5][27]; end
            10'd228: begin conf_c2h_d <= w_in[5][28]; end
            10'd229: begin conf_c2h_d <= w_in[5][29]; end
            10'd230: begin conf_c2h_d <= w_in[5][30]; end
            10'd231: begin conf_c2h_d <= w_in[5][31]; end
            10'd232: begin conf_c2h_d <= w_in[5][32]; end
            10'd233: begin conf_c2h_d <= w_in[5][33]; end
            10'd234: begin conf_c2h_d <= w_in[5][34]; end
            10'd235: begin conf_c2h_d <= w_in[5][35]; end
            10'd236: begin conf_c2h_d <= w_in[5][36]; end
            10'd237: begin conf_c2h_d <= w_in[5][37]; end
            10'd238: begin conf_c2h_d <= w_in[5][38]; end
            10'd239: begin conf_c2h_d <= w_in[5][39]; end
            10'd240: begin conf_c2h_d <= w_in[6][0]; end
            10'd241: begin conf_c2h_d <= w_in[6][1]; end
            10'd242: begin conf_c2h_d <= w_in[6][2]; end
            10'd243: begin conf_c2h_d <= w_in[6][3]; end
            10'd244: begin conf_c2h_d <= w_in[6][4]; end
            10'd245: begin conf_c2h_d <= w_in[6][5]; end
            10'd246: begin conf_c2h_d <= w_in[6][6]; end
            10'd247: begin conf_c2h_d <= w_in[6][7]; end
            10'd248: begin conf_c2h_d <= w_in[6][8]; end
            10'd249: begin conf_c2h_d <= w_in[6][9]; end
            10'd250: begin conf_c2h_d <= w_in[6][10]; end
            10'd251: begin conf_c2h_d <= w_in[6][11]; end
            10'd252: begin conf_c2h_d <= w_in[6][12]; end
            10'd253: begin conf_c2h_d <= w_in[6][13]; end
            10'd254: begin conf_c2h_d <= w_in[6][14]; end
            10'd255: begin conf_c2h_d <= w_in[6][15]; end
            10'd256: begin conf_c2h_d <= w_in[6][16]; end
            10'd257: begin conf_c2h_d <= w_in[6][17]; end
            10'd258: begin conf_c2h_d <= w_in[6][18]; end
            10'd259: begin conf_c2h_d <= w_in[6][19]; end
            10'd260: begin conf_c2h_d <= w_in[6][20]; end
            10'd261: begin conf_c2h_d <= w_in[6][21]; end
            10'd262: begin conf_c2h_d <= w_in[6][22]; end
            10'd263: begin conf_c2h_d <= w_in[6][23]; end
            10'd264: begin conf_c2h_d <= w_in[6][24]; end
            10'd265: begin conf_c2h_d <= w_in[6][25]; end
            10'd266: begin conf_c2h_d <= w_in[6][26]; end
            10'd267: begin conf_c2h_d <= w_in[6][27]; end
            10'd268: begin conf_c2h_d <= w_in[6][28]; end
            10'd269: begin conf_c2h_d <= w_in[6][29]; end
            10'd270: begin conf_c2h_d <= w_in[6][30]; end
            10'd271: begin conf_c2h_d <= w_in[6][31]; end
            10'd272: begin conf_c2h_d <= w_in[6][32]; end
            10'd273: begin conf_c2h_d <= w_in[6][33]; end
            10'd274: begin conf_c2h_d <= w_in[6][34]; end
            10'd275: begin conf_c2h_d <= w_in[6][35]; end
            10'd276: begin conf_c2h_d <= w_in[6][36]; end
            10'd277: begin conf_c2h_d <= w_in[6][37]; end
            10'd278: begin conf_c2h_d <= w_in[6][38]; end
            10'd279: begin conf_c2h_d <= w_in[6][39]; end
            10'd280: begin conf_c2h_d <= w_in[7][0]; end
            10'd281: begin conf_c2h_d <= w_in[7][1]; end
            10'd282: begin conf_c2h_d <= w_in[7][2]; end
            10'd283: begin conf_c2h_d <= w_in[7][3]; end
            10'd284: begin conf_c2h_d <= w_in[7][4]; end
            10'd285: begin conf_c2h_d <= w_in[7][5]; end
            10'd286: begin conf_c2h_d <= w_in[7][6]; end
            10'd287: begin conf_c2h_d <= w_in[7][7]; end
            10'd288: begin conf_c2h_d <= w_in[7][8]; end
            10'd289: begin conf_c2h_d <= w_in[7][9]; end
            10'd290: begin conf_c2h_d <= w_in[7][10]; end
            10'd291: begin conf_c2h_d <= w_in[7][11]; end
            10'd292: begin conf_c2h_d <= w_in[7][12]; end
            10'd293: begin conf_c2h_d <= w_in[7][13]; end
            10'd294: begin conf_c2h_d <= w_in[7][14]; end
            10'd295: begin conf_c2h_d <= w_in[7][15]; end
            10'd296: begin conf_c2h_d <= w_in[7][16]; end
            10'd297: begin conf_c2h_d <= w_in[7][17]; end
            10'd298: begin conf_c2h_d <= w_in[7][18]; end
            10'd299: begin conf_c2h_d <= w_in[7][19]; end
            10'd300: begin conf_c2h_d <= w_in[7][20]; end
            10'd301: begin conf_c2h_d <= w_in[7][21]; end
            10'd302: begin conf_c2h_d <= w_in[7][22]; end
            10'd303: begin conf_c2h_d <= w_in[7][23]; end
            10'd304: begin conf_c2h_d <= w_in[7][24]; end
            10'd305: begin conf_c2h_d <= w_in[7][25]; end
            10'd306: begin conf_c2h_d <= w_in[7][26]; end
            10'd307: begin conf_c2h_d <= w_in[7][27]; end
            10'd308: begin conf_c2h_d <= w_in[7][28]; end
            10'd309: begin conf_c2h_d <= w_in[7][29]; end
            10'd310: begin conf_c2h_d <= w_in[7][30]; end
            10'd311: begin conf_c2h_d <= w_in[7][31]; end
            10'd312: begin conf_c2h_d <= w_in[7][32]; end
            10'd313: begin conf_c2h_d <= w_in[7][33]; end
            10'd314: begin conf_c2h_d <= w_in[7][34]; end
            10'd315: begin conf_c2h_d <= w_in[7][35]; end
            10'd316: begin conf_c2h_d <= w_in[7][36]; end
            10'd317: begin conf_c2h_d <= w_in[7][37]; end
            10'd318: begin conf_c2h_d <= w_in[7][38]; end
            10'd319: begin conf_c2h_d <= w_in[7][39]; end

            //----- w_out -----
            10'd320: begin conf_c2h_d <= w_out[0][0]; end
            10'd321: begin conf_c2h_d <= w_out[0][1]; end
            10'd322: begin conf_c2h_d <= w_out[0][2]; end
            10'd323: begin conf_c2h_d <= w_out[0][3]; end
            10'd324: begin conf_c2h_d <= w_out[0][4]; end
            10'd325: begin conf_c2h_d <= w_out[0][5]; end
            10'd326: begin conf_c2h_d <= w_out[0][6]; end
            10'd327: begin conf_c2h_d <= w_out[0][7]; end
            10'd328: begin conf_c2h_d <= w_out[0][8]; end
            10'd329: begin conf_c2h_d <= w_out[0][9]; end
            10'd330: begin conf_c2h_d <= w_out[0][10]; end
            10'd331: begin conf_c2h_d <= w_out[0][11]; end
            10'd332: begin conf_c2h_d <= w_out[0][12]; end
            10'd333: begin conf_c2h_d <= w_out[0][13]; end
            10'd334: begin conf_c2h_d <= w_out[0][14]; end
            10'd335: begin conf_c2h_d <= w_out[0][15]; end
            10'd336: begin conf_c2h_d <= w_out[0][16]; end
            10'd337: begin conf_c2h_d <= w_out[0][17]; end
            10'd338: begin conf_c2h_d <= w_out[0][18]; end
            10'd339: begin conf_c2h_d <= w_out[0][19]; end
            10'd340: begin conf_c2h_d <= w_out[0][20]; end
            10'd341: begin conf_c2h_d <= w_out[0][21]; end
            10'd342: begin conf_c2h_d <= w_out[0][22]; end
            10'd343: begin conf_c2h_d <= w_out[0][23]; end
            10'd344: begin conf_c2h_d <= w_out[0][24]; end
            10'd345: begin conf_c2h_d <= w_out[0][25]; end
            10'd346: begin conf_c2h_d <= w_out[0][26]; end
            10'd347: begin conf_c2h_d <= w_out[0][27]; end
            10'd348: begin conf_c2h_d <= w_out[0][28]; end
            10'd349: begin conf_c2h_d <= w_out[0][29]; end
            10'd350: begin conf_c2h_d <= w_out[0][30]; end
            10'd351: begin conf_c2h_d <= w_out[0][31]; end
            10'd352: begin conf_c2h_d <= w_out[0][32]; end
            10'd353: begin conf_c2h_d <= w_out[0][33]; end
            10'd354: begin conf_c2h_d <= w_out[0][34]; end
            10'd355: begin conf_c2h_d <= w_out[0][35]; end
            10'd356: begin conf_c2h_d <= w_out[0][36]; end
            10'd357: begin conf_c2h_d <= w_out[0][37]; end
            10'd358: begin conf_c2h_d <= w_out[0][38]; end
            10'd359: begin conf_c2h_d <= w_out[0][39]; end
            10'd360: begin conf_c2h_d <= w_out[0][40]; end
            10'd361: begin conf_c2h_d <= w_out[0][41]; end
            10'd362: begin conf_c2h_d <= w_out[0][42]; end
            10'd363: begin conf_c2h_d <= w_out[0][43]; end
            10'd364: begin conf_c2h_d <= w_out[0][44]; end
            10'd365: begin conf_c2h_d <= w_out[0][45]; end
            10'd366: begin conf_c2h_d <= w_out[0][46]; end
            10'd367: begin conf_c2h_d <= w_out[0][47]; end
            10'd368: begin conf_c2h_d <= w_out[1][0]; end
            10'd369: begin conf_c2h_d <= w_out[1][1]; end
            10'd370: begin conf_c2h_d <= w_out[1][2]; end
            10'd371: begin conf_c2h_d <= w_out[1][3]; end
            10'd372: begin conf_c2h_d <= w_out[1][4]; end
            10'd373: begin conf_c2h_d <= w_out[1][5]; end
            10'd374: begin conf_c2h_d <= w_out[1][6]; end
            10'd375: begin conf_c2h_d <= w_out[1][7]; end
            10'd376: begin conf_c2h_d <= w_out[1][8]; end
            10'd377: begin conf_c2h_d <= w_out[1][9]; end
            10'd378: begin conf_c2h_d <= w_out[1][10]; end
            10'd379: begin conf_c2h_d <= w_out[1][11]; end
            10'd380: begin conf_c2h_d <= w_out[1][12]; end
            10'd381: begin conf_c2h_d <= w_out[1][13]; end
            10'd382: begin conf_c2h_d <= w_out[1][14]; end
            10'd383: begin conf_c2h_d <= w_out[1][15]; end
            10'd384: begin conf_c2h_d <= w_out[1][16]; end
            10'd385: begin conf_c2h_d <= w_out[1][17]; end
            10'd386: begin conf_c2h_d <= w_out[1][18]; end
            10'd387: begin conf_c2h_d <= w_out[1][19]; end
            10'd388: begin conf_c2h_d <= w_out[1][20]; end
            10'd389: begin conf_c2h_d <= w_out[1][21]; end
            10'd390: begin conf_c2h_d <= w_out[1][22]; end
            10'd391: begin conf_c2h_d <= w_out[1][23]; end
            10'd392: begin conf_c2h_d <= w_out[1][24]; end
            10'd393: begin conf_c2h_d <= w_out[1][25]; end
            10'd394: begin conf_c2h_d <= w_out[1][26]; end
            10'd395: begin conf_c2h_d <= w_out[1][27]; end
            10'd396: begin conf_c2h_d <= w_out[1][28]; end
            10'd397: begin conf_c2h_d <= w_out[1][29]; end
            10'd398: begin conf_c2h_d <= w_out[1][30]; end
            10'd399: begin conf_c2h_d <= w_out[1][31]; end
            10'd400: begin conf_c2h_d <= w_out[1][32]; end
            10'd401: begin conf_c2h_d <= w_out[1][33]; end
            10'd402: begin conf_c2h_d <= w_out[1][34]; end
            10'd403: begin conf_c2h_d <= w_out[1][35]; end
            10'd404: begin conf_c2h_d <= w_out[1][36]; end
            10'd405: begin conf_c2h_d <= w_out[1][37]; end
            10'd406: begin conf_c2h_d <= w_out[1][38]; end
            10'd407: begin conf_c2h_d <= w_out[1][39]; end
            10'd408: begin conf_c2h_d <= w_out[1][40]; end
            10'd409: begin conf_c2h_d <= w_out[1][41]; end
            10'd410: begin conf_c2h_d <= w_out[1][42]; end
            10'd411: begin conf_c2h_d <= w_out[1][43]; end
            10'd412: begin conf_c2h_d <= w_out[1][44]; end
            10'd413: begin conf_c2h_d <= w_out[1][45]; end
            10'd414: begin conf_c2h_d <= w_out[1][46]; end
            10'd415: begin conf_c2h_d <= w_out[1][47]; end
            10'd416: begin conf_c2h_d <= w_out[2][0]; end
            10'd417: begin conf_c2h_d <= w_out[2][1]; end
            10'd418: begin conf_c2h_d <= w_out[2][2]; end
            10'd419: begin conf_c2h_d <= w_out[2][3]; end
            10'd420: begin conf_c2h_d <= w_out[2][4]; end
            10'd421: begin conf_c2h_d <= w_out[2][5]; end
            10'd422: begin conf_c2h_d <= w_out[2][6]; end
            10'd423: begin conf_c2h_d <= w_out[2][7]; end
            10'd424: begin conf_c2h_d <= w_out[2][8]; end
            10'd425: begin conf_c2h_d <= w_out[2][9]; end
            10'd426: begin conf_c2h_d <= w_out[2][10]; end
            10'd427: begin conf_c2h_d <= w_out[2][11]; end
            10'd428: begin conf_c2h_d <= w_out[2][12]; end
            10'd429: begin conf_c2h_d <= w_out[2][13]; end
            10'd430: begin conf_c2h_d <= w_out[2][14]; end
            10'd431: begin conf_c2h_d <= w_out[2][15]; end
            10'd432: begin conf_c2h_d <= w_out[2][16]; end
            10'd433: begin conf_c2h_d <= w_out[2][17]; end
            10'd434: begin conf_c2h_d <= w_out[2][18]; end
            10'd435: begin conf_c2h_d <= w_out[2][19]; end
            10'd436: begin conf_c2h_d <= w_out[2][20]; end
            10'd437: begin conf_c2h_d <= w_out[2][21]; end
            10'd438: begin conf_c2h_d <= w_out[2][22]; end
            10'd439: begin conf_c2h_d <= w_out[2][23]; end
            10'd440: begin conf_c2h_d <= w_out[2][24]; end
            10'd441: begin conf_c2h_d <= w_out[2][25]; end
            10'd442: begin conf_c2h_d <= w_out[2][26]; end
            10'd443: begin conf_c2h_d <= w_out[2][27]; end
            10'd444: begin conf_c2h_d <= w_out[2][28]; end
            10'd445: begin conf_c2h_d <= w_out[2][29]; end
            10'd446: begin conf_c2h_d <= w_out[2][30]; end
            10'd447: begin conf_c2h_d <= w_out[2][31]; end
            10'd448: begin conf_c2h_d <= w_out[2][32]; end
            10'd449: begin conf_c2h_d <= w_out[2][33]; end
            10'd450: begin conf_c2h_d <= w_out[2][34]; end
            10'd451: begin conf_c2h_d <= w_out[2][35]; end
            10'd452: begin conf_c2h_d <= w_out[2][36]; end
            10'd453: begin conf_c2h_d <= w_out[2][37]; end
            10'd454: begin conf_c2h_d <= w_out[2][38]; end
            10'd455: begin conf_c2h_d <= w_out[2][39]; end
            10'd456: begin conf_c2h_d <= w_out[2][40]; end
            10'd457: begin conf_c2h_d <= w_out[2][41]; end
            10'd458: begin conf_c2h_d <= w_out[2][42]; end
            10'd459: begin conf_c2h_d <= w_out[2][43]; end
            10'd460: begin conf_c2h_d <= w_out[2][44]; end
            10'd461: begin conf_c2h_d <= w_out[2][45]; end
            10'd462: begin conf_c2h_d <= w_out[2][46]; end
            10'd463: begin conf_c2h_d <= w_out[2][47]; end
            10'd464: begin conf_c2h_d <= w_out[3][0]; end
            10'd465: begin conf_c2h_d <= w_out[3][1]; end
            10'd466: begin conf_c2h_d <= w_out[3][2]; end
            10'd467: begin conf_c2h_d <= w_out[3][3]; end
            10'd468: begin conf_c2h_d <= w_out[3][4]; end
            10'd469: begin conf_c2h_d <= w_out[3][5]; end
            10'd470: begin conf_c2h_d <= w_out[3][6]; end
            10'd471: begin conf_c2h_d <= w_out[3][7]; end
            10'd472: begin conf_c2h_d <= w_out[3][8]; end
            10'd473: begin conf_c2h_d <= w_out[3][9]; end
            10'd474: begin conf_c2h_d <= w_out[3][10]; end
            10'd475: begin conf_c2h_d <= w_out[3][11]; end
            10'd476: begin conf_c2h_d <= w_out[3][12]; end
            10'd477: begin conf_c2h_d <= w_out[3][13]; end
            10'd478: begin conf_c2h_d <= w_out[3][14]; end
            10'd479: begin conf_c2h_d <= w_out[3][15]; end
            10'd480: begin conf_c2h_d <= w_out[3][16]; end
            10'd481: begin conf_c2h_d <= w_out[3][17]; end
            10'd482: begin conf_c2h_d <= w_out[3][18]; end
            10'd483: begin conf_c2h_d <= w_out[3][19]; end
            10'd484: begin conf_c2h_d <= w_out[3][20]; end
            10'd485: begin conf_c2h_d <= w_out[3][21]; end
            10'd486: begin conf_c2h_d <= w_out[3][22]; end
            10'd487: begin conf_c2h_d <= w_out[3][23]; end
            10'd488: begin conf_c2h_d <= w_out[3][24]; end
            10'd489: begin conf_c2h_d <= w_out[3][25]; end
            10'd490: begin conf_c2h_d <= w_out[3][26]; end
            10'd491: begin conf_c2h_d <= w_out[3][27]; end
            10'd492: begin conf_c2h_d <= w_out[3][28]; end
            10'd493: begin conf_c2h_d <= w_out[3][29]; end
            10'd494: begin conf_c2h_d <= w_out[3][30]; end
            10'd495: begin conf_c2h_d <= w_out[3][31]; end
            10'd496: begin conf_c2h_d <= w_out[3][32]; end
            10'd497: begin conf_c2h_d <= w_out[3][33]; end
            10'd498: begin conf_c2h_d <= w_out[3][34]; end
            10'd499: begin conf_c2h_d <= w_out[3][35]; end
            10'd500: begin conf_c2h_d <= w_out[3][36]; end
            10'd501: begin conf_c2h_d <= w_out[3][37]; end
            10'd502: begin conf_c2h_d <= w_out[3][38]; end
            10'd503: begin conf_c2h_d <= w_out[3][39]; end
            10'd504: begin conf_c2h_d <= w_out[3][40]; end
            10'd505: begin conf_c2h_d <= w_out[3][41]; end
            10'd506: begin conf_c2h_d <= w_out[3][42]; end
            10'd507: begin conf_c2h_d <= w_out[3][43]; end
            10'd508: begin conf_c2h_d <= w_out[3][44]; end
            10'd509: begin conf_c2h_d <= w_out[3][45]; end
            10'd510: begin conf_c2h_d <= w_out[3][46]; end
            10'd511: begin conf_c2h_d <= w_out[3][47]; end

            //----- w_x -----
            10'd512: begin conf_c2h_d <= w_x[0][0]; end
            10'd513: begin conf_c2h_d <= w_x[0][1]; end
            10'd514: begin conf_c2h_d <= w_x[0][2]; end
            10'd515: begin conf_c2h_d <= w_x[0][3]; end
            10'd516: begin conf_c2h_d <= w_x[0][4]; end
            10'd517: begin conf_c2h_d <= w_x[0][5]; end
            10'd518: begin conf_c2h_d <= w_x[0][6]; end
            10'd519: begin conf_c2h_d <= w_x[0][7]; end
            10'd520: begin conf_c2h_d <= w_x[1][0]; end
            10'd521: begin conf_c2h_d <= w_x[1][1]; end
            10'd522: begin conf_c2h_d <= w_x[1][2]; end
            10'd523: begin conf_c2h_d <= w_x[1][3]; end
            10'd524: begin conf_c2h_d <= w_x[1][4]; end
            10'd525: begin conf_c2h_d <= w_x[1][5]; end
            10'd526: begin conf_c2h_d <= w_x[1][6]; end
            10'd527: begin conf_c2h_d <= w_x[1][7]; end
            10'd528: begin conf_c2h_d <= w_x[2][0]; end
            10'd529: begin conf_c2h_d <= w_x[2][1]; end
            10'd530: begin conf_c2h_d <= w_x[2][2]; end
            10'd531: begin conf_c2h_d <= w_x[2][3]; end
            10'd532: begin conf_c2h_d <= w_x[2][4]; end
            10'd533: begin conf_c2h_d <= w_x[2][5]; end
            10'd534: begin conf_c2h_d <= w_x[2][6]; end
            10'd535: begin conf_c2h_d <= w_x[2][7]; end
            10'd536: begin conf_c2h_d <= w_x[3][0]; end
            10'd537: begin conf_c2h_d <= w_x[3][1]; end
            10'd538: begin conf_c2h_d <= w_x[3][2]; end
            10'd539: begin conf_c2h_d <= w_x[3][3]; end
            10'd540: begin conf_c2h_d <= w_x[3][4]; end
            10'd541: begin conf_c2h_d <= w_x[3][5]; end
            10'd542: begin conf_c2h_d <= w_x[3][6]; end
            10'd543: begin conf_c2h_d <= w_x[3][7]; end
            10'd544: begin conf_c2h_d <= w_x[4][0]; end
            10'd545: begin conf_c2h_d <= w_x[4][1]; end
            10'd546: begin conf_c2h_d <= w_x[4][2]; end
            10'd547: begin conf_c2h_d <= w_x[4][3]; end
            10'd548: begin conf_c2h_d <= w_x[4][4]; end
            10'd549: begin conf_c2h_d <= w_x[4][5]; end
            10'd550: begin conf_c2h_d <= w_x[4][6]; end
            10'd551: begin conf_c2h_d <= w_x[4][7]; end
            10'd552: begin conf_c2h_d <= w_x[5][0]; end
            10'd553: begin conf_c2h_d <= w_x[5][1]; end
            10'd554: begin conf_c2h_d <= w_x[5][2]; end
            10'd555: begin conf_c2h_d <= w_x[5][3]; end
            10'd556: begin conf_c2h_d <= w_x[5][4]; end
            10'd557: begin conf_c2h_d <= w_x[5][5]; end
            10'd558: begin conf_c2h_d <= w_x[5][6]; end
            10'd559: begin conf_c2h_d <= w_x[5][7]; end
            10'd560: begin conf_c2h_d <= w_x[6][0]; end
            10'd561: begin conf_c2h_d <= w_x[6][1]; end
            10'd562: begin conf_c2h_d <= w_x[6][2]; end
            10'd563: begin conf_c2h_d <= w_x[6][3]; end
            10'd564: begin conf_c2h_d <= w_x[6][4]; end
            10'd565: begin conf_c2h_d <= w_x[6][5]; end
            10'd566: begin conf_c2h_d <= w_x[6][6]; end
            10'd567: begin conf_c2h_d <= w_x[6][7]; end
            10'd568: begin conf_c2h_d <= w_x[7][0]; end
            10'd569: begin conf_c2h_d <= w_x[7][1]; end
            10'd570: begin conf_c2h_d <= w_x[7][2]; end
            10'd571: begin conf_c2h_d <= w_x[7][3]; end
            10'd572: begin conf_c2h_d <= w_x[7][4]; end
            10'd573: begin conf_c2h_d <= w_x[7][5]; end
            10'd574: begin conf_c2h_d <= w_x[7][6]; end
            10'd575: begin conf_c2h_d <= w_x[7][7]; end
            default: begin conf_c2h_d <= 16'd0; end
         endcase
      end else begin
         conf_c2h_d <= conf_c2h_d;
      end
   end

endmodule
