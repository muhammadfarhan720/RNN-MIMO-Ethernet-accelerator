

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AxZSYlrqWjjbM/ghGgP335GwqxDgV3HmMQL/p5ebckAQyJ+kqJFTPj58BKjOX4mpdCMv1bT58Fu1
qGdZGqaeUw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EIaioRFBcSeMA6Aux6hZm/WyyYgPDWVHaRtKbzIwL1QTiiAUZlNppzkL3bbmZ6KUvAn+f3bbBLZv
nI1at70553BjJ/f7JWSLFqvUyJvDaz1fb/ElTqdB3VheCofSfItuLq6wNAf1eaXg4UAiQMs6nSeP
bYv5xrpdIQrLt1D9QHA=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mb9yHUsW7uBsE4c/OKrF7NiKsfxXH5+bboQS2NnscX6YeRYxm+eBZvwT3PSD9ibYiQFnSx/solW3
OQO086UdWxyqMUFLcczGEx5Tqo5CpVbQ3CRAT7KgWnfq3Sw5pAuNsxwfXjN6luLSyUceI44YWnvZ
jNzoi8aSibopmfyW1ySUElOtnOzAOOsZpW6FBPVqwSIV18HJmOORpq6HJ1huXP6kFt/P0LgI4KNJ
0SeFy/2RlRADetCrV8umpxarjaDfW3dkNCeZIu0mWy7n8bNc/glh/qa2/i5v89Lt3neYjpa7cMXy
ICB4vX0zyiAb1G7xomAPECN8BfyzZeKkXU3L9A==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gBaQZNFSH7Q+cY8yvr3uGZIme+w3oCQPu8RtICVgaZhAcjEo9yTTeID+H4cca0yFpRdgM0pcus5J
5FJKmqOUXCBailX6awFdkRbi8P+qzd5LZWhXxCEFoQCAWDXZdantxf1Npl2sva9dLV8+XevpyvWw
na2fAJSEp/lWg0rNz+EcKnd11hmCw3Uq5A17kwqrW2kIl8yBpmqhRpwTKUaeyi1PlK2yMzLkDSj3
g3L9JraXIHucFD5JDVMs31PKB0bLhp9xva2XeqGFDomux1ArgEU2GMtksKuFBZYWi7EM3MnZ/210
ICkCIfO7B1+tuTs/vDrpmr16T/pcZfWjHD8i4g==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
X/0WESaoHNKE+VQh6wiFQZUGC/wvvLyzJWa7+XHLf9u2HGK/wbJysf+svmnB6pdyOjRcvCdqkITz
XwegHvpEnCL5eBSM7wrkLdsUEF3XcNtNuFXLtFkrk/zKPfCV+Cj5+TdjprdgEEGSQyiJEbOirUGo
QfOyWo4Cn++z8sGq6DZemWplV82dIQad0OMeak7WWmG7Pwef65b49WpZp4VtkmzU6zP3Hq2RKuc2
JfAEvP+4m1AKa1AIvFYtKkIno5azYqCR8icyJj/aAeFkwKgmw475EaivMmiwXI0CEGgGhUaSatGn
t78rUSYMEB8FycWJ+tnZkr2fLD603a+4Ea82kA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y2sBFuuYPz+gbw4FP5O5GG+zlVJ0DyXBElOfyt3NhcumgiOFXrUdbEKBNszNLNHqdAfX83DQlvFe
dmRFhUTrp1zAwODtXOHbgp7OcQKFuaGIo+poJ6g+migbsS0N35Sw+qK4xtbAtXQz3HjATWd+gz+S
zCFMgvYoG1+WYEUj2X0=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sOc8FhbMR64uyLpKFyrXkbouaX3PkKiNHTHeAKNeDiWbDAV3jythTS34N4HWRYzf/duBai4EaRTQ
3byQC47/ahfN7MGuftFmc033WhoNzsfTJkqu5w+sXclPKETCwWwBGCfd6WDcYwA1EaV24NgJqZLO
VytDboZOGxpfIwB2yEEPyqHZQZtat4wiSyi5mDJ0GF7oPhDS3s+HLx50a1i46WdrdohQl2WaD1sL
bzITraqPIVbRdj8G/0aABIIWM19aF6l4O+1DKGIRw/F86DxkXKS+zA6V3SGO7M3LwyGSWxhDz0AL
KBu6Yul8QRtuswKo8lHHQeNt5xF8Z6yRrWyGDg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 132688)
`protect data_block
Qo+8CwaZrt9iYaUQz+wHitsLoskg/dNlAWkcNt0ujtMwCgWW1nCQg8w6VJ1u1loezzUA01XaZ1IL
IRoNG9zORqySb6/HmITpyw1f8GXB/3fYn/NVfRSgoPHX2pG8KwFgmg/UoIQO6rw0TISlQAKTlkz9
Hoe+jI7UaBBJMYm/eeQ6C0XDTpNQD1lkVqcYCxsyn+XMffeRcKvjdlKw0mQKhE+PlschdvsbEhts
zPxOy+Wjp+hwE4gkFohbTonRvNmNAkonzgh7bgLo2RZO1PXJ2GsuOJlrYAurTiB7zecZcyHvXVGS
VQxGP1QVzid/HT8SZ7Tggb6VetY5zCvqd/9f0nvrm+BxiJYct8mSAbu1ZOi50GWCAJF+RhKExFxe
7Hb3mJoib84Uqzz2KSrh+hBVkbxKSWdNb80Lvc1GLBHJwPEYklKwHb+CPjHnJMUJ5atwR5uSzGcv
Z4OHDDBApqzP48uaWsv2H5LcuaWgVbbecJ3Bw/vr5vY58YozszQldVIgwt607n2/K4Gt7gHqWkkw
bwvpQb4X2j0IevMOLluA7/nLFuv/ddZ+3Fuzjm/VzLRjb/Mp1fHd5EwmVy5hqHiD0qmAFJj5uFt3
McJ1VENrXjh7xRVIaqh2/UauRKmkJOmgU+xx+ujwscBUuRKAAdKBXa2jFMwbucaG9KzvwuEDsDMq
ZmCAGzB7ke3xbJQFOMABLeHdgjtVwUXsRqCuNYOuU37+PXJBOgT0LrhFJ3pmX57cMnXEwPAk69Bq
ITZmQmMhKKxzmYhs8yiferAdRXWV+DMPmmg1CuFEp0ekIuONie1M3JQytYSJ6E1yrcsckdhi5UuA
naijHAerHsn35x4+qD2kAJn0T4XSaI58b3HRvle823M+q9M0Bx5ujw3GUHtYw8feHIiMFloVYrBD
Rd+ERKm79PovZgw8ttpoxwMNxp3VxO8pQqWyYekHDz0aTJrhYXXZlqktkwScWKrJMdTY1ljkeOjK
uEbalEY4Acm2BpGvuh3yKMvz6Iu0X6ESaS7tOixyurb2arPNyKxwg3/oeZsCI3U0uPiWkS4i4TQ4
hE0JyQ7V52bexhylYfBJrIiTYwE8axuqYShDsl0xNlj4gXTfUFzMhuAUZJe5xNKemtiOr2yHDnj/
hraH4Vzy+CUFtL4qjsiJ9nebb54f/SfdZJGVxv6z++6XscYjiDAn7WyJ0uYx9TVQbQEqlbj91NCN
Igv4fodKUdPr6xjS9hKcOQSArmo8Q9H/zVez4xVXP4Cb1vrMw45GidMj5fv0vFoinb73YXe1X2u7
2UKUuzhxmLTHBE76QpZGQTa85OoPwLVyupoBPw7He+iDXaoyObREoInoATZlrDSeXCSK5UQrZTGq
UEZ8zCzLGtOt2CgOaMGskTiL/+X+px6iqF2PLTdyuB/Q1alobN25vW4v8BPdpx3Ol/aDa4QA7/QL
jQk5uK3grz9ms6gVNKXQ3R3B8wo8avlRvS3P2c/MQZ8yu8Sm9ogO8hWYYIpELStf91AJq//Htq7i
l3ulIZy5yY+SL/zOSxAj1snAHHkvsy0XDS4cx0H/eOLO7YSEvdWOzgDgVjlPcrII/YBTPYBXmfgL
VKgsyCb13624U80+/A4Rew43wyGjXXq/8IcQloJgncJgWPykbbDPFHnSMu8Wbcq+FrBuimqIp62W
meeoYjjFL+zpVNnHgvvSO6g7UT9hf1xevfjo3fmydvjeRYu1a1x8eEZeMVoSfMtApYHSJhz2Ll97
YedIGUODjnXVh9+7YCFfeUFqLtMX1SqFbsnDm8nflh4OtD8PGYC9qqoHp6l/boI6NrCiTo0eIXy/
po2NeeDLd9j1qe5Ei5oeLRRhtjKxK1yUtF1pEdLNKvLN+mcd7k1WlXjn3QIzuT9+f6gSmfqs/7GO
kkBYTtcdyYapJ0OiKrYHX77ZEwT1UaltzDuhhmbxqI8vyevtr+CjJOuyikAaBpI+m+iNdgtqJTjW
uPzhuJO7tQC/6ICaiPLVdqiqDa8OtdDtgf6nHKHD4u8eT2tqQbpRebW2r2CA8BB4YXzU1bmp501H
xu4UMm3fd4kc0eFtKKOxYVHP1FOWgwpAlFyRjRe0YpI3MTVvYVy01BgQsKb+0Jx1lLwUZCAVYM/J
hPmIsp9m8wk9nAvk861e+Dfn/J4sVnf2MPx8b4OiYFcyL4IaSmOBrWztts2Gyi8X+eLdnim9q5vj
oKugegZoxINwxH83TFbWQrUOni2Y6aZHepLZA65Il7nN12qll2dBa/m036DVP2iGsJEsH5QG/qfe
duvg15AsO+43ewYe3bfLm2L3jI8mz7lSII6OMtdNBRTLwKvvcZD+Laa2P2xptJHm3NP+fjJn9+vS
8znfkubiXsP2oalagqNhYD1B3oamDfUQQV6TnRm2D76iiVTb6/RFh2jueDYtaipqsPnXQlTmPnNI
NL0XRiy9ByZ2g3mA76s4w6SDAgL0QAAhlUiYW/5f+x4Ln7JWvCZ9PniRpDzcFvwQ7ajlO3XatOvI
7vw5v4dMH0HeEud8/daj4q2/mT1iUDVHW3KDtoUmnzYVJ4idR3zpA68fqOpa+SSnTWmFH1LFMzPe
wPwHj+wTQBDRc7QcvHzZ9AIJKJG6vQtGeefFnkow4z8YCQelioL37vMHq1QFumse4uGzuP0qEFCm
4opanXw0cUjs3uwoioA1alTYfIuECjeJFqJkemT9zCpi6RuqVo/3rnLE2Gp2z0U6RSZ3nsdbfS65
QOL770+OvnrX4Z+2D1lZSX7xC2pyz2raQQgIGuRLip+2cK+/5TpAEdh6D5ngZGqo1qE9hZKXq8X9
z+Sy5JaFOeZNGWFTOvaf3L0Ahksk2+H6B+qUmEsMspyP6txk+6TDrat2T8e9AexcSpKpY37s1zYU
jfORsBk7PwtTAb9Tcuf+JCWFXb6Au272K/1r9o1VehlEQbNUitMOKIpM2dsz1wAxUX3L0e1pYMys
eRWEn7u0ZvRW0onuCg/en5OxNxMEiu1mkgDfQOFozswJdSqpaiZgr1D6Tl1Y8SlF+Mwd4Z7Wpf4n
H7fhsFnzHnIYwHdgKDHpTmfEFfTpsKW79xGI0cwPjyoSl0r1pf3F/T0XkhjSaWlCAtFaPU4CSdDC
dGFm/8GCZ2v/X8/kHGfQSb15f0eNUhqyRPhAxnb1d8HFN34oJF3yJCMVwoydbzEt1OfZT6lodZ+1
HNGefp/BimaTr6D0Q1SRVxbTUTIiayLhyt13SY4UKwqNpNO/Ye0p27RmZDcd+YWuJH+DKdZfl/O0
9zdHAGtNL0uJ/M9BkETdxnG/3DTc2stZSdjgRK+oetiE2w/M9usTMSpDWDNfW5X6Pb0WmSFBS2O8
Sq6GaN7lf5ZoftGsLS+bXNBkdptR7amAXZK246FAxpKhTYaklcVFg5qo/pZXv0w5xsOawluNt5GU
metIY8v2nq1yHSOxGsCmGQXodg7IHR97b95ohI1JyelBMRO+aRuzIDPCaMKkxSrhzURWWGiuoLsn
rm6Q1iZJ6vvsvloZTxI+VOwssb963GqvODpYNLxqJKkx/xEskwDylX7LY0Tsag/eYmahSjio4M/P
GxkFd8XAIWDUcZ/rHy0hMvjXsbhNlhajhKzHS01POevcVUXGRaQe8g0tFrbXeBDMeY/WZurq1Rnw
VfRa0sUv5fGtR5z4dLm8ZTcLxcT8+hPZKDoouy1V5ByYn9AVTCcF9/dtuEH7vyIY7oeXyXVVATgM
P9NcelY4Ne6LNFuvyyvRSUtKi6HeXYWD6NIx/MMVZskcGp22f+490Baqr2RsEz0OwltG1Mr0tXRi
VZCWFpQSrUzkvGRkXj/g0IFxHcEwFVtkvmK12hSzBOYih8sUoirFbQu9r5AWhzsHrsdZ/vyJl0Id
VknF5863aB5Ok4OPVLpDLwFsEGTqwKhQzFQbYciXp9/6+l/JPGQdu2VlaXc7MV9ieS74dlc2nYVD
0Kw5Hsjq2qhPx3CmK3ipL48r6jE/CCwHDUUWMl+UvpBqDfIhQfNAvIcxuFLwYx84sYFtaS9RNzTB
ol/TvjWGjGjZMezHfP0+uLfliFcGoXnFUZuV9JW89qaoX4eOmGlUL4/V9Bj6R2Bo6iQqfwRvw1Yj
ath94eSHungYzycOPgFA0uw7wolfAAuuAMzxjGy8twlFM2NI3K/KqrM5heUSYjUH+4dYNPQEoyOM
fLwLt+M/HqO44+CdNuugpQ/+XDiC5QGURQcGhtn51lk73DdfiYBE3wVuSFGNIQDUcdr8mU7QVatP
lV7fxqGZyO9i4x8S7tDGC1CI7KbrYNYtasTeqFXeUOxCIAW9ZKn+BqDdC2UysbYVLb38Fk7ghKoS
I12ejyQnGHd7+4t8a5ynD2ePXHMLAhbnXurCCvTbLO27uajOQJwJlL/DCVcb97oiQSKx3lNZvSQP
EumHpRTEWXwfOjmS10nfTvum/+sMTCeMP9qI8RZ9eYg4xmsCeAVAGorJrT3TP/JXRLuq2Gj+bz2X
3QfXqTsPzRRU5dzNPp2NU6ttgHjpCe8TSn0b8vNxFnmm+LqyKcAimR/I5x7K8wuZk0BbVk/z1IdQ
t81+kdJOplOzojbq8KnplkacKdztM2qtUQYCPCe9RtBnMuhso5YgPliZyvCrkb+u/XKYI+1n5yl9
bvq8so0MNJw9toKTxB2RkCrEhFk9t41f616c5MeiW/Hb8lVTbfvnugKyFWxSDzC29hadwaChGtU5
HXZGO4Fu6SdpOUr+Gsg2zywNcyAu0IkYVF1ZFMAsnYUeI9hkKj9co/1hF7DfMsJ5/m7FrjJNfjUO
wday4Nn/egJimfCtmWYMbcnEv7sIo/P/D+sjn/YT4XD/yNSUlRJfYacQUIoB081/XKK4wkoJBnuM
rHHuZLmjR2sTjQQlRsoDuh6Ls1JR6Rur1CiM8B1PWHGgtUaFKWXJ4/UqM6GN/KLQD6Skg6Ele5uY
EnCaYyDSSv0FgXG5uidRlhr18de3RyMCT9OEvLL7p7f2VBvTDoMG1b835Srr41DRAs1Gso7jJqB+
+f1lgOB2cgko3qAhehu7AoLQi20i0Xpry5C2alUAWJZm+mIT/LE8qp8M5YzzWMsLG5cRvbAocYhq
OEvle0JiiVf97g8VxIhw5lYJZbE2amjGA2k5G2UDWFBASjdBCj2Bde73cuiTQoexwUvrckm8TX/g
oh+zR5Z2rUsps8VLRouaczkJrP07fOryBlBjc4MU6a2c4Lr/HVQ0D4BDhkEoz5AxCEYXbkjSMJDi
guyIn2mCQFYv9ECW3kBTcxSyoDPOwcjbAPZobyLyee/9tnXmAzfWuNwAwTVe/EnxMsuYOXQ3DaNw
HC3ezF1DVC1fMQncYn2BpcOzSeeSipc2ikBQU2MovF3TK2DpHhmCk4VxKGkkcrQHe5oqdvvipx1l
TMiCMrXYih8PC7oliKVGakV9lzgZFWAlySV5cgvnuKMBtD7i3u2o8XGUTNxebxsRJ5tDzKMNfCuC
3H4shXHMZFYNDeRxCUjmw74Q40tvWkI1aSfumqiLSAn47ieNzRe1K8jErdDneydQuAyeGWkIH6DO
xFxfTD3cIFmMeWQEzxrr20VFe83OWR9NhUasb3SYYffd6cz1N65lEgYn7TUYHAgOCKhmxUCjqwZE
te9aKr7vE8Znng0AiWv7UHw38Z8xP6iY392gkXuUadmxb/An6vtmZwC/lMLQxudsh2ZGqQrHCOoV
ZZ9Y20I3HDgaT79y3VeNaUTRdPdgT+RrDv7MJfo1KUpNKuy53J2xF/QbVNXvDbQ+15FCZ8MEUixM
coyXIVBY77udhJ3XpkD9CsZpIzRKhMs4izI+9Q8Kldu+8rwehNWcQ+jx7pDbA/BHWPJhQOow9eiZ
TzMsJvDTfJHCYyTOsZifvZ0/YdFhQqFHSllFFMfRP/qv4UAVXHEMQJAj6Ee+LBTCldblYNOBoMbU
/hcN2ZtFejzlyD5Oy+eWIw5Pv33ts1F1VA23l+zAIIJKOs07nUVnBf8gGAG4vrI8Rsdt2h0wNDZv
mnqCL31wUHCeQly9LQDgDtaAC5PbBalALcBcXrRp4FHQvWEqdeG3SsvSO0Gd3ykzwzKPjli1oYiB
pTpSt8aCvC2cz7tAS41gN1SaPzk41E1dXjt5+bLtKWuhSHDGzrZuUUFFZddH63juQyxB9pD1AAxO
i6E63Vf4veiA1n6etg2gcO+9v9VFhCxM0HY8YymerPtDRcQTzfo/aIjJGZzg8jnMYpM6w1IfhdEL
bUcmPc89j0NeqTq6zEKf6Pjy8fnSF0VubitcGAUXqkrn5bBLwNGkXui3ud2qZ/fxEhb69bV9hVbj
F2PiRhc4xs6m1RPQtPQOpymG1g+DGrgq21Me1RTQWmkrElGu4JUfkIz+WGVmjCzD8i+/bnaXg2TU
dxB/T4w5DH+vtEmDHiG4cBAlH6GZslBvzSLafYDuS3TxSpTYwqMf8cZehCZcmqbGiAwsVQqSLEH4
q8UACtBTDsh+AhwyNVK6D/EIX2FeUrih9YK0SHKu11jLZa/W6eQZZsWfiXEw9cMzWlC4rPqA/oZR
1yPsZ+itY9VTZeXBliEclQN5DbkihboCcjbHI2IMr2SpcoW5LUo/vSPY77MrtB40mGP33mCI0jbY
cxzZGVTRN+RwNURKzeH7sl4U+NOPvBFaJJ5LpcEMk5uO9ogdRxrFJmyKYJB2drPOUn6UxI812uHW
JdokpAWC/zFWxsOIxdioXceZatv2q97U3u6qtkWUrEXMI8wxy1w+lT57s4XbCFCugpMbWsGl8Fdc
8YnbOBdwavfpt8KnLnNEEqLbcNDUlQU6yIMj18QDrtASBSbekbNR4YwUMShN0R4sWKvtDAhS8sAm
T/L1/rfojKV1BQXsdqTCnFZhF3nrvP1qXr2JetMTyxCb660hetkWpuMNxEgRYBI2zQryy9h8fPMB
07f3b5tD5DVDUpsYTDXb9sgwSgzdYXVS28kvxIiES0lNtIbR9JR39TH6HnqCIHpNpv6Ydk8NTF+9
R/C1lmHCTxJcorg8KPAd6dLk408R3K++xAlFIUU4Xb8rrYZyMkmQxYvPSLy6PS3SFa+jTPt3dVoQ
nrjJ27W1ECAE/KzbtjF60LYQz/YKI2V1ofW4RR2FLvWGePzLJmkNzIRMVQxCU5Ck+eQO4TbGWo8z
NjU3ekc6q0dHJyNL4ojK57dYIiuZhLmKe8BDjKp1Caw8nC9nw3brMRlXVIYND0GJZLSXTzP66/8c
ynq4EYlNj9zTjG1FgcSNPAnkA92Qpg3yl/SDu5Y2W42NL92kHw9zXPGC2N6Lm8WRWW5fFOfBaulF
Nw/t4hBentsysbWclOEGJks45kg4SS9H42eacwQHiRsPqHELPuYTSsxMQQpYpegAvMUclNyiH0JT
P71NJQUVBkDtqUSv/PyFMkXZd2JoBdw3rT+2hLpSfVS7n8PJYpsCQmWlPaVI9bHi15ZN6sT778UJ
mWG/xHGe+xvb/OvdAksJPTH124XGgwMNwEUoeuScVpuZIP1+gdpdSDNy+Lbw/OFOmkajqWS/Ebeo
1einF64skfOE6a0voRa/G9SSE0eTcKIarsnl1B5cKMVgkeqtwokLpd8dnEUxaFYwUKcQ46u1gnVt
z1sD9WeH1T3MRdIDor4/zuuxXjViLv0B5qa5YpSZ4F2vdhJpHiojIuJf7LFu/8vxZhjyxxH5RYBN
2Qw3mGCLgckp/faGZHmsk+p4mbOSItIbxnnBTpRdA56pF9mID6n070A6fNB163u4lICHIH3dTK6/
MurcJ2BPmifFiMGQAHM11IgzQJ8jQCeQO6bz7KIManqljB/4vixih3WNRIGhayy3GZ9GY2kJvG35
2GVey+yVUhBbV3vgHnPESTDJjO/OcHFAZmqTLaK+Gxk9o/i/I7uXoZQDPjYx8K6Bl91c2Lw1iEaG
rbMXqOBhI9fN6O3quQxRFPLTIKkiaPRjissW3E0e7ENYYKu0CK9kKjlD7aQGsdda++qvET71vS5j
q7UpFKI35lHuSLbXtqSzzcXqBDxx9EQHDjLAenn2hjj2WeHt4ub/3yTD8OzndVm2aLtrjmUfZX0u
O9tRG0TUoi5tUGr9qdJMkkuOfi3qLGk1lTRON03YS2z2RRopt5JmJ6ky3hS0xqkRQ3vI54ZTjtGM
Mkq+ZFLAOozy4K2EOcl1NKrIi3Pbrul5UeoIgHAowTc4q4b2q03MHDTA6Lvk1Y49vfga+m68Dgru
TqEzH3it4Yxu+rHw8zBvsNqjPBI5UBVWUL6HJiVFUYc5GJCucvYhFXkjR95xRTc+sLSMnUfJ+9WN
LV9rofWa/b3QvgVrmESZ4dTr80WcddW/8/seEQ6zX1ZrnFj/1ew1hBrcF2zLP9UXMten4AJx0Te4
TK63WMQThXYJvRSCAPgUwQlVOGKFN812Gv/94tg31R6Os6qji4BKwdimmHaoXLZ4bUw6GmUpB59S
vqKrtQCzPdMJrIr1khZAbzlYSQ+EU9bA1n481lmdiSZHHWnGLqg8M6dUbq4kutiJVZM9yrAHTHjS
50epy/IMZqqvDtkxIsY1UIhnRD6qN/SreNdwnFhZ0SWKvTStdH1AadShwxAGgkQfUTmjKmgFicgd
dAUpCvjV42yQ7nM8KCyPUZIZp1YQH2ai2HCk4Y+Ks+tzwoU3u793I0FTeFNuu4tN+WHIC9HeR6eC
HNlNL7aDTwB+TbWIIqrzbiPsqnOJE/Zs7RGIJBVx1+yJU7K9dPA8zJHj7gnec1poN0maU0dFam+x
x/ANh9kLbm/HVQSmkyO5ZLQQxBPQdvAme/iw38pNNnmmFw8lK27xwuz6FT+ZzzE4xB2q1rMTitoe
WZDEhcyekbt5xbQ16lsD25QJjiyB82+U9RlrOJREX/Mt1jvED93BFuKGE2w/q4k7ZVVGJO8sOIzf
MeewsjTDLCnY7Ejieakcq9RqqymcWM7fE6DSzOy53V277CCAtOb5Wx/GHdMd1MMCtxT4HuJvZCC3
9spqxmrCFVdrTGWqZ8HT+/nSzgbyEKbd3sx5ruZUSBK+7zeXaNxpTQiz1QwzEBmHgmYTBWu1wzjw
P5UtG76hOPr/Lnn+kD+NAklxsSB/8cyUqEnyNVdcrTfUlWnTQ8/1X/nx+vnhJKvs2oih5S7zQ5pA
GzMvkQkchvPTICNfD6BfNHBMl5YxPOd/Dh0FC6aK08c5S0UuR/chn6Fkgyka/YFVLGIeRNWkykcV
r4nSByeCbbXTVbr+AzQn3nl/OFSWbHhTvz6+KQ5dGW+GRRcjOSd2SvuHEHtM8X9jHqwZP61iI/nO
T7PxvCoBLYIlXHtgatS854Wjf993HSPxaTNizGVoSR8drnGTQf8flmeQmOtUFpR89GtrAyxkPfQb
HfRNIWc4dLBYTiPmOQS4rGOEQzUkzpQSsZfs582xuU/RF9zXm+BO5bOxjtulIXOXRFQ0NhLLQcff
eyuv6hbOKxzxgcAUbDfSkdQxB7FK6w7FzowezWsZHV240qEXzEZgwcsIXzdS4Qjp6g4G1zA/gNQo
DNyypTxZS2KfxBEPF0K2+q726aEJmBBLjUHtShkT6z83TjTI8/+6i1E8KmSDmdJb1Z62uLynjfQ5
G8OmgoiDJLHsRBZGD0PZr3BPTPJHZiXDfMfaQKIpLmT9jk/pIgskZ2OwGqTYmO9iSHkmntJ6WrkG
juMYkMRmTFWvhCZpceJY2iOVHOcdvpIiDWw8ed4iw2XX+ruYxu7lDvHGuo/z5V8ZiEKlNeCgFnLC
hvuZkPNPA3tKJ5XuMbhBTf3ug2HiFrQa9WpjJOCaQhLUlmStmHNBkMvrdaoah6Cub9m2XUTOtfTa
/n51qgDKkvZRmNItM4ghVWcEmRk0QmL0UmtaXI2jbukScZpJLbZZOCUn3BhKa0LBMC75jf/LxEpB
uFOyr3KPb6cTVJf+EipTzPngTsUHlQtjDfsgI8fQNDqo0dn7c4rLpsAopCc1umLBb2ZGpMkJZ6A+
G1J/ST+3o2DvVXzUEoOBomajZP9cxzFYomeMVSFK52EUKZghJdAnTi3ZZSZYIZSEQosNIscsAFd1
vAlkT3fJqkAKABA+HFArb7eUNtw941u0iph/Qbxgwa9xa8phdo80oD5pgAeacni9qd0hRpaB+oXm
X9CytXa4+eaNGReDEcS1J5B7WNwZsASGAwV1Kz4WQXYPcl3XRbqCEUEowGByhtC9xpdVEPHnoZko
fOoVTDt3rSDw/V3IC1/wuWUnq/jVRNtV0noLezTIMbKjkt4CcR2cOCpaq7kOqgDblHQVt94hK0sV
ZP+rVh5QLILDHov5mMpoyqoEDNzqQe/NEzVk6PwwpMMWmr0+sutuRitUYMZLS0+obLe9FjJ9qUwV
GLg3EiqzQ6cU6isTlQslqNKrjljHWMbkRFM10w/7JtCj1joS8DfhjdLp6Co8nCMGf4aKQkKraBv3
PKjKy4FSXvY28oKwey8CVwgSPePGbTxqTfZDKVWG3xNw9HuYXBWrYlx2FHtkhjIMMTAqVm3j1va5
kpuXReCxOrbUuIqFObxNvWrrr2zSxbCE0+hwcoOWm2PrlFP1dgX7rWEeKxEUnCqqpZdwUq1q5lCV
j2RKbVvb77olD2orZAqTtRPpsf8gYjtaibdJd3ElWRkVusgTCxqVrkGE94G62UsVqDAes9tz2h/6
OyQAoIip2tvM0bIkBN8OhMcZRN4d5hnqauSpNCOzF1aqpLFbVpAtv9FC+Qwdd3WVAZf7LPB0wlpF
NToHcDSncOMq1zZOAor6HRr8WA62DznqWR2oFpkuwOw7wYHCqutUygvrj6hg/f2mbCkoD2roY1+D
E4fpEUhv9JCUoa61pHrPy1yhA8f3qrGo1ia2ahHdkj/AQxAZ8nNxpTaPeDhx/1M3eGjgZRGMAwrr
t/n8TqeMc4+nXPLtbJRa9hiJ3Ngxav4wAgWxbwpri2Hc/+Rf+HFI0KNDsEplx8tDfKjwV4SB/pa0
osWUMm5SMMOXF624Khr7Xmkzz689XAmF4IR1XtcZU7bdfPHN+8+GV1UvpQX8s7Q8cV7hRX/tZ16l
CBXfyv/+kLM98arUEjBaeTLPwg/2S9IDT8PuOqaK3+3gkydsv3pUMiKyXccDEnkhDYajri11uMNM
GHxkbtQQKacbBI4AH55Cwa3eHZ5ATIHZjfiK3RgH2xzE62UuIov+rcS3OodTkbjNPU6sv2iuS7Ip
X9b3BIhcXUkE7P3PY+JFUpaIg9Q/H85V/7az8I+wPaZZZ36etiXh+pdyD+Rd+BFM8731A16yprKY
B1bfT27At2Mc1aly+rDMQ1rHX3jFwmom19yLNUzhd2iptMwvOcdb0AckOyYtOWrtwDexqBM6MswG
zvDFRGLMoykC//Rlbz03TJWWiRRNsckc4Zw6zo2Lj982+0Om9d6U80O80EmhPM3z3B8qM1NVTm4V
9ETZigcp05FzJ16fvlvJrtV5DcFYwke9ufG4QD85l3mMrSu0/vBOSUlzfhU5NGVCRkB9kJqjUloG
P+ewIEbUMZHbCOLh6WXGqKhdrOFX3+BwNzDo0J2Z6hZUq/1+rXx4c0sLVB9YdTn/CiIkJEoSdg4U
amW/X6abBZUu2lHs9fqm2wRHLjCR7HtNhC4coZ2nH4wVypZL3wbuxod3OWVqjGWoXy+R/3bcd235
DS9G8ojdzsnOLqtKSp+inC2PRjGsqtWENrCnj1c80lp/kRXweKZYwcImvgGkEAHLEg3NM84RTIho
DGelPHwhTo/Ef7essmbS/0fasi3xrmi1fCXjAuNPLC3gNoik5EYmlelCUdq+p5d9c6ZVEh1ia/GO
dq7k3sgHaUmsk4eJZDlwNGNZNH3KJ/FarUG346MPBkzr2mQfjEpbJ+l7lPAV9xhmoIgo2m0kFTcY
jM04FlfHOcnRBDcrhA44M73ZG1vnq+Mz9aV/hk5J+zjgHbHTuv81y6ZiDJ9KUfBQcOq6IQ4CAfe3
mqbhwvylMoO9XWqSGPDYmnk7/HjQbU6DQZfjnwyYACQoxR3o9U+funX6IqGW6TiRFQ2Ia7EOpc+Z
IrTjvEEBk5dp8eghKSwpqrrHhquDcvIFg/fjLqhKVqPJ8tIwyLTn3vMco207sYPHSxzGPRFYzLEx
XpwHYiAkuhUCHN9m8OJGo6YuhPCrD1b4HnSXNubSK5EVoSBGtgz+Ar5g0mqC1fGQ7Ob1YqhjBMiF
2m+Kf610pwoF84/8tlG+IPjx3JbJaNl1KBHAJBrhazKZet0lLNa0pngpor+Z9nxGLbL1Ujy7RaOO
amIPvoUYMoS9N5Y5GY74UqLNhZ7EMyOwzg2H6FNzy5wN19yqCAGRjZ/e5wRXa4SkFktznu+XtndF
6BvFflVuLcMwYrTBFHWZAp8jvKc+WJW7+qwdTUg2DL53GG3gcCRUcZYGUttVd58PFSMLyGj7LAEo
FmmmwA2ZgyW8uEhQTKWpXv4wBwTKTbTHNzbufjESBTP4tPI0C1LDbbtet9jpNQt3GFKJLhyUxrP+
5C4se4eUlpz3WqK1kb7jeYkomBk4SrT1tmy8EodV03NHNdjN5z5eSYBDiysVUmWvQarc8sWqjBwk
gPk55tpBKbuCfsSImlZcbBuIh09bTt1tmqNL8j3rH9HkOGkkVXRZ9dbxFfFHBccAUwvsBdseoP+5
PEg6SnyONUXVuaAZI3pMiQiP1z4ntQpoRsF4Z/S6qonxzRMkhlhC0zE90bzkuxtEsFN34ZlLLPeO
QiC2WIqMltk1guCFXGoqseojElGdeli7lArpkAzm23JPJsjZHjzHzKOpJhyrlmZa+XTBa+poaHtf
ZJD+qSSIJlqSKy7NO0E8BnISdtu2sB/dLaHbQQud0/JW31DL5XzCNxgSwurHVmj99iqVawReWpgP
YcE6bWIW9nw44I/p9ewh+VAc5P0lBqdjJyp8Lt5DkfSdN0k9oe+uzssA2oA6R6lOgwMg0VIu/qKf
V6CqqpRf1QsK6foKbXS7i3ZgYBAOFaA73FI4WXl2JddIuQ/ynteXaTNN4eRLNa2+MT0tbWCINKwl
NGEGmDEQau2Qe/5PiARAlafeJ5UiklSB7Q0G4kEz6IvJhSv260IQKSMCirXjDmigjUcKchSExaq5
aJjfm7X7iHXpoDGry6Jwyqu4L3dRSsFZleo7SRFz6wdRH4EoSQbfFYMQgYpVCV5UhZWa6AP8QGU6
c51faX4SAk9rKTydNc2CGBk0vPKNaQN47yGahLImvVQZ+bC6bPorilTkGCDJzUIW/knB2UD2z+3s
IqJjfNnLuD/k73GVVh5TswAq0TXfXkwdJ9gOb7gYvhkk0aATOYmhO/xJbIWWORJVANjeQgjYAtuD
GIdflCp3z/zzAsucbhqRWl9/qpomGr+a80c0fX1mypzSxC3eeSqX0CmYRzXj7CWMvzlmpwgnuAfY
vYUUGpwkeTRdw3Beoz9iYB5WI6ZFOr6jw0uJc+Yj+DpBg3heeWWFUc7ojyGBNl7HZrnDSyJ0CRQr
Xs/EEaOBf7ugXHFnfaauDTr64Mx+La+ukuzYUjePlBWuxUmWKyt5u2/wUZ93ZC4Io0T5VCF28qSM
s+TTKr5eT6RsIHuJFAP0u5S2UzU8UXJkHPsMw0c+wucB91k/cXKTBALvuNf8QEOtdNbjzVQwLJ99
pzfxVyVm9Rr7iBpW+mN64GKVbBZ1SXLAB9jcsM2XMwPjAHqgW2N88+rFL7m+wiypUKO+6r7AkEl9
/miPiL3zMUECRbIDNygw6SqOeS6h+4TKoGWk8ja7wN9ZpKEVwQ/X+pZExpFZ4SsWzB624Q681CLw
9gduIWhcLKhRLrlMpJ6EAs+AurUxpL8MoadzGQ/+bk5m1HQnM6eZf2fBGF6AGqNC6qSWrPdybhAM
IE/KFHbqU086GNm2g0CT/qEUvtlaLC6yZRyOks4uLqHgW2GXDOjV7kgKFJ8V3V6dz8PzLusiHomU
qMpe+0laljQpiWoWlOV+mAjXPEKInrYMfEDcVLOJ1Ca8DZ5QCoNVz+i6VlqfjzUZn2AkkBdwRp/D
E9NqKFwR/+iU10W1ruiXzVF08W5mICZgY1PHnRreWIjWle6XlJgdGNYieaPpp6P9ESCyjivv6e5G
2RwcQ1EFxMqVYL/NHeRi3KW7eiwjneh1xe2u4r91o6n7zR7zuOjpPW7PpKGQbUUdbStT2T0w3Ll6
MvrtYEUKbsLtmMOn+cdwmld5Mh0mCAJbQH1CxY+Z9EbVLSnhrLUTEbjNFJ5ByIBZCwPTmcFlAA7y
Qy4hacLTik2CTC1f70/a1yR3dexNbwpd2EdSOxxqnQgxzxp+DdLNIiA+XNwzsyVc2rnA8PzZhhZ9
17lwurM68QtRKei7kQ2peA/RrVRfJ5nxgM9LKryqvXpGYkkY+jFHGpi+wIYyUQI5u9X0Lui1kNbT
pn6I0XJsHgU+XE5tYQJb6adPXHepnnICadkSU637GZ8lSgRzNroJJVVRljbcscc2PlhX2qQFKG6C
6OdHHHiTqFeIBFJgn+YDx3LqjnPV/QGRYLzH+JbNXiwYjhU3ZP12tuIlv0mz4Amnvt9GD9amwckm
taasXT1TTWcopaZ6cEslH68mBirAb8yGRXMA5EhPYnk2c8LdmBhLhbhOs+dlpzdORoXXAQ2GPyXY
DtnQaitZpeyF2LXTNn3duc8nwF/V5LWA6gxxcI7sqzPtQJge2Cce/UozLzFsLTIAxiC4NTF8/uaB
HIE3y81ENP9MoIjm5ZQ+hZBiau/4MjDeA2NK1crMU/AUZWUu/cRPYcYYLf5yICZMtcivc5GNjsib
A8pM+C9weyzEavBWLtn7fkRz/WTwtuUBd0WQKV4QgysSIvAcxxBHccuw0kr745t1Xiie8jeeTsJx
69hCDpPyzmlS1LrLTSjrfSzIjhnRR2naNQuW/Sj159ODF8Qw9LZYtbVzt+oA+LkOO0C/xYTyO837
pE5BLPdlejUtNf9NtN8jlKfdpFIsJhHygU2qa4ThvDJhJdfG0VKgz1KTicQvcLrXPPKVncn4Tn6w
RkxLwADfJwn8MeAfTGDszh774tSHU1fRgq/PNUC+EfzRPwaGTAKdy8CLH035tnlj/MYKydtLrge9
pXW4wRa8VZddqmtfoODodch4R8GqG6hzUMYNY2Z9g2jtFZjd8q3yH9OC89maMhpixDyAvuxUYeNk
OKLwbXmM/h7cp5BjEw63wyNoXT2wajwjcwOE9AvwwazDo0Fnm2kcnEbwdR0JcVj+WK0Ms1wDU38Q
lBPGvSiyysRZGxmpTnT5oTqbNOHt5ehkel6ne7Mrs7+f4ga5Kt9OimxcfPx+F6++e2lPZWrzgEkR
wiufZtWMIxkJNkTF4+5YysT2VA27NvTJ3WKUDioT2cS97NAJn2mY6Fkz1DDQrAS8eWFMPm7TnOHq
pH6hGrJ2OVzJKPIW4xZXNsLot6uyNNnx7ODavDl3vcT7Uo1iaREerzruFrmf8alFaPUE3iVMBiu/
kSKh5VOATB8Qq0Tx7vl9XAuX1y9dmOmP0eXxURFYJN7+Saidz9vNq0n0w95pJim2+Yn+X2F3ULIj
eHKenKT5bIqUwZJv28EVJlbnBwQo1+ozZ10Z8S8quA08j2n6FBnkxq5UhRIJLALv6j5sxrj9HlCY
rit0De031EBVowSlyGeoRXuJ+5m/b3oThyX0r2Z12PWI00EP8hn+p/5KsyNrUdN0Fpx96Ch8ZTFE
rfw0LW71c8x/sfQA4Ae4UVDWPngOmisuw9WNt5YFXi80P1ePHX9F6mzWfREnfYRziY8GnmJm5nRJ
2JtrIcOMtF18SrypKqVIHPoMFCbhWPYHB4dEiYILK9daDNvS3JzTFi5RbzrxxflLoKcrEKrpdzor
YHaeXO/Ey4bWiSvdTpDNfddPliDh5ZAYokqT96yNZ7QfLyl8Ei0zVNdiSL3TFK1SWBfNL+5dM2jn
rTnriYrEmkt9+e5t+1uWWBQXCo5mMr0PIH3OWg/kUje1XPfOmN0Z49WWlV+IrRSBbUdvrWjAkHJ6
KozCixN+Vu9o9dwGHXfUPdCeUGcXBnDKiMwNfKFUsQT799QG0PXwaaOq7KNlY7QT3B+QdTTpbjL7
Pvx5LdfVz3FLzSJ/wI5bPf94aqNAh05tn7r+I461tmhoIt609+CNsBSIsmBj7AjzjYCKBsXjCqs8
6GGMcoFj+OTMEUurX1oF69dvgEHqHgbtSXQp+LfK8MingGkY/jREyw5jj2qzi2gwiRdWrXW8gsLi
7QpH6b/OPas9U8sCJ9lWOyUB0fy0j6w7I8omXIsKA3lEhZY2/CaLCFrbQ6AnF1Ay85rDjJTxj9Ku
76ox19SwMft9cP4+q7F0BtBUy2X0Ckg4S8nuVHgYR+2PhuA+YN4xLgV4QAvuHCh4hLwV+8ZcTVH1
uyxd0FTCFW3+o9Fgi6HPQvzbbbPy9JcWJzTbNMgf7de7YuGCTGxh+b9qhJifqvy+Fsq6aTC7a5g5
WKHPAi1Fi1tup7NmXft19pOn0yy4Gr7m2iEcl7Al6D+e6nmgu/dGFf8K2dpIw7sxAbQTH5uwpV4W
NXpo73gDd21+Cn0So1o0HsRuoAyLDl4PU/8Zn763JRsb1g6WxetU54SsvKkZeqtexzUHHUd8PnDt
0f2JVuQ/qrZ/WPm5mNJHzJg6xPmZcq/TyUwaqMV09Vema0kqeCSyXnQhqodmlJz/En/XqsObDJcV
9UK4rINUwekj7Ees2DJTtjV1CIp8yxdC+HLb42ikRXUPhQ55VXBfuoG3EkWoAwX6qdDDK+j7yfRP
oancdqg96h5Fz81FNDaDTdialLBFOZYjx41UDFR3kcYNZukwE02ncDGoDZbQqyjuV7zAM9E1195+
X51063yMFJQdgoKQgyeKLP6vpVyGWmMjywEKLM0wBRNJ3k6wLwlywPjdr6KVWBIT01+uNyKNPhj3
EJUUPDOdfW4RItlPaMy/N39/7yRfOUOh2JWp4LA3NR/3ZSTpt5Wr7Yr4t+Ue1lOUN7keuioTNKUA
ZYyjtLqTxq/lFMUbxeMFoR//eHmI2K8MsQcA8CrWAxMAwFyVJmAzCiLEGl9MRIrRzP/U0/ZjrjXF
TyxwixxhJT1P3qxgMOkREsGEd9AkDUT+GSnMdTZ3fr/PipXgxztuz7FfH9BZzh7lrKKuq1fD/nNg
dEKffsyqRsJFqzKzAWRmSskB0IOFtv1Sh2tUYeYx90C7t/yj0FY8Zk748Y/RqB91l82SsIsLynPq
lIecrRZaIv8t/MK9lwN0yv+njhFTGZI3G8xq47QNwPtdKRVbyao9GhZCeX225wPVwnb19uQsEzno
/HqA0qgQtyQwpLGP9+eAg5wa9RkD2v52w9AwmttJOODX7qFX61FuAuI8tXZuFuyzK4rOJrtaTr6l
qk2Z7mnV/LnvQ+aRwPIV8rLz2CArr8BV9NIyFrfzFBVbIEpp8Wu46zVfAx+V/paFdZjrWUSj1yk/
BBSpGOX7jY5qMioXzsIq2nmuzRou58ptVQPA2cPbvQ8rE7xITlwoWzAAVBEsiBr4RPzEB+2ITieL
wT3bznVRo9RvLqdu/ulgzMpG7Dl/rQgLo//JfdLXqiauHpzG8pXyiseMqNrztK5wDaLCnpvi8HwU
7p35afqOZC0fTcoNJQ1LVTxBVY94iy0OqqJ7T3eptFirAa00BQjEnZyO0tqR3J/wcEoOYuZ4b/Md
PBxADNDHFL/1Gn/zUUjBEjfBTnxjRu2SpHWRAM5C18e/o2yT1/oIgdjiPfr9BKZRFPQy7C7kJL4d
QfNTvScNztCsxwnJKa9pqCz1s/5B13PqiE3BYdpW762WXBMA88p6cIrey8fzP7GXoJdHOloiLG16
M+RX8vJSDoXgM8F6ntDPrOveQkLJO2/zkvfm2ZYJPEvvm9LXktwA0vpbGurNZYHQLDYHeMPV2sll
UZLPKc50qsZIYTUuJVYdi6STm4lRyXb33jihoTC7vT0A8xc8bHUKAb6jd/uf5l2Mol4VX1FQ6AG9
PA6KtauHhaJbvQRu6n60sKT1HKmwSwge0Qs7d+ghsEPKzYPjf/f7g4ups2n8oowHTrbeJRbCSPMK
ct/JGm5pouVUGawZjvu2czqTiQZ9hQXCM/Mk8wYfxwOu9gmtklHTuVsCUlrs4tCgCwDBl03na6gK
+KqrfBHMQycoGr8xeZ+4UyVz0r4E5nnxpv0idnVxaUjwUPzRNtNEQ9cGoDdkml/id+T4KfVF/jBe
RXQK0wJSRQDKaAelUqZiQJBB5xb9K2UyJ/N9hAFKgrNOCZfEWLclLS6v9cn4lqLj+rWsCJ2pZWH/
NI6YQWiZMwRdT0FetWE8ZDuiMdl/9lYYIQ6reIOQH8yJeCi9AMs2KR1QmPPkXPmtlj+5F2CIE9Uv
vaMus369+FYYJskRyZsH9Yt4sTNUMGTnduObFfjvtl2zC9hgMRBYGijJIDHLWobjPtQfFmZnT+tg
Z3ya9nsWwnLfMPi1WaMaD6FC8P+9cDlG9uglDooYW5J+YWNpizrUKLqz1QS+Ckz3D9MHcmJx9b5Y
fXezyb81mPzV74OXzb2JKLjYBDuzHjx846fC8TPLlqAnwXiKXWiOPmLDqcN65Cn7XjcuktYuE7kd
wvnbrFwgAG59BWu8xE5uDwSIhrjKMOyjeUaDZXQSCEVWwovfNSEC19UNECVu8aDh9tgkWqIiibKH
L/mhbgxYjNyJK67mC2HZTGHW3AWNyKHDEVt8B8QLfsAAyppJGPmveVDcBrq7XZIcahjIwUU/lycd
WH2EvpFEVhXQqyQkQ08Lx5F3WqOG9EPMy/zja8GO5+exbKlJqE/rAmEIrMi9Uxo38bf0S1xcFoWE
Hegfu+ZanZQ+H3O+5qwxyILOU6NRfa0wAFhhhflS6tQFhN6guTE6EW8/r1SEW6nZfWfNaW2CoIF1
u4GuGn2sHPPX6HfUgtyBpsjNbNblCOTwQwOST8UtqU4sA/l/UtGTe1ymmyaFnu22cYlxqKyTIor2
PWfX30WB277Tiouk1+bFzyKhtasqJ74HEpDINg/5dkm5TPqn9OxXorUosGV7rUN7lbFdpMFZjrgy
Pz3g2EslzD1rhn9EshgNVMRHN+eJIuanXBsZQPo1qNLtr/PVV6JqFS36BlEZEsYtgjvURbI+Oipq
zaAmD/QelJ6JaPv6Y1YWy8bxntIFJSxV/sD9BiOREaUnfI8qm6PbVwp0SHZ713OQyXJmSmkdgdea
BsdBBQ8Fg/Vy9l+zzTtu4fjmnI3U7zjvbog4lItLhk2kYDc98BhJv7v/lwlJtUHzYi0t+iZwMN+M
jUccX4hNOArVaUjtOprvW4pC/P290l7TzNgJ1yYFOVHmEn3rxUueykXHcQw9piYZ/z63reArEAVH
G7TsG3LusX9ny2Q+Lh5b584O9MlrQmkO6bjZyfphZoRpOay7RiFOv0NBsTJF6lhXMJnqG1j710QE
HSuDp4DJYBQ97I6fV4JREHiVVGfx/UJdBJknybS37JKPBLVv35WWt7kK81MSq3DWytWj0PByEI2a
uktJikOREjUQesyvn6GjdthToWRSgNcLUV/pSLAyAIKWxARcfhFy8sC7vJk+LTAqGwGu1hWc5+7s
QG6ODwDuvQ5XIp6vRZsesYW6ERbEoNcC0NIrWi98HH0b6nCsxjtCzWG8rVXa1dY6WyTeXxCa7FHC
nnhRqTuPhJj6prVId/lyn9wJPyGcxNyjVBn8qxnrTOyzPX9GS0d+QO74RzA4OhtnAaZrIgcesTfh
WEWTZV7h/NEnyDpGahtOBjw8XJrnyW5BFJ7ONPkFaizgMQGTy29f35IAo5ZvhO0j/F/qQAGVlNgE
hc8q4ZlYrvZsSr6L3+34D6hMIJoUgfPtxOYvR0keBUKwQJfnM0Jx1+uF+3pgwp3x/Ue8qqU9kDJN
Ukeg7v/FAbowX8is2YFBxebbfywd/GzjksvqbP/8cCc1xj4Ky9WhZjJzdZQ4hUVRiYrAIYDF6STo
/gqe26y4u4Pvl8wsQkckZkAoWgAncEazb5sMrD+X/I1YZ4M9o1d0YIiHOfAYpZigcLIpDN1e2wf1
C6KGjYHbmLAbTR9RTq8IScQIoDa7VFmJ0yN9N//hEUFQe6er0GsiB3v5ZrRoOoZUwNKaKgbh0XF/
riILkZh7fjE+1yGD94HE4DozPz6Nuq0W6gKdeNV1aiXtar0E/gw8zs5vQ1avCgj1sargzNlghRI4
2uqVC06PwFaV8rAcu7jifw0NJlp2vhS9GjgZrSN0UGJW/127FtxjcG7VYF0pggX0I2G/uvotGi4e
2PzfNiMJvoqI7JgpLy6mbGTNjog2xvX2q7bgMZY2PpxyONFbv3hiheWO7qPsIOaFwDEuzXDRLzdT
nAyGpnMyhaynvJSACD3Yye5KKfejY1dAA4z+S18k5nzMp82BTJ9UbvOWMrzR8G5UppsEEpelHhVF
pQSvZMgGy4bNdBrBecZw8/N4f3T/XojRLjNjSFVFR8yoL46C8aCYcZPr754954odoGhMDVsCgGuV
mTl8U9Qmy0btYU6hPHH3VerC/rF5HlJT1+XRdKa48rclkh8PjDZ/QviPmQ7GcX0mp03k2PeD61Ry
EC2huQRkydlRy1Im5mgy3wEGiTHoGXAjyWM/m9Qa15bpq+uce6mOgOPX+2ib37irhSzGsw4PQGpl
SHwakec4T+CbzINEv9XlNyFx0pJoit+PjzCDB7SU+/itX8ZWBShta6mFuK9MQExNVuZH5866DT1z
A4HOH13EgQCZgI0Qwfrmy1S/L2mVUCMk72OXFiso5Jw4+G8kTuoniWy0o/UoAEkKxYXYGhxbBcab
ZSccKNsdeZaQJc7oeFkc+lGPEZo/akV2NS9pcI2fII1VyRrwkY7RThB0u3EzQCBFPFShfhBuyoSg
ngNnxon5oP3RdsKf+dLqjja63JwctI4HIbnXA9LOmt+nPYWVJ5z3dZGSaIz9wVGNDVR/eijCpi37
A63XId6+mZ6xTc/d7dCIdYCYYp/iOTtZ84+EujSfuknbEnMVHR1aT5mEP0hrXeY/MW9OyAusURg9
pzKpHRwo4X8zvM8ifsPi/u/tAFjaACe0COJ0gA/usGrz0VhoX7IxjlcT5OqV2uWGSC8j6UbJapNm
PYJV/Ggy9GZOm/lKuIcX5Ex+muWao1IvQTveeKQ8uEmV9mB2anwigOINNJqv4y8w69TZr2Cq63Cb
Z8bJ6WkEIl1mAtIFVQXudiGgbpabY2ZWWS0leLGs/f4CDlJqXUlEjiXB3jBIkruAkgx1Iecmaps9
0etZIvhFoZjpsL1X3PM1arVva8zwQrvhCSbrMJW4AXA/76ekV+eda9VA4wwnJ38x8s2ETCCgrhxn
cJQIqOF9nF+DMRgJ+i4aSoSdnrmU6MjGDaZ0IqT6EbMC3CbpoxTp88CS9FEbOlDV4lJw1JUJme2V
S9vKCLnIlK2tiQg5wKaZ81j4BQJ28PXzpDx7+3qfeLuBlSHfn8Pg8TQGz8OgYuLTYMlNetCKWDpo
OJ4Q58v7VSfmLEKz+RwH7BXQvR9ELDEcOkazJx0Ji6Zlxytpl/UWBF6X2SD4yNp6lVwXC9vYkdLO
NAPMVbjM+vnSayC1b52LPC1oK2t3llexoBmnxhUQfpI2vLqgiEpiq2Sx+gq0gorYTSLamy99l34q
p59JGoSofRCPETtPUJuy9ScUvUkDApX0kQ/6RmUeaJrPJA2KAfI7nBgzQh/4XLnvSpGMHnFOnp8W
tnWXnE9gLC5E8SGVpz6qc8L1mFkykiKWDp3dCTbYGUXCaPduJQReS4Zi9oy7kq5ERwnzbaPdzzWw
mefykTYS7ehFGr7BHEfiSC74rhjM69Rj7kSrpidrLJwaNNMZqyYiZlQSPDgxy36EoWtcqFfei0ij
TVmGgutfOC+BGGQih3p/tXf9yFtqSYXbYUtHKDjUnWBrCZMMTX2WdeDwyqwy3r0B8JTKBH6zn8up
3WFW1EiKeDgGWFDWcytQ9ot5PJ5+bV/dpsESQZIrnAAsr3x19EbPBBSvIWjWIY8SygQOogf1s5mM
wP2MWC3jSJ5fyAwdwqFn0bI60heuPPDnJQFZhaMQJvjMtnDfZasPn81VpiHpjs+K1ZWwjKdyaR+l
6A3W1AcRC8jP04nJzCg5cleSkeb3/B1aFEtqDlGd9LlD7961GVp8GCfziiR1MmLzx7wF+JTM0etF
8FEK9/nK93wqWSv/6zpECEK3ktO4za2Ld5xYhfUUC4bB4KAvAHxwIDxvr5zJvNaV9eIuxQ5b7IJN
gpwcgnuJ38eGiWb+nwfeubwYs/Y7cRkDDajBOeYzcBnCpIuNjxiZVbsVeouNz3/ySkZbLYe1ALPa
gZo0r2M8rf1Mr1r8wiP521FGxtyf08Qf+286r9tOdsKo2MFArFECo/fEtB2eeje5uPzVuzCp1q6A
7+COAK1ya+n0kbvc3HVmvjotIO+AlipNrIQGvIacdAsV66d/28NEmvusqxAy+j2qaS0WT7O8b6S3
XXP60e/sls6Ks0JdrXKmS0lHyptmi8PtE9bXglvLyHt5LMNJLy+nwX5H8LEdTP7GYV+bD4ulcXm1
5kXkCgHc/+cHKlXPGXfXDFvriywqscolWdogHsuSnOVh/xZncU8v/ZsVchW2g/JdZYTVCaQjiNZx
MSrRzciEFlgvV4bfgO4S7FvMwPI4qohzI8Xf5I7iMBpHmkbGEQoUCDm8AqHX/xqUNKmE/I2LYr+X
7/Ee6bWNWgejJTAxcnXY9a4ss5lYGHAzgS1U6k4GghJ0BBm6DTM9F9OflELZ8/a3bSEFCjGkxQlV
luRBgwemvE7qFocMdxcXsplw2uxeH0V1GCBXdstCDVy80D/5R/FLonI7b+XolSLuC3KyFzQRXDsf
/05o9kLVybZZd0btgoOELDVe56Syjx3LbTPOFOhiFpo9eKjVsnIqFdjMWM/Rr/9H4jk7PHuRudMw
X7KQU8QQxcH8K+BPba26BixLKFfPxgXj+j//CwD3GMT5BmTyYoasJ2Qs8V5653LexCgKyFPrmYqW
Oo+JEzAwhFtwBr0dz0GVs23VsXA9XP3ggKKBN6azMmUZE7AKgPT0LM6ttOsIFcZOkCgC13CxuV1F
MZlYHcRrxBuhREfToNeneAJBddG6a/CmfnbJ3xmwQBe/dgJABZtaRpMTsc4eu6msZqPVmI4+BeuH
U0JP+tzmGiLV4TbLxhTAlAokUsBW6oNzY0A+XPXXY90GKWs8k/lnQ7zQ1Ia1yDFbQE+CWZX677x+
PvS7ghwiGlzgOoAaO+Z0KfUPKcS9K6XJ3dBnFKRRELaVprWN4wtYbyqxCOdnr0AqLvjgOc1E8hPK
MnKJQ2/Qw1xNsDI2OomhyPySD6HNbP76feh4RekM7kKDnniLmd4sYPGlkvoUfOJctaRHZJ2/o9DN
cGxjUUBV1wXtjB72HiT1pgqowUKAjtq0LpCkYteeJgBwEAXQnM8ex1wX+Ud9JRHoasj9NBjwfJBn
ARPqBogceE28tJpCLNYV0vcQI2u7alDjX/RxItYVH7WoBhb09nFrLZKMEYCWLeXfCp/6718PVLhi
1tWVOtp/iI8xtK5JXHxW7l23xb4FMyz57cwS2N+89aCSo6dZw8Rr8vElhWDqKYIZIH1dz3MEqOZg
imFqKITsY854oF+umEtZg4D9lObuH9OqnuYWV/ZU0GVLTs/oa9BGC7tkXEJciRphJPJbOP4/3sYT
Lm++vmbVNj7ULCmJ9TCQnS/U1AXZEC5qEBhqfnbXN/gvHge17F+ji36Vk/pGXpgPpp/Dp2W2wS4K
mxC7sKMGhYJyXxK/2/G+V0Ip2acuHHnLrM0aX1B+/oC9nTk9TdJaDzCsu/eaPe1YYNc5U/drOLIN
sw6umYl3YRTGADAfSZuw9Dw6PSCBGau75u69hy9yiiab1Ul+FCTzoeJm+0dbcspWPx+VEtEPN7Jw
mYTsQ8RUaDdGvHAYB2Ksaf40JLlBt8iei5hBVQ9VjBY6MdFCkwj09MP9OtpilTyU9tlXg/jW3hfU
kB8Qclx/z9NRvb3OX+21bYqg//3DkIn+vzVem6Llw/Qd7+7DxSY2oenI7+EFxSXbU6VO+3eNAsw6
Da2HFOsxdjx2LeBxWrd4RCfFVX7IhLADcnYoStBtBWBSMIGzcyOY5nNl32s5psn3TPqMEk/S/Rkw
Lg7nPDEXOnK6Ad1Apr90rMZk2ybKWfvoaRZwpfCJjSVcePZNluHYYRk4zLA4DLdk8BV4ebxjDNNU
ir35rmHHcLcZoTgyVWNzBdrOZWA9AJ0FpbYLY71KyTZGc3oB/S+3yVTFx506kTfiKiVHsktyviox
kASzTJM3ZqDtMPElglPu3aGsmce6ZWFE4QBRc5zvf8geVkZg5ndn2URWKTwD/4uxU+zLBSa4suT4
tnPXFSedvshAO2vWqwFVawk4FJDBHwJ+tmu203iVOMhH+S9IO4qnyuZWwxGLp30RB+AbRqlRo1lc
0cwCOtZQ8BIVruU1dMmyJrpO27osa0WUhQfMB/0pZPXxD43k4eNTDrc5TGtsW0A6+orWLa7ZTWU4
VJkSxjHrdHPuECsS2ArSogQHzMqQEMrvfd6SNNmyXvrmTkxhJ0IOjc0usNgNHULe+jQF7wKwMQAe
EHJ7Hz0w+89mmpKAKfn43QPPQXfqhrKupXVLGQHhjun/ojG3NwHkdZOo69nxRWnvY6KoQjq5lUk4
a//yNO5eZLf1jdGSiNlylZRO0tk8EurXzxVqmuVoPZ+Ew1gBbEWAorSasMvy9ZmTNHdp5bS3FuWb
IQfcTZbQQCMCNN8zFTrYNx2l6oMHk+VBOAJDqEpChZPXNB0SqWjjcO0O2g5ey1bFZ7KxeZSw9K3j
S8S+Dz3AKp17U7v2b4dtgF24ZtthhmzVm22LwD6rhfKgBOA0mHFaFwMhI3VFglkUZWtUBvy8pmOv
sxVZo5//u/UsiXTTFMgMXCJUS1G6mwmrKRuHM9RqWyLY+PEgKGC1jZGpgrXkgdHA2wXaMKALDauu
rnasDwdsjTKbsGLDl2s0cegnZatKcCdZf9UYqj2PQ2oCkXb9DMBzBPsrdBQCeRSVx6974HequFHq
9KHyRTAl/HV2Ej13ftswpXfFUvAecO8BO7r/DZCViTFQFhjzGJQI0konz3sLpuCHwKCoGLChe0GN
0LaWsNhuzMMXvf31ANHmA/bbbTis9vJ3uXaEQMNBms4QnUyHQzb5xhmnTry+20n0b/vXbElz2bNB
m6x3JWpO1GkMIVmwI+mPXHlcH9xb1GM454VlecnHz/MvVqLwThKKtx8X3exi5pkONn18//HWG8u5
JQmreyxUqOZx75gZcvj/adwRCI4lMt1reqFysFO/91xDPjgy3w8gnI/lgPSVN0XEFJVIkR4G8kXZ
dF3R37H2NwQcZ3M7KuchRbl+qAdw4pweCCTqBSyt50Ke6BdshPuX16ZeCMIoB6n9+lPBIxxePGZc
PezsUMfumQX66kElvVUXx3GM9hvEiO2oYg3LX0SsWWecgooaN5iXm4mvROMruTn4mnj/Y7Y2dvfD
RDT081UZmFo8HUuiQmaXqI29sV2aCNNu0B6K78e/Mn6GBUDx4MpIQI4os5sdkT7efiXkUuULMV53
PO+o/YBoWoSm5h51duNj/Ef77iOP3ieepwoxv8BBpTGYZ49/3pRUvnlmtacukSeKMldhFIKU2nYP
piq6zTDTXkvRGaKOhakkKdtKSQnPVt8Iuk0KLYTfbppOf8zMEYLLcue5hckghqbj6m779XGZPb/o
uUJQMtUWrkPL2C2OL1VddUVgX7rQEOpfsBXJ1wCFfiKHtOCxBvJEp4BQOou+1EZyDd+m1gLelipf
ju1XYnEAI8FYy20Mb+KIpwqGLjF8B89cSJS7/HKH7cetgHH74rl4LOT05gJxW0Bn50a2V7pG2qVG
AJBqhxUQMQXUw14efNACac6YnZWrN0V52Jly/wl/9F/7EpO9QcmarWvAfA1ymRRM4BF+GIg80diG
7Pp2ELHn7eqLKHS6dqB8utwWzNutBtQhNTv/HB98uQ2ju83FqqHEwg2k01yI60XVW70035t5bQIw
SB9gnZo2Rtk/xpAJQ40jlbsztyLi6XN+Fa88uD6rz0wxKEHwotWxykFPL6qBp0VQexmzY0V7nVUC
snZdihzvzq6UW2jb11/szh7HJLgt5p9Yx89UjxqXYMcTBQ7moFx+bIcNMt4yQo1iWx2RoWA9hpwo
XEf+ub0XVwoG5er1wR7mp6I44K/1parVf0vH5RA7sbWoRHL9nYiFSmMAT6p6h9UkO1rmJkDh1SKW
d3kSBxeN0jRmKnZGHA1srztqsKc/bkFc2Pc0v3JmPdVq2c26/kqxz+6ug3pO3KQtJaqnOvPnfhPE
BH3fNr8Nwy8DcBI43A+wEhjwydB1uk2jLiwpHOP6qux84J3GdQhUMuUZhHZfccembrxDPl3AJeX5
ygDA6m+JtO79d3S9dwJklp1XhTuyLErEsieFT6LfgA3dQGm/VLvAbQQ7YghgcqpIpagxdFs4za+6
05o1xnq4g7OduLwB2qxu2ul4Qjn+WWAYux9K0Ay4rPYN6IPFYRaDluCBXyBDw4VNdgKgoYOvHaS/
P8IxsEG0T94zmj8y34Qwxk7M37PdJGd3aN6kROpKHo4YcXVZOdnEAECW7BcEIu/Rn24W+uamGEay
WnH1c0cTMnFZ65QP9dZzaC/woPyv2G1Sx0+S/7SUAntVZ6V2Tl56MkvUFWXIScfOmhL0sgiL6hLm
grgz5HHSU/2HEps1e0USNWVkgSjqCHcfZSTCwkgU1D0nbjGhzE6YXQbLadeoMcmEbXN1faQnZL6i
9U3NPN3uk9eZVhCSRuXJ0miVpv7SHaz3pMMPxOBZ5B+jEIzr79IQNPWFDVnkams2ATISAiOmmx8D
BdSHWjdfivJoQxYbUoJOoo+nnI8H8m1kdBfbFjQXgCvI9u/nGlNa9sqpjMbaC0d/cM3DASzSEjWP
21CDJ/SFNEtwAkuDdozVu7Uzpg865mgrX7cztQqXb1kQNCj1bwa2dvczBeHzI2UUTmYQ3+cJz+qj
1atX/AH5NfXCKRokT5G5IMAVhvgpZOMQp3uZrcepDH7hScP2Ppd6JLPBJgmWathsfMiY5jZcjxC+
40WR5nETOdIZr4AAWE3D6elwZgUVFIdXGWt8owQ2EX1mQ1p/EFxExqsfh+1uoLUcFrWaqJwuGqYx
g9dYDNgdkcjgs7v3M6cOyzg3zlOeTYlSp4EFFOPIQca2e4AuazCF3peLUTPalU3Vv46zpukl0vKz
9jUvkEEGqZgJYMTIjRH19V2hyKn+ValnIaaF5ZtPWDVH3YwNH2GjPVSlzchki/2QLgXyKOSkLUWp
ccD7jUKrCLTS4tZPcrt2a0/FpzRNjx6jBv6KEQBgvMPWX6takF3JwVRpGz7799lucfshur6DXoZ7
kOVhblrECP4o0hY4VOrFbY6kXLsXaI7RtnVL6+Z1Z//F/DPIoEhhOw3rfnqkg0x11gkR4y1HCiCH
bViSmVqi3y7sCt/q+1YPDhFHtbpAQeo5wkHTobJUE6WHHNdc5SDz19mtrQY8VqGFXkwp7ObL/NbD
zuXMQV9rihsm/Gq7bCBjP3zDgX/Cg6Cme/CEBwp19qMZYiKerlEnR96s+U4O/6yykf57w8g4aLFd
Zzss8r8cHEr0Ojn5oNVB0MIqoFBlevPY/DARC8V2XxY+dfbKYTyBlydlYFE97zLETxnbvqf1NHtc
hRyUH0XFkira8vHbR3gpU1bzXgPFedNVZ+MVPBHb0zNXj4cpAxC2gQG0xuvblwjpU9muHLD17/qV
DF883Nng3L9XW9dejEPJbICFHcpP9tF3ilrNjTHp2JkxWKhQWuOpT8LWUNb6zL3sQ8iszdMr2jd9
jW20mBgUlVcEBXpV0acYWwAfXG0PzlrYr0JLSbej7ruub2eOlXF2EAjy+xZSpuLumkAPQVX3ri2Z
P3Mya/kpE+pe0olUP9iGdnJZnQprB8gbRY7whPFKczr4dA00Oc3e+5QtZOidMm2Glmqa/6V8Zni8
BtacZA+WnGAYqJA2e0uKbh7TTZdL4OrxqW8fC8BIMitWfU/QukIaw2mhPf4A/Jzpi7B7zsApVMsX
zpWJBoiRBKKIkb0PN80cbe95bH2+PHTvRemg26VsWZcGrY3DnfeSLOA5YSiWDkriHRo6Y2LoSewy
3VjIsxO3PtKg8QBLB/lpg5KimqPVUnr1vWXc7JiWacO5JdjPkdYlixJW2oNVrSf9+LpO5SaGo2fi
/ajtGr/7CCtduXnI6dVCRksseoHQXIJqcauhqdrmKwHjHD4ZG0sXRIvPzpx0u3w/oz/xj5PfrhMb
hC1lJMGdXecju/+/w97hGDSH/avnsEIbiUSqsDTgyLgB9WLVa85HHFo1hwV2LkAP2ffBgCXHr+RG
fDD+X99sLmHIJJ/ptZbrHygRTse2ldCst+mWD2/sGkZt3coz13MCo4g9pdg+qa420HWAm7TUGz5C
RWm/aBk4+uF/S5esGLU64IUKjH38YMQdR41bbJOKbBW2jOsa31Dw9pA2OYYbV1vszpkzjxefKQZP
vfCLv63YJWJmKvaEbZFckNQjqB3EUcnXF3jW/wKGpzW8bY34jnVXjpuQ4lvKhCYUhbUmd+yh3KaI
1aJESEG9a7QcEtl/GzrdNzmJqocKGw2piBG6JXphjGfAe+6AEXdju9OdrfQ/LKINzb5J3zCFmum5
vZIPTm0G49bnm8sVV76YM8HK+Cbt1b2r78wh3+416ygPUnnVHb+YAYmZpAwlIvbJ9rXeY/NgdFA1
6zSRGy9voe5kOGJshUCGgZx1IfcDe3VrzXzm38QdVs/OZ/jW9HGQ3vNlxzU2XRlon230/v6x3yM5
4w6qohErUdI15HCqZ5jZ2WHrO3tt2rccQtEWcMOpICKMSfa1G/sYww0Docbn9p1qSK/sv1Ra+WVN
iFYEsyxbUSEWuX1lpF0C0XIhSikBzO40TKq7dlZTMPhXPbEG7w6XDy6HX6Q/YWfgplgHc2WsEUSM
s8sS22I2sftFK7vpZM1yjfEiNPPrrikmsS1gs7UvrwUd9Uf7I/OLXAbmEudSpCDjwyLASFbrzyR1
PZNXbn4x8EXYlLJeAXot9+d1PqVnk22S0MTTX4kVKLf17wwZZLzVaPx6mrO8hsVDrqvtT+tI5lfi
TeCwwxPZuwYLZvQtgUvNss4aFmX+IMbc9cDDelZEg7OCalU5J1b8780CLmqp7u5ljtOIdGpKBet6
+XDEfBk0ND67vnZZn0v38vRI/68sAUaH7+1YKCxQEN1F6SsanFVpQq5CVfjf8UyYX94gaSbDlpYy
DGgqM7gUFKTkFSeC0Z4wz6/lZI41zxP8hnuKCzZt9nqaAqcLhLO3SHbwZbo84Izuc6TjqZTI+r2+
xnXxEN63XXx6lLPy4pAfmopLVxqYUuGuYnlHBaepXRbQBP2MIoTYGdKr5PBb5KmnTQ00T7GmQVDz
B5Gw4+Tn/Ht3h/gd4NYMNSO1k408JMwvb40trnqfQAa1o1cuh6vdu7GJsU/cRhRfsajD3hsJLOj2
72GIKCIj9xrsHuuZ1WerZJ/RjZ+J9II9OHHignWALA3PM9rVxf+NdtS8cyDOBrhhNlgv5TKJ7tx0
neN3y5WnfnsT4DEqdanTZqzXRAEdPCtSsQ3SB+B2NwBzYiz1adkR8mild0nR3FsEIoSe4rf7LwXk
wa/iaHYDm3fX4Lasl+1iH4yTV0ptNYoEyAoDJuJWvbOuEGMusEdSsaioCcWucWy3jrjpI0ZYVASx
BnrTskz7oZTc5Usx2bcAPv1NXkZn0gWMI2rIvVZd26JuTcVOU4mq7RjYQDSVLmLq1cqxN7I+AtVW
y/Pd7I+B22GoQrs6j9cQuPVTIJ1qJfiK/zOa5OYARo1u4XWHo/FWE+A63+4Ylf9e61sLSXEkuEOD
b7quoiMVuYd8/Px+3a0/OzUNuqzsrmILYeX/4zy3mge1y3gDODr7SUlxOPmlekfcpO1aVLTrXNw7
oq7SvFTsR6R0X13JBDwmBdBKI1s4EAcpcGi7zECzODSk9qtPcW/E6UZ6DXSHu1n9tGsQjmYDZJBP
OItpv0igYYN8r6BXfwOPTagPHJJkXrz+i12eoOcwtCbIBH4jugRkFVYJ909FxquPiVmZdL/PisbY
54DttG1yXNxSzNdm/l8fszbXJ+yCvgt0OrnvE8y9xk6t6HVHjGDOo5Bd8aW/0VGXcoeuvU0Tf2FV
+KLPP7S4IwsDhM3F5cFDMk2hVhDPaR2640dxCnY0rkL5J6KLa2CgFGgdVGMh+AbHBsN+xW/hTYC2
Zfry9dndVKIoejGkXNXS3L9oMoBz6w/ybAZAhYSmcqw4GNltEFk7GomK+gRVNE9x01U3zQF1z6O2
vik3L8KnEOspWtoP7b2XxGp1KJeE8QdW8obSNfWHdXyIT1B0V849EaFAmnwWaAU2ejKSlcGl9+rw
jY5kxbpdA0ttAdck7iUjzo0RtxH8NS5yHBGDSK79ih/8LXixcD7Hm/q42aBUFxrKifPFDqlTGXCw
OEHEy7L4Ve9SkOkKUonjjuzr79jdivKkskXhWyFlpZn21E25fkCgnsBBEK+RuiHTEjeieqleCmTf
scwad0NgRjr/jVtFPJKtH2sLrPOXcacd5z8MlKwWnhjVCFZcRzShIFeXpKpJKcXx/Ul84cyhkIhu
C3whIwrnQDytSKtGvDTpdEy9a4p+69JwkftUd9zDhGhbZCgp2Yn0jaI8AJHoPQesNwcUhvklkM96
WTd3Ke6FoOdC7tU93Lw5ZtiM84cU/AQG06QDPYQhJnMRgmuafPhA7wsbtxYPjj9Nc/bSnCzvHX3p
nenH8XDRUnEDbSpUq6ANmGLXRt+sjJMrDN5ddav6ZcwpiDOOGCfpCGPf4ST9/z7Fkxk39eUJxQ7s
w5y4qEcuMeJAde8G9Fv61r7xp6EAaElMulCMVicYHeEAbAXeIQbPyuK7XqS39Zzk9EXPCC+4qKtE
+VlMWxdyIJobpCSczUJiq4XRoihgarstGGWOje1Pnptknh6ESGf2iamuepNrB0oXs/wMMVhf7xuP
PUJHzTRHnAD1PjJMAjSzbfILTGFP7KP21QiL8P96+2Orh4SvgpneKQT4+2g5VdvvwKCL8sD9Vgg2
iJQKUacxfmJiwazM8V2rjhDxarhsb3+jcbb7K+jvWZSAFCmq9TOjue8oCqMQ7VE/bIsagunPo453
/Ym3kbQcc5MSNTnWesh08+ZNRKJLn0LU/pGr4H1EznlG4iKMyDcJz6yqhhhfxvwQbiQjqHIVzQjd
NMCd1+IB02l9vXswa5BeMiW4mN1KMxdxCeT0Wzg49apOj1qurgBTfaJ3GmrHcdnm88bwpUkwfkXz
/7MHaR1S6r4hfJ1ux4IlX0mhKMurVccl+Cvm7u34QPxr/Uy7c4SzsbseRxqXvgahUDk1P69c6k7f
EDP/8NummFRfzx6fdTINq/9I7aR35Z9RrpcOLOQ/7Ims3g6rFqxh72CIaABQkzCSnaZ5IZz5j7Xt
9nE4i7hMOaiTl0LlREQVSZPOvcbAorPiBsD1rprm4ji0Mi6jV/UojUXHaGjGL8TTdx+N//iWDKOn
FN4H4isYdVOGc6HfVgXWDYgaaQzqR3hxSnf/2Yurr23xoi1SzQlVkfOHEwCnbkpN3d0oGlhCwhtI
ZUJJnulJpcOZ/uAbo47cxvOmb9HzQP9B3sAJINLXlcCQC7L64xKgsdE46PGVhIFrCxixOz3Qcj/B
Xu4nBqeTXoc5/Bopysgnren+5U66ozWX4s/cWeCylvdvuoyXmIrEhITeJr3Ec453rBOQpNk4e7o7
zue/LBfZblgWD1I7LK1l7iJvgimAJpOfSoJ2zgkF2R3x0m5k1gaQYXHne6s9PnWq4W7+QcMX1pbE
pJawfNPRDl1tYuG5QdJOwh1LNO0d5RKkzH9S1OVDFaZkwrmmE7Is2CRsCAoZ2ZMqwrpPtZYtiwZ9
XkaI64nxseEVgqNpccWVA1KADD5yHH0OYDFvU6zIFf0WBIF1qXBxC2QxbS2veBpw9ES3w7Qjsx/A
YKzSwx6AOb24/eJi41HViG9iYR+Ebqkje1MY8M5Oww/O35Y9gPisWXfxyiIMlQOT8l5kU9LmijYQ
lkaPmTTYmPl6w9LNQN48hU5PW3RzyVHQV0kit/iUIscSbcGc/cnMEgIgmcIVtEpV6cVHfKJ43jX3
k8xLt8KaIp5ZaYqRWZTtMbQw6vrGJdcieZeTGwbPbMo05EKgu5UMX07o4GPSArchwxqb8I0G0xXh
N+W4gtH/YgBDeM64GKmYtmh50wjBSxCyqRrkEjVb9vhm+Vy8sOxxHDzqdyYI58PUAfAoX3nVtFfH
bVRcjqP8vFQqxjmBIi3fIvlv2lPSbkZVYmBOgOP1kfos9Ub05BNIzJh8kOS5tal6QWrfFxWNVSxI
7zlcqfTVqAiMO5qYvxQUP+kBuwgs+TPkr4g+IjuSEkrtaqvWLb+XVfp897h/YVlC8ZewsujhSwHT
PwYGtZa23tziHYPL8JoYTY8KuEdFgHYT5pgITBoyD3NDVVPddJ00IjQIOI/fiUC3CPj6wrab7zWR
24j6r6qf/SgcpGFFZqBt06g+L3vAGh+ij2mkVUm6pQo4ZaztQqa+vaY1kijXKoX4yjlCtQxbmrSx
/sPt0ldH5LaVCYr+ujr+l/FdvfsjL7lX+jVRELz5E++7seZdOYffimxiSFtF1e3RhLQ/vik+4Y7W
QRdP7amEQw3vdLv2sIHjrOZVZNHxbkrYrZa6M1nNzSBFy7cHv44YELxvDeeij/1UK6Tic1dmq4+D
Zg77LwLBDv3pNmm1Y3EMdLPl9XaM8m0ddPWUhzPfwbJtCXXMm4vqR9IK/8uNQ7Tj386y0+kwsUIN
CGJ/daVmVSJNw3xReslcbVgYujtdSXkNue/S5B/0tcBKSnhR0TyQhBWW94woJCnugqNl88k5eoFf
z2iz6sHyvWtTByB0rzyH5QTSMtPA6XagqvwHfowLAU/z8eHK3lSc97sJDpksoDfyUDfu+wSVNYJJ
TQqNU7qf3pJWeo/I/m9o6tdRmemgwqZkLPlk5YFIe7i57VjO5tbq78iKMSLoXVPg0eErT0o+dOLm
8BtiLhegj8Wyy4zVfpaX7E329I5FQIOt4CUYG4apvaiwJhr4FLr9h+R7jsLfk/Uuk7RYKBq9BUXn
gwG+8+u73YhvOlWFQci55+hdJwbcW1JaTYG3pyCPmZjQGkIDfvIG99/jBqEUS8GQEfcYZyHS3xQ9
c7ObeVZ0swjsvlqWTOx/QxGdtiDXy9ctITj8xN4vY/9HVexDWg47LSwOKgaFDOBuxYb0P2CqTZoN
GMyMs7lAqRi68rw0wGQ8qoGqT0v7dRvakfpkb34xoZxG36dKMASdjoZhPreEQ57SXryp895L1bk2
GRJP12+Y6CVeppWXJN1IvQcFb+7WoglZk20xjK8mOiVe0wzkTLy7qayOTeMt4jqAUn/4+I6/zvFO
iuhrzBSjr7MK6COARCPQ0koX4Ks/xpOBgzJgsnYfpUVckYbeniQ3Oja01gv1VwLPD0FJERWOdG0m
5EZZ7tLgHEpJ521qcB7UKILvkMnSDVgHUznruQAbogTtKql49VVn3Tg1Sd4Ut0ymvBU6+3strurv
sVywZA2mtO+DBIBDsGjZAQjtQzs1586ksulb6VY4fp7mI1m81L3bjYpHYbRgdibvmD/paOTfIeij
Pt8ZGw/9OtaqaSyjPv79pZoU4AY+5T/FLYs2LMAEfPtgeypkIVRu7+NNcnnzFaoV6kJkIrdt7WJq
Br9VwYMeVPWYapD7A7s3mxBNHtm3ZDBBM3TV8OxqpRFs7BE4yF45Fmag0w59en1Td3DyYmu1HhLq
CB+3XkWiO5utcCsqtbhteyg/+AyRc3j9TptOlxLfDsDe7wAJ7ZbLpuAmi35T5wY2k+1iqp1S2knY
8ChqcqBGx/cEA1ncv6TzVijsiU0Y1Mo/6z6vxE2eL/AuBdmVcwz4QlpnpSqzKasOFM5t/mJ9R7Y4
zukiPK/3BmY4cNo2lXV98XverJJRZczj6ud5jiMTYvCqojT6ESK2itcscWIrbjuEpnFMFnjibFKQ
3KF7pGdoQj2+gBP02zh3qZ+LUkARdahIhTnmHCieK4bS0CbAtTAiXwMsAAMI/AtnCRO8193qIFC+
3JJmUmH7sd+qM5QlO2eY1GBx0wIf5oH+8HuqaC+D9cNEL/QVFSm/9IlRar7b0dbCMTPPmCebYeG+
xXK4796E2eyM6rFkuI1+T4kauYRpkHKJ3uD0Lg30dU1ZO1iOd4hRCh+N0BphoKGYA7gQLexLIYhz
uY4LLnI0M7Sdqwkq9l7c6mMDR9mBsCSy/AuUWqdcSYUSok7ei8U6VCXQED2HQVXnGFw3lhitIBE1
6f3XlLVpVRKSi2S0/intVlNAgG/ET+6aTkAXmviGFdF0GkJ4m1V94b6cOVGED8OFZlg/JZ0c/N8/
2pflbn5QGHBtgRd7tb8DokbOe9jeEcTK7tHhDc/VziMDG3ERTpWbww39APr5zgbrYVj+B+PliWTG
BpQS0johEaledTGjInTVL+4M233YdiOBj+4nPvcbWatBVDvxLA4FJJSd37vNBwmqXxIISi0PD3Bm
rLMJmJ74j852XULH++lFMiBYBCqqIqX6rHTv7BJjVgz1nAKUsuPXQVlaiOXPUxcC9TGfmpQOrXy0
owJDfja1oCh3rJ56z2oRmHR+ja842j1PicBJ2R2jidPSnOMUSD5LUmRN5F3QBfFXbOfmxjudCP83
KiOk5tYBlAXLPdr9G6LObhFTLdqOspyN87HP0LLvQQscqwZBCeM1zS2M3pLny7Eav5BObtyyPSPD
w8vtfX1Ej2D9/XXkq8t5WtGkEYrOGbre5OtwnndP+vTCzjgneDkpnvmEYh2zzQ19Kl7P3XBZZ6cO
bYg2zUf/VQFXXoHxkEH8gZBKDRd1IAnO7ANRvMUAubW4iAF1t5BKO5UH3xfjacU7RtDX83ynzvp3
vmoVihRGwvOP+MYc6JgRQIUHoOTpp6zkMBGiz5xYmhS0Q4gPitLXm1uLd4n9szsdrFeHvTQZuj0Z
9XQWVLXZiiHmV5yA9gLXMmiqtG7n1F4pIq5aJvfSZS13WQJoNGR1lI2Z2Qvto8+QCp+Z4YY+YnOQ
5n6iA25zjmTfNOk7x7Vd9m11cpgm6WRJJCT9pV/IdmxoT9SKs8Yl/uOqSS+V7OdWA1nScdVz9R4z
2Gn5IhPw91i7GG57JcBOzxRe5BzXm6QC5zrWCrHm3qPMz2RLttXHj4jp28rAuGUxNCnx39qVTvwj
hleHyZ6BmKJ/sr+O3TV+DCc8k+nAZ15EtF2HzO83bzU3bpTlJZSv8NrWtxOTUxUVqLZFznELU3jR
ASJtSmSjrjygdiqrybsnbLUIMp62Xy+YZ4B+k6Mnn9Amg1oEkEVvOJGIXPTuWNH9waUBFgevEfPb
oduM2ye+cj6iFQ4CrXk76S1002bGxt4wg1iiDaSdtDHWOQvcuNf56JHssRJE4w/1OphAQ9QONt5k
saETuzao5MwF+oJA50FO1iQ03lbLkpSxWJJrtbFVyfSFa0JTLSjmfAPERasztq62yo+2o/iVGq6m
RWDtobPXxiubdxqYd14TJlxeDKveg83edV9NEtUzLF24K5a1kRr0gMaDxxhIyJT2Sl8JNN7hTRbZ
SshFaOl5LKWubu+GuXIOEqAwVnU9hoScpGp0eIdwv1cCvEdEbBQkDh4ynW1M4c6Q9z3biItMX2Li
h5jBPotwIc9iRXnIWoSjRRIBfdJ9vZFN1uQpKXw+MK0R+vxsZdTkutna7ziHamw3iMYkfb43jy6c
m9rTCxStjBM/xJjoWalc3AABVg+evbCu8AS4UQulshsDgceU5UGr47gs0xZToRsKpb86UQBy+xXJ
zCp9EJNvmFrIAjC+mknZ3WONDnwiO05fUOHQf3NP+pFxZsrJB8IXrf2SBKhQ0Yq4aD4y8Le7vDa3
or4CdyjsckOsnFj+SjVAk35PINJoKKiKXPbR0kDj8Aeghi6vOfAnhtACDQ8UHzNvJcmfrnkMc2On
kQljoUElnnL20PkFlBfHnwbNzzxhJGNsIZHDYjQaTBcA/AgUmKWWzHPPveqrP/o+F1wt+/boLgLv
jgk26czBQwMthMXseJ15qSMXc2ijlqdE1hDmjEjYLFAqcrS3oMTc7brQ/JIWxX8jqDJ5gxUxCXKt
BM1GZR3llIPWstnMqjpSkQyAv5LqmwtXO7Rxjt1mkTyfdUE7l6LgIwXLE2PP/bRhJbEjxDACdAyT
IUY249dea9mG4x2+tjUUlpmK1v63mKinfLzLtrcU352rV20Zq0S/gpo6opAKvibdbjjhKawYS2TU
DZQgodEH9sX+Di3+y4ND6aGItNCIWDs/hmp0NxTZ/kV3i5gjqm0Tc7Q1i/YbPe1vozXy4j7t4jmm
ExtE1AWyuaSK8lZD0M14ua4beznvPyqb8hawsJQrWbl/b/L+4fyHYC6g30o7n9gaC9eRlCTuyNXK
eZDR+YK08zHYRAqzTmvpwwRTAzUgcb9wwzvCofTGCOUW5ued056CYdDdfbeJdRtlJLdh8DG9KxnI
Lb+BOv7SEnrAXPSU2hHn70vRPRz1oa3fKtsqFOwUSEe1fYCvaOjc+W1Lnzjv6/Yk5xTcfqrwWyYO
cHWR1AFI3l02apJWGq1aIllieotBfRu+x9kjpXCDugAUYJtHUfkMbzYwnactQRFsdj5rF75FaYmq
KBu2Aziwnh58UKmign0GZBcdAZnVXGUipydhcG32Fq7YSG33P5hltmbYyqGU0gnBfTtLzaOm8/UG
jnvnWxMCkJmotf62GXPeFhyBm0vgGnsZ1qtT7gSS/+BKVGPAzUf9E+d+UgDKobf3MaRVbMYWtEli
oTtLuIP7STr4Ba+CJrOdDBLxM+d+hIWf7ud3HQ/6MwUbE7XhS5ec/TX8RRNGSB+LGDzMF/POrseb
OZuLYDzqBmwuXiSH36f/RLiuvzFnQpnCAphTMEzkMFiMnEGctbQz3I9veEjn06YR3JISeTRrriG+
hQqqrL/7m6NAOOxk+DOSskurORbe1ejFzHhj712JzqFOwc0+CJ4REaoc07uVX1Z4TKd1uFM4FqOp
gg1rMtGMecbnwBSQ+1kGkOZkC51p3C4mME7WoRZ6ugQSs8JzGW0uhgHNLkXedGVKIraDwmkDj+t6
5aSwE4tJ7u+u9hwkBCVx49sZqBs08JpUWi7zLjFirCitmmK0hDf7GXdLVuIg+LHvu0AON/WeAvXm
/veKvxxgXw1HY7EDS4gruHaCRO8k5tjuteo3/MuW21XYCPaPBiHHufcCvhpgsYjbzBdDbgGrvzVr
hslVaWc6NFPIQ+6JUdJLMw/tB1/n7IbnQG26Zz9l8NHr+bD8tIg3ght6c3c+c+Oz0qQmrJVwKp8o
sMMTPAqkG2IdWF9HGciyBRSIU+OvYdGR2Cdv/ssx9aQWhm49VN1JgFR2lnf5LVGxZp7NYilqXsSE
/3zAXSSZxP1sQ6keHIZGtW0XrWTQ8toUG2JIpXsRr05J7/NTfnMyb0w52Md8laKz16ouxYCVxgG1
5uvx1k0KPckSMPpMjzLxd3OyFx2epydPpwrcilzmpJMZUv5tvkKpyFZX3CduI7QqYAwoKqa4vSJv
ZcsswW9ZI9Ple7+0b1dglYf8pNwiccKlCQ3dzUuRTedL+QtaNZQNdUortDg081oI+hGuTQ27jFJZ
KhLuWKNSVYOmKorU/zrOmwuRHQRcUp/U6bznEeZ5bWVyq6a/1wEhTCatVXiBpFObzADUi2QWZLMz
mdUxciRovGz5iBS98W2riWRLnyf55ZUzYKWkGiw4jmv6H9fdXZRdEEX8Vl6P233d1X/LEIH2FoPt
QnFDrk17pWWw0hvoRAsAXRffzPMhuaSZvNvFqZ6VlpB1Bl/GQqTCeiBAPk3Hel/WJxxJ1MQy3jak
njfaypgKd5HlAj7dt19+vXkVaDPS4u2s+8AbILUv3G2aWgw7q3X0LqnQJ6TWh0S5IevPYzHaGSMa
aMxAWp7egi4LGbtFYcEMzz4eqdclBZU7D1JQUIBOZXaBYHVe8Ni5ICfs/GnzC2phzfYMcZ9/IwxU
TPC+sFFyKjo9A6PmHtrmQtTkK7aXw2yyDuvChpTUtBtI4FS9CKkXX8QSIzdYOJgqgtrflwpQtgtu
gA2e/yxvo3ms21ttU7WvJLeuuVg9c9L6115L58hhQZeA27Fp7hxMsN87oB/yaHuvKrqG/PtAaz8P
QBsuRbykFqeTfNodGn1BEo/i67uGcGNII7WEvOrfU7bV4dAf2dZS+cfRdCurzVBfBaRANYpmVQz2
1HERwWFw1K4lah0C0J20iafitAC59fTzmsmqtLcV5rGObO/ojgs43kxS+jJ/lwdA0IHTN/GVnm1Y
ciDey53XMHBfhI0Enpt/EYkmqT/aAzHEpAAKaoNXw5ufB2BgiDJN0VdzCl5kxEgT5ztoFv/HHkXQ
fO3CVdCiVrLn894Fnd6uUBi9UO/JKMhIInp6DNjEhiX0Sxrb+CO5DtQubHXSs5mONuZmk6zYozN9
7S1WGwNzzo8bw1VhhksEGp3+bFvw6ETOxkVJiVE9E+Val+GsPY54yv3HWB7qzEcPYwWwwFoCTASb
jGDwU0Q0HolD0IL6pm5ir4NTI/Pm1j3ePuLAJ6QVw4fmdiqvlG3wowudo5tVIyzW0BulaZquDZK6
A0xMH8duLzGg2L78LlFkGssWkcIwaIRzqVmID0EKB4nCK54d7TfPGiGLxYTD6A27AFJhv6jFvdM1
QBMXqCVLRuhFWy3Ns/zmNErbhW6+KQOEA+QhJpaLvXRPCsItwvZc+pK39QzbTBK3zsH71ceiJUIZ
5gh2t3vtB+43+pCneJmUvpgQVXbh58WusdfdQmzIdRiazPEK+BT4QI+bGW2LLQGOu5Z8KAcdO7M/
f6mXgcD3tU2Zw5wwlTm52jw1RkT41Gs8zMjUcAuOFWQNvWuayif8ejALXtD3JQb04b6414NikEMY
lkwThrYvjQhhEK1ZA/Qp1PcgfaAlyvEgTYe4A+9bh42ml7ZkMBOEWS9NnYpWn1w1ndVXrIsFGXhi
4eEwIIG3KrjdXDi3vQ1M8KuZBUTX9c2Myct8FHEVZBBGQHrF0VJClnVsZB9r9WNLndulcpCpuHk3
FCaoXuIbMV8qQ7xY7f9crNI+5c/UN0QHGC1Og0o6u08g3uiuDEVYn/LtHts5ctYDmtzB77m4gw7t
EDjCOYA6EomF1uu9ueDftJXunlIAiF+gY9Oa+MlSSWl5qoYx+7d2W2XOUxS5RZ2vzNRckt5LxVcq
cpnxZOtGxqxCkPawe2Jn6kLPukd4465Xw9+8hI5OZy1FI2gUv9su2Q1D66Zz1cSlGFtoAoI7wxXv
875SW4Vey6pRrreORvDSPNNwZRqrzn0Umd1mIcUJWSS9uUHw5vleKciGQMNjreymUCJqC2YrT9xV
jXfGh3h0dl8v5luqzPHDLlqHhR8ORnXt92GlhPJLVFmGX28rknDc59JvIfiUiSVsNePYmi5x6y6z
0t7FgkD7W3DFM2qVg1VEg0T5PfO3TMJN0/X4vnL03rXFdzRput9PVnDWpRKd+ym5PtWChES6y+Dm
PUaRAkU5fwFBrZ4GUO5dibyty5hnNo53/lTsrGALyG5peCrafiQIrqY2WeecCLzcUk677mhr/Sm4
WKJfGWzzKob9g/Va2gVb3U2kNdY10uQ8YPggJmBnnbFCa44Y1kmpLSwF7CfHUeQXFtHy6fRFqu3K
wXVSNZfIJIAnClss+PLBHcnYlb1UperdwoI6lm1QoxyFbZ4mVgE6AOZ8su73ZXdxkjlsVS4j7G0Y
YPyG4+GmnVQdBRsi2mphNaohXQOWrSSDz4FYfxU9k6uvfs6yx1P25MHhjR26cs4rCF+CtXlTWMb6
obbtrYOBGWGh8FPQYI4oeMEsJ5w7PbnZpe94Hz+QjU4qfiEa8jxvjM6GP6raVAYXEjAQM/Ld9fRQ
G/cfP95rz7cR7/glRUR0+h3fVaZJhyouqsvlirb9l1cKBseqH+lcIv5a2oCjhwDZXV0X81pi8g/F
OXFQzFBzS5hGd2qxPBUq39h9HV5VEugdQAq0fDNa5c1tJyj+ZCWVeRwrWgGc7B7gqXA57UkAzZp1
O1oYAKUSvKQXAVwykecuoepLMsjzKqD5cfdiU/uZACwdad5xZK3KgFtYprtCjjlfEpJutMm116m4
aO5AM1tH3gqoKzBAMtTkhtQNr99NlvEqCtzvJlmKlvFAfuEgCIKt6l5uyOUoot5RvNPG6kKq2vD5
tNn6f4rb5HzbxLNjPSZBhOOi4M2xSp0cwcxC1FZL0Uxsui4Xw0fVrOFqIvLhgUOzHvkduHRX5t7z
Ut2lbtrOl3RJxrNZdQ/eY/n7kuAAr0T7tc0YQ7NPNmroIVi70QN7qf/Er+2d44E2V96xB67KIJGH
Tj9TpMdreLZNHgwSVBnYoHNSDQabwVgcOZljFvdREZ7NzUzd7JKCFoYKDUkKZTCg7tHSlRpzAGJq
8VGIuurPgZMWlYdgdywi0JhrJqJpHn2YO/HBxg4+Kltl60KNSe7jLxMesxo+ITFRcrvoWshlDdOn
JlZDh7Hyuz9T1d7tAnM6rfuUIxpGiHqCuUEcya38TUbkbWIqibdGNZQkEuzndW1WuY2BJs2TF436
bi+Rr561mf/lTkX8salaQWt1HcnP+I1/JsLwpQQXroKD06TouATEEoFNvWFNXYq8yAYA4lUkXt5n
jS8Q1momv6h+6QCkDiAS78r0f3aZ1lmFZlNsliejAOx0asWs7SDLx5bBZqH3/BIB6IpOQ5SJWx0o
XW088JKdmFMxkwNqcQ1iO0DpWWKbtbhs/50oNY5O4WpJSq8WGle2MGCoBcbXQwcoSt5stXinHNrD
iGI5F2W4yOPvW0fO+SSYaG8AVPN0Gbf5tSgQYMtj9DnHolCTuStYME33eCwOtHs5oIA9QExjo4So
f+cybSqzjEpWW3zuFOczyj5Khgxphd3pziFN1U3z94Ax0XN1E9qyAzrSa0A0h82/oyPKiabaf+VN
ONCZH2TKi93JuM39mlERjeRJPC8mj73Rocp6JjM582yys8y+YmQIYqaJfk9T4QM4PBbASJTezvIP
sBZvHLSXXMw8NaOC1EhGvURA1t/HfqgwflPnHJKml1o/JnrpK62vVjgcOcfCTLNX7y0Zf40Vamc3
R0ai8XhZZT6hCn2eskP8AM+ecVo9OJ8wy6OUPo5ZEpufWJWzIy2dfjrmI59gyigLsrGw3b7R8kJx
5Tr49WNyQRQShdPDTxBHyTmYanfRvr72HR/ZTpcaEqD/6PD4HOtBHfQt1Wwofv46SDv7djE9ZRbv
H6L31UnhIE/T/T78n0QuiVxrf2C21+fuz4MaK3togwkU3Ck+ejlnBiA8I+15hfDFa28TGzkgpZf/
g4RyVLZE8M0/o06i48wt2SMCi76RVGmBxdM1qpBpE/IGnu353cebskLPQTmLJjKxny6ZH7RM/SmM
82Q7FZBC90Lfs7OP5Sw0OUOlMdt7zIFfiHosWN6t4qNxARhtcmw9PsYzvaR7hIYg1qnt9iAOSggF
GDWPE5dULBshRRTyeB/c3IKeYrfg6BVRVCajd1u5wB6cWNZ2TJmB91BDMxKfvxxszhVKNFZlLNZr
4T+1TGNnYhBWaq7TA2Pve3T0S3/oJbjZENXmE5ziY893EMvKeMfaXta9W11VmLlvKX4iEY7DUx1E
HfDRKVXdQ9h4yIlYfEKkc/P01qe/EPFvGowAb/cMM5qAdBeVQQgKDxmtvJKrHcO2+hWrvCD5Qxyj
A/aI9e3phidT0zPClrMi/iMiIyPVCGD2PGyUmzg0YnjkgpKMJ7RDztJOdPVGXc3iw/hXLXb4hdZK
5+/UGY+28q36a5bX9+2E2RsyXnAZNgnrUDWdXtM1iBHIx4CfplADOcpOpp+wy8sI2z1TPxiNjHqA
kNY3AkA8PhdSSfw1xaSV8tpChp+pG4i5se+uzj5kAvqd69Voa7TD6S/GP5y7YuO/Air0pNlqElPa
dvtIWrFLdINHbsYLbnHDyeE7pXmz+QFK4PkDkjlGdJlJwNi4doS/F9bWqufl0i0VVx0sQ1M43PHh
HuEQXi+smEMdQleZn6lplK76+o9mN2o0dnqbTBxDFVMa6rJa0oYwLwU9R03nj5hxVt6825icGNei
b4o0s2AboWnmyUjVBrZJwqbfDk0n4Sic/TCBZ/LUI0JlxgmWDGHD/DyvjGGtclVkAWLWEobdsCLk
A0OKQi0/Eca7pmA20bPqRqAStfB1sUv1qjc0fUSYvtsQq9VOm1XVxcWiFC2lQbOj047oEicu8MTq
/8U7lM6OT1zb+JmWg5kEdsZR3nGakJxrV6d1rp8obVxzpn+eUNFej1dFfLAeOOw9HrQ3gEvCsKdz
G29DuIHKVf3bbboNmWxrGMCeoqQDTXHEWYYJ86ohwCEoUPPqrts7BWIaW4IqLBR9XWlchgdPg92h
q3CnacfKRCVeGpOo/2HtWnPG4j4FxGhe/JlRd47asoxo4LIMUmwjoxJcPFCaYruwzvLjM/bR5CNt
LmnSibW0ti2zM9iu+36V6v8WsCWKVzFC8SRoRbEWGhW0a6EHLfUvddXffZUrLyJ82cP8gsxQ+y7g
bGivgV4nIvJw1T/klldAKV7kDxKV55dQ924F8gNR7tLvYRqvRe7TS5ASrvQQyuVMH+PuzyN3/1Bv
6zjGFTny/d3eR8siUw5fsGCCnMJslzNT4sfOKYoWszRC5VXYcGpTTJYa46mxgiLUF9Z9aB12wl1T
dT9zBNZU4TILkXPKFT8PQW1Oax+bgl6tQzneeUjk5Rlemk5Ka+ROnrxM2hIDe8hed+zuxygmZ2oz
C97GH8s3tcwQBEUWV3EKGrY5W19bHLGyUxKdnIbsST00P5u0CZu5Y5JXGg9FS/ymxNR+oMfNqKJ+
TJOaAIb2LYB5Psvv0z1QI/tyZbDgayhCCcDiPhckptyDrueJIaI1gOorYplAKNZ0MSHtxIcV2IYu
2XayzxEAF6CCAT6Hu+cNKCHnmLUgCRWRjJZroifOx3r3EeRjEb9JZYIAZoTqTTL9NI4JkQXpkotJ
fv0QEw4AUr/bRj+lbklVA6oUGx62SHrcAvUGor6nCEX+OsXH6OGx5dMDpoAY7mrahCAbXyrIVlXj
AnQVzBNSBQmuNuON2OeWV1pxo+umS/bb+FKlSc0K3oZhwoRXIJsQ8h0Fq6XPZbcMoBe4PJ00UGpW
7zRh9kd2zE4OeK8ys6z33OPJmv0wP7fLT1GY47EQU9CszLYC9nZIgdodvLkE5nAinT8Oiffnu91Y
gbMbmLcI6CQwIENVsFEx39fJsQllth3CQjQnR6FbPbdhgbnsTdW2R9CT5nCgskjcnqZtzQPdBrTE
NDlGw3cBenMllUhr+pYSmI8S663ftSDs2jTU9+gkxXcWYT9sUTjmh9pQ+CiPPRXguIisEEQ3/xjW
wCHUOuTpT0j2+4w5jeGY5LboIUWVaJXiNSXd6Y/I1QGfr4W+Lwmz2mCJHz+aD2OnxkhhizkL4psu
JLZTDhR+EOeHQ5LDgh5d3b3aQj6ckDipGfIlA1WbvzcBNyi8Fw8JEu916rZcDXGSfOewCMDwgNLb
20Zl3ymASZCbL+ozV9r/t8crYzo3pVTt1yYBX4sbJnThwpX+MdqraQtApEUysD0LBpmZ/8014H2R
mkXTvCe8SEQ2lnhCgdl6U4w+NfHqNQ/XBQNb9A6Aa/g6WMWNYvg4V34qBLDuzrlevSgqaLdeJQYP
ESai3uDEYM1c0Y+mcBgeVejpdUhk7jzUakyTOdyAn//xuFi4WfkDiGHPD5Di+k51cphLgMtCyJbf
hiRJr9JBUZ7mipKLuX2MEj8uXpwji2bksp/tgVE638arIKHS8FKlS/9NBEfdQTj/gyYSjtGQB0cf
4quygJEq9pHp4XSIKH0cW2aCY+UWrKi59aMoj/zIC3+0GeEaKGfc2JLZxTbM8oIePbeLBcgBqr0s
GkMDVmaetLVU/ydrsouppvQ7JONMkBJvNz+dQl1sRBlPmOq/+Oao2bXQHSLk/S9Jal8FyLE59HMJ
KXq2PtgZ0+jfO9QuqAf57vcpnNIjBEM8759wmzTd972kOfy8jmmP7vdlFwBKzfPcn2SXEjW63zYl
oRGJFP9RqshPDkWqHVhMpd30I/6EfKVm02y4b6xkHxxxaToYnKBYBmTtd+i1F3BwK4D0NEjNpl3u
wCe8uKJdT192M+1RXshUsZi8RCu+kkbLqK28cMPF20F4/IgdCDmnUi/ahnvCInPTJQm79VW0JvQW
8dNQPMfPNtyf8cZj8hE7008NYZFJ9+7P/ug6O9EkdB5EU3Cs6VUDjgejudtno7SfqfMDmF37RihO
AWPYvjfjtQbAKuBhvlfH3RxiiRPTtL0Xudbz31bWPrMUlNd20Yhwz1111cF5oLByE1Z03W9wx8wE
NyY3HjvryK8liX96kc8tkNGd3jO5XOnQftTUglbzy9O0naf0xvof7O+ajjKWFuEUyL9de2G5CuxP
TB16Dz3MYlgkdgzJWRAee6zUsfSEFDsxMhO7LV+1/UXFlue/tJKePm2yw4XT6ZffAd3jTeUtAlEG
TLJnFig8vp86+gulkg/tIURIDD35N1xxTwxgHHq+p3zN9Wd6UF1zEHS7PqB+kyRl7wBUUV/PSvRP
cc+CoNdDaPFUzGkNLoZNT7Y+C5PFJS2gMw/gZZGUdX3VmOtTgAv37lH+dhMz7Lma2GVOhkD3vcbY
a0mHHTx2fxz6tfo2TF4+HFiqgCkY56NZlb+CXmSQK0FWFAIwZIGDlSeQ/1cyYsNum51yCcZ20ou/
BELDaez3do3MrQrbYHSQjwGHEkfdOptVCBfm2MbcNivCVy75YRdZVVLNmgPiIV4IL6J0vvOfgGYx
O0IjJh/lUth+o1mLWALfsWEViAkzCaZTEDxAJ2JskKcsJjnSMc8a/LDBrKoCc8owrd8rvUCkb2so
zW7QNz779zQJ9xH6Y7xOfa4Fz7ythucuyNGQiLXwGLcHWjPJ0Zq4clKLVfz4EX+mfOuhOj2RVWgI
2BIXISVw2hZ7UIN3UMjTW1efrqG2rfRj0rXWULa4jwQipoBloHud5c6E67ANn3dK4lLnNhXPhhZi
GApEfyzm2dxxa/8DLEeuJTjyaEiV8xLta5PsWfklUSje6Wk5wJr4JZKr4FCpe6E2GimdKP5QL5cK
YMtmXbCycMqqMjP9MPAPlCd+NU/M+r/rX6peCgvqns0W82cuaOkxpdcjbnWlxlFrRhBs3a36IPjw
5YY9NIUyY7YZnkR3VcWnUumwuAtIhmuJ4q2eSIAInypf+B5Rix9ixfH2a5VdI5zTfx3k2b1EGO+D
GsQZTWeUZGMvlnr9eFN7CmihSUk8fEOUeHY9H37RYvQOv2gjPIkJCOhc2QlXNCyfCPD22/gryN2k
Y8WO5r5ke+gr6VT9FCHoah9DURncFiWLRKJ9wRKvconlG3v39W+JCkELkNaI/v3rDXgdRmJL4mye
DyOFmm0v4lc26AFqKE5VUD6/axIANkuL44cCJkQ4PRMiL4kN1Txnb8+1lbmvBqnjFHdvP8j/aA98
Bsimg4RV1AXgaKkIC7KNdYhPX4Ik2xnzL6SoBAwiJfCerGT17aicY0B1xmeutc1QjCJ5fCRT82lA
EElHRAw9loWLgFc7eyu969akeTfKDPBK+G9LOmfWlqhZB/A3441boni80Fzvy0iKxEjCELEzio6L
PWp5H/mk7Mx36qJ2xPdG55OXs6w81PoK8WrIQjNpoT2kkpsjSob7DO8R/zcPid+vY4vwzU1E9Zct
i9JZyVuC6mkjLA3q3OPm8+5UyxY7J1QYWDln2uxyd/Qwa0jmE2dJweIh3vQpESKtf+2Cm3OoHwEo
TVGX/aYG5280dedFiOBzurji4qFYxxiHWf4BbnwBTWqVrmoJxCBICzdpOxyqNx0Tb5cCmQCTi3/E
eMeXmhidAQnrIidnulCez2Uw6EaWoVUFVD4iz3MyvuiCjL5vefvSzyVYj2s7EU8eJ8VJOwNS/r/2
k7yPrQs1QaWsu8OPY9GqzNpWSvGbG6vSkmB29IaNsjoskFxU4S90Drqf2nxZuaiKJ77mOCMTf+Dd
WFJgD7upuw0KppPxQnjh7QFxBxYlOck23Wgftmcp1pHTe+aJfyyEGr2BTXpPywaP9OsDiym+VtAm
GXUi1oaPPLGQsD4+kuWRM4xwnxCETMvTspkrNDmc13eZQ1ytmHZw13o7mi+C5JpDAc4KY+mphpo5
3sXljqiF5rVlFfp1i2ees6XLz7G8F/jKL/nWamxsFnOWjATP6DzXNLOj4HeeWUsRQhZypibkVLdS
qui90LFWxOJc7GuoksdbH0q04f1zvIe08YtnaEjDVws7GL7Yk04/vQjwHcipqapoghsC1MTVWpA0
umLMsqeIFa+y0nWx/HpOf7QMQ2SYZke29qGWyGDjDKcB0nA7X4L/SiKMf2Bcc7jb9hoKpPciV6ze
DOIlruWZUGS20d7dIxF9TjtVN8xWV5V2Ejfr6wJzYXILMzwev5gQnwC5nsrVsp0dJhs1OCGQY9w3
x+PzmPNJRaCN+pE91ptKw+HsEVRS/cKchWM9DiHAHLmKKKrnF6P1DIoKMeYuBy1q0NlXA2ksAqTM
zKCOvH/a8s4pXvmrMahsStM1EmRyK0fuU9rH2nxJTVBOH6SrcosV/8GKrHfVffU09wBw73lUc7ck
9LVFj7CdXHVItnwUmxoZkvbhqqJvRSFWy6+20eIy5Ruk5lcxd2SJaYy5XvXx/rPVeZpoUzFQjzGh
ZwBwps33XUwxS9EcNc/cfHLaHPwy34UnaIkVMXEMYme5P7SwU8S5YC3bNNtJTM6tKCyDJVQdtJXb
Vr+qfajJyqp0VOyO1aCC6BOAsQ8vNqnpIeQzjhCGDHseZzg2ATK5jM2AM60AgntjYHAXSKPmM7I2
eTaX/NQSoIM3Sj4YqLJSBUHRf4NCT72OXZK9VvMyh8OAD9lwfwJ9uSqF4frs5L2r6CwuO2lBKai7
/085Misd+I12yClmh3onVzpfpoCcf3LG9GcWWZziBTeqQNo1VSfI+IfUMw17MzWA6ooSXpYpwKUz
zhGpaVUU5zSZt1YVfbwyfvqiWw6HxDLnXe4NzHCBCvukwygNMQpvdSszwe83lWq0e66gS2HQ3p2u
1+tDWSRK3Z/q4S9bNledpKTuW13mL9BAIOkuNSRh+ERIy5wrvRliDE1r5JzAiKN0s8TWGHruQGCG
TiKHS+0nbCl2JJ80D19Hs4uKS1+w3l265o0JhcH0niTESJftdf3UFPUYia3ji7mxbX58Wzxz1J3z
BBLVD7djxUYFureFCpG48c+oDypCFUZ5gKOxZ6nBcn8RpOOk7W/fBUlaoJjytA9F5LG3YVFO3B1x
+AgHgYnLbl9vuTKAlaigvcuZIyFh3XYvIlsQvAMeCYv58l2sfwU9qOzng6OIrYxqdvoSlzLPQVw1
kcnS9JjpmgKFVszOmVbNqzFaD+Yar2hyBnE8BNNzs0qYT9p1oOYRRFFvlN5F44lxwv1AZgyg1ABG
3lKAbDJp8pIFSrHsiYqezHzoK127KoCkbx8IklauADlW5NJTLeXkobknii9o/sBHnt6VwkUAXWnB
rrTMCE8ccfH0yAIfh0jykqYL5TqojjMRu6/Ln1UQHpynBvxvecuZ8nvGk6MqaBt/AQXcrYIL6T92
LypdKGxLpcPFg0JDNtbtYpR1Q7dnid449B+e9Tat06eAG4xLWneEeuA7+LdFOqMseKX8/FHH974t
48PY6j866Ey12GbGePYI7u4teb4BskrxHnVJ3+MTpBH+pc3MG05/8gPpYlhWmvSNAABCWsenSG/g
zI7Z+hFzdlqL+DkPOCDDVd9obfFnEf5CnmKx6G3SKLDug8RrsfMxPtArsZc9372IATtv7/C+YBAq
clH8Kjwj6b7LuRPPhGFTd2HWm70zfr3x413Wp1Y5I+AYXrgt/6LJicd0Y24uRwaSPf/jJUCgClFS
RHVq74GJch0Wq5QZ9k7RkACSLRPKEuyzAOzkE6kUDr+sCCLc1fVSUsJ+abNptumxs9CXNZUyx+Yh
kVzywYpi4k9aD4D2wJH5kiDplxmz+VCCPiU15Fk/3/2QCM1H8KWlbJShyJA/EQM5xclXEjtoHfxf
prpEKuMQCU8JrpY67ZC8/Z9EXBoQIaC50fzEYb0n/gTS6xNEp33wEguRbwd6jUNM44bpClSdWk/p
uq1DQ408XzYfUPJWKyPm1ajEsxTVI6MG1qYza4TH7mFRN2Q7A/e1MRMnxESC2V2Zf32IIeI5/vR+
JIghyR6EFuu+2FzwSvVVBENGR4IQEfrBlgWd/6Or3WbHaeSHWtFT0FJxtDj712RcNmoMdGuKAt12
iiQCrRtaN8/h0quj97ZyAxD3HThi0UgPwQV46Pr7rntxYw8UbsPAfNJR7aWIwLEHTRihfpE0p9et
2lgM+MgexX1lEYfZcyJVIyF/dQJzyh5ldUmVmo7AgAYMZCKK6mIsDDohepKWwhtEBf8esKqy5Imw
POSiwwxJ0RxUwLT6H16e8IJUcRjSKcytAR4q+go83sBawQW7sLmb2NJwZbWZvqlIEgDFDfzmgCM6
WrW8l2WVOmmu7pxsI+ilvXFAJG6L478Wx7e1X+2tPGt7/kOBfN/dRzhk1xWdOYrE6gcHNKYRwBMN
U8XIvuDol8xXcGyvpdg/TUwTegMa1Jlo5Di8vWq9KPU7nO4WEYhV7+oMy3UkshkXIJtCtTFszRnw
D2CYtUQzpkHGFWaCvEFsVRxdfyNtTqAERLOgymPOzjmY9SmdsQB6JKOjlYIRJUW5ECO4HI+g1pX9
AmMqf6T9s4AEFFhAjrRkZoAh5kZllk99uWbvCAbHrHtoa9P6gE2W8jvvF+Cu9pOYP4pu4Vv1OcVz
t+mZ83AdtPZZ/6sTrB9FrcIHWWB2KkkgvUINW2q+JmWu4p5KxzMc7IBgzLRpVtSN2A9VXCNPh5yb
iJyl4p/MvYmcYTJrNtxZXnetzRtXffa/OO8S8TEuaCXjlLxhsosUzNIhN4bNuiFTVCRs+dIpef8z
+mAbMvh9aooP+eewCWDsUB4ZjmyJ1IaPi1DtF+zmVnU2LDn9avyoNNnU5Yf+mNYRqV2siEpluchU
b45aRgPDnjMFNHqftDSFlDyvW/piEJ1/UT3HjpS38uYz9RymasgRuV87Vf+NfmuwGl8+qvbHAwK0
eW1naqpnQ2GA87iCIduwjNsj5rR57xDQ7y5uga72vUG/Bicoy5xEN32IaHNrrDZvODjsY3rPSTMD
Ag1hFA5DQi3yCArkHSPXmfkCRRbiHLYIAi5MdaS7j+kgRz6D7eT74n4dKcsWuhzXZibFNCD4o4I5
j4nRCJ6HMSrbb+rg3OrR010k4kLBMsOTiCEOfhqgg0q0xrkIOwSEDHIpm1NrFhtCuf0CJq9i4UmT
GnVDKkM0I8ODkaxQY3BQ9KXAHLj3Mk/ZdM39RXT16jP2JCHV7vVceR14AKmcZxsJBWb2gH1Y3Dik
NfnrAvrUO0wTJEDrePVrMNzQuE1wTJmCuYzTmFQXTHqcxKP4cZQbUhRqBF2qaF1vbGgLbM3s3rBt
E3DmT4G5Pfl02qsR4iBg5Lmr4u3w/D+JGmwM0Bn4ABn3goZuFeM2tGYEgcI1xYA/MKSh9fC7Z3rW
O14vBA2i3Y2lEX/2dHdywggestoOaSOq/iA+KqMB31GzheO2nEzsE5sk4ZSjx53tlD0ieUafSyNw
fA5dwik7Q4a0ephHZYlv+XAz1npYQ1oDl5Ny1oXEIVhH/9DLz/hLb3ri74trUK/SS3qqOE/6UWPN
xHndNDvMzXbBTyqqOULthf+aWs1idxGzsBiyYYK7PoLS8kd7B+XO/7YJWhGKL53mBpr29MqssjpN
GdMaFBpd5YQxSSr6rTbwIOf85Wsn/QlJr5X+KXF3LFQqV2jEnxmTwJ/f5x4CEteXvgstg/UcyrGq
DXMcYX9peNltyg8ykuT0/oBvBZF2VriZ8al9nRHsIFH9/hQXHTT3HG7lV/+z9sPkFkqL2IMrp1Rp
I/inPxULlijUfW41O69SWJyoJQzp3sI1Nw/l+dvRMexeMCMXxScmprhCc1Q5oozmF3Oe6ygCsn2Z
Vr+euVsNCQ1+CyWj30AEFi2mUyVCABdQu6Ku8qHULhDTTJBDjgAdHdyrDvA7utPuYhJRo+xq/pjL
aHIOcBP1LPtcpze5j1sHF1oG/l6s8etOZud63lKV/XpHZ4846xE/aLblXhXAbMvMrUavbK8QShCv
Vw+MwBAQZHPJu0yKkQDyHDoUJaDP7xyo0WucyeGhS2E4ia6FQwq8s1nK/oEKe2kJayEXN70YeElc
E40SWi11Jwh2gR0CVe9v+lab/VwVck3UJcZc4ECvPBi3XaMXVsvJ/nhlRvh7XSPoslYLSoeGx8Au
ZKWskGlmgA9vldY2d6vaQcVGWBVjOBkCKLxGCIBU7HriJSV0wFhFgwcA/GbXL7v6L8LR11x4Lv4t
C0WrQiYGfXcs9FFzJQVcApn8yH76sWKp78wvnyfVY83jrxfOjplbig9rH/2c/2n9Q1AwgQf7jeQd
+g4VXlCiax9DI7D1KjU0WGdfFDKH5PO8jzZ/SJJFQgyPljoBz8THmJ+MpzVrEFb7So5fGIGZVE1Z
MXQgWjfhYZbMESxh06xQGRNZnoVCR8CoBg55ApL9E/13c+ujIUPkbh3bpzdznHr4K+QZiWRWcoFr
r7Yw9hIV0dNv38Kju6cS/D8go9N6emDlzAh1fZ6vzNH8Chbc1+ZfbypNQciaFGif6aUeOmcCM2bh
r4cSae+vVI3F1bDplhA5RXL8SBvMkBnj/GBoA3gq2r1Us9jTp1+RkbIwT3wiYSJ0sYnBaeggSt1V
JZPWNgRuVe8WwY4yLCuJfHNWLNOD25ri/ZVm5mk30ysK/CKiTSuj1dKdHCw+Ohel3DEgkfK9qwaU
Eeg2bV49Jj80GPApcWhGsBfsUH6ZxDAqs1KvLUHdtZRjrKoTu+9M0R4ChaG+VuV9uXZXXsqunm09
0Ik0xWHbnztMVxPkmUaVb5bpstfHXMbQrn1ZQ3+M0yh1iK8ruGaplO6pDmspcLG5EMxxWKPNggtA
TBs8Ob5AzTziWPI4vPeI+jdhNqBEKrY8ztt3sgagIQI4hkW+l0Wz7k/HZGJOHbRXCQPM3DAJR5l5
Wj1HolkplsK6gHlgvkHIq1azQkTSSlFNiEcGiI6uKRoRDsh04pInDlyVvZuisYVTQHYQwFLzs5F/
R+DPN/rXGeadnBIpYLoqiNbZtdKijVgndXh7Wk1U9pTh7mbClYMqESCXHdSXCNomtcH0CKWWnzIQ
wuEXczg2JEyrUDxTbtpyfi10eIxgI5VAnIYP9BAlmOClifE2jTXiHutNtCvjsW2ge56nhOlrxlEJ
LVjMT90IaKwL+85PohFHI23DH4t8lBON6h8HPygIfV+KLccMP/p/+xtmVNObedCmS8Cocc2pLYCz
wnupQUEwanLPpU/BKQrgUwNa+ocX4alzMUYmFRLDNRGweXrrv9/F5GQcnyjU8r6TjWqOKwDPx4ec
8Ov1HXEXTBWVU/De3vSTJgNY1Dd8lGCj/7osXuzKnqRdOf4+uY8JKI8DzTTAuRV8FjgZz611ss7u
XDcJthcF7U7iEUMHLQMoDxKeQ6+mpu0kwoS4KDyoVPEF3E1Pqp03lqtlN92JLXLKFzh4M0XU5kr/
CPD2Vm3z2Zw017Pqw26mBwYwMGOOptpz0hOgpMv54UZw3QCyYUTTg2fTrVrhWxt+5EBQXLjwwlvp
md9r+VsDp8MBCsQ6UFwNm0MI5lQLw4CqmI7JlLgMo9scAfiNzyyHYmTieONI3W9Jyaihla9P/ZG8
Uv5W5gCAtryOxI8EmEAFZhDZNMM7gDWcEkESM7itUiTgvaFYTkN/3CGT4217oPZ8wGtPRnV/OTw6
RH5d2Frgx6hAIOeaXe/4cJmf31KG4mQ6IQpVz7LGJd+bwJYhZrihZHZcn/vztZedifOZh1XcXh8b
06GYuHUGMdA/UykCx/yM6Ndd/YNsB9rpY16CuFei9KL6xBWAI27pur7dfJ9WaS0mOIDVCcWrSwZ4
5fi0e2AxOgXM22h70jyuhobuFyyT1J8APfKt4mUJFvTRmdYdz2p+N4GR4jl5TE7/rF4Y7PuJs7/H
Xn4pcBdtt2L1SmtyOcwIMW6mJ+xcl7ukhM35VrRvnL/pj7LRRdJUFlJ7eOChdgyGmLU5BhMzI9uw
NYDjjzs1D5D6nHnGqDzD/9lJl3+X3DMdEHUVYkDABYAH8tmvisNEG4IKqd5R/LHy6SSOWbrKpDqa
NtplY3FlrhXoZm3pwUbfuVXwO73Q1OJeTZJ82Omng/9qlmbY2bVu15R4uaiXSBSclVKByDdkByiJ
gR09yl/VN5ZYco+pnFpECXPKUoQStfVErYVr1GsoyEIcfl4N/33LiOFSHKLC9NH4VHcSZcpKUMBZ
xjWpSPgcyw+S8yzjVW4N1FWHjvy4w2WW+xjJG0znbE0JhmvBdyNbiJMq76ZgAc53I6WRBY+ZaBPh
WnEoPoRQ5cNwV2EHrEvPOfH8ugwO1uNHJOOmAg9Dr1xGycnRsDNfwkmh/teMBbfVUrCESYugs/yW
LXQyscUWzh0B55vriAzX56vhdH+SudJudR+ptqDe53uAzbISCf6/01lvv78dTC5bkk0s4I2jIfMc
R1PQxiqXKhRMykHfyaJsaRujlPepQXu0s5eeMY/RNyrD8AplqKgSaSTGFcNx2j7w6kKRCvKKEVE0
aJMcIP77ynq0cOF8Quw82LkPMxn/Qt3kjiTlC2Z8nyhXv1sXEQh7Swqfi/0pfSW3K+yYO4W8ZWn8
tWcFAOOwIAvQoaGLgegxx6rrPZqRx6takoItHzW1gKXkrHGh34wv6hXJJDOvvJXjFPUWG/71tNN1
KUdtpESmEqnWdvC+hNv8bkQqLxWwgVqklCuv9xk8hIxzh1j9eTtM9MhR6SHXu+AfSV71cds0b7eU
yDPS92lxjaof5Y43GMqyVFIqEFE1tHjokImPWJnBvgrkmoKtwcN9or3Li0VHKzUnkR1o/aLd4n2I
I/X1OLmIvZueIBQnxAheplTsh1uLbKsY0owhiEhPosNG95GnKGPhw/gZ9VClrz2Bq317rqTBeOZJ
TZuU3/kw8ONvrDiRjxplD7h41UrQ31UkeZuFMDiRHb5fJJE916qpWpMj1K7/xXo5io5DM4geVfnC
zoxdcWcTXWIWHgNmgaeli2WRS4x8knelX7ptWuPecQ2sCsbdRlS76SnEVb+9ZyeFzTnVW6DeIp/P
xc9sV80HnZgJ6Z51Z5Ttp9R1GXhiz9YusFXd21cKii9XMCAJ/kVefzx0SN21BUXfQZZWNPcbEx6R
x2gNBdh9itFpshskvGQPGu7tlpAfyYUIFb9m1YHxr0brSIzHm+WzkofGFxRJaqzYGjRlzrB2Ef7y
St/eIYcPYZ7iIdQWYp8SLEvRWA2+62mHUM6nNunA4nxsgeySjgvM1VuPoidqgdkJA0XSN9LfkNji
hO5hm3WXuLPg59obTIRGISllE+h99Nc5KHb/Ajw6m7GhIA6WkO9q700MMNk1c/HPM4oDgTAv3hQH
KOtBjQQB5cJyDU7Jb0XYlDrMHxVQmbhmiH8y57BkWLP7y1TBVe7T2tzY5H/Khh0uwaH7i5eVlkht
fYWKsRL8zEBPFOVEpdqcYRxM3QN8BqGdyjg3JNa5kV+Ze/vKVdKJ76DrcxOO//ZtZcjBmLXlLtM2
tfnlXXz4X7GuCwHrguoXdtHTpukPwtDqM6RvGUfo+oi8qxxNRdGtZ/hW+UGMb+MBdXsy/h0CMhxC
ZxpcNDamD0yB/8wRzRoXldjvtfMKq7Q7UO/A2CmR2SqDpFaZSkNH5yIEOzcdpxw9kLYgoaCld2TT
+vqgD+Z3yZdUy3dXsmy7B/Yo5P4AsXfVY5iqSeKJ/5+tgji14a/Mn2bNDLt0oCvSGYC02TXj9QRf
YIoLoS0xh344KrYvyguRB74YBvq13vGgihPowY7PO8wGMmj/pnmEe7C26ImntsFOzrUlr0sLa2Sv
G3wQuzWblLf0G43EFI4pZDU3/BAkiRnlSQjyfPheqqCv0A30j712RwB9mUQD6YZNybqtB6SoUSS6
8H8Q+gOPCK11lU3y6S+upt0HJxrAGPFBovaXEK3wQPCCBhQJyujURR6a2JqiLv8b159tx7tBjYvz
BuknqzBKlY3RrNoOSbJuLH/ng420n9dFl7jsD3FvbWGeusHr2bbEPOSkJcMnR8aDkqfguJebKuUG
3nWQCHhI6wkdAHUme231lm58x3nWpqq0g+YFNLQF6HS6+RPUsUSEvjdkfs+6tHQUrYtmP1zxvkfS
OL6BCI07l33eWD7NiYgRlvhVQWzYklnai8o/xPqUXM3Npcmc7LkYdN/ari07NuVWLGaYvO/IOXiY
khLyncgCV/UdtY7KFQVS/Rnb0BB4vvgJn5JnoWoE6Fe6ffcNiosxnPqelxp70ZwkXq1zVZwd1IVF
jyUrdKTZt0MXYbDG3ygEE795mL9u/OeePeX04NmHn5czYz42KlUHIrgBj0rkbpAsS9JaZFXG+Zg1
sdkRhaZsKYOA4JEXtoQOsa+6qlEvFarv2duKKj48jkiXcELLDEgIdkzmhV6djAJl8RHd+10lHgEF
wGG9kuNUnutPC58MMGEKPBRBLrbPJqy/ZzAQNXMQ58pS32UgUmzNADA12hvxs8HNmYt+Q4gKLM5K
MnDSREakpg8sUi9TJa56dhGVXGqlbB2RVtZUmalttd01jF6LZ62lVCylnx5SmGd07asCNWmbMU0d
FrLFMjfkr8WUXHxV7lBao2cTiT7wF7VD535X/RxAJDMWiZGTAAKGpnUBqlmjJWsNjL8AI6ek12Bv
U4vClklOuCTje+KD3qVTMyv49c1xx263p6hrJmPa8dIx0pKs6ylRyPYuz3KysLJcHBOdOK17q0p1
BMLO8brWb3fAeLcWfptsbdaJ5m+Y5plLsRxmduoxCKwglAZdDKkyjV390Q4/X4wgYU773JLhzand
dRlaRp6+nyXC9aMn2O9EtKywLMtzaec3eWFD7vJ+xCyFfRC0svfspDYj6IxFtIOuF3Z3AA+55Gr7
ltnGe+kX6fFXdWeak+8j6o5VhV9TR57i0VVKvIeke2LiCyIzfvcFAveKr5z24LJoSy4N1YOZqGwA
qT/2pCKSOis8GrZpU8MvlVl+uI8k/jZfLagUZhVq5n/zcVvgpdwH6aXGaR4DLEf1WhGfGIlXx13Z
09nIJcM8DSU2MLLQBVUsgxCVk4BHHQ5gEYqu5rS9T+1YEKVFzVY/Nj8x404KX27yqVhR538Flnxc
qojf1VDlBxtrz3dxcek7Y8BJO1oQQQMFwMVXRUS2l7GGQyRN4TiqNJpJ4dsxSRE/qtxsoXj2+YKt
AMzsMGcVFk7bkpkIWrib0egUKG73ahNrRCvtxRI4+ujuzQXwHEdMze7Szz91RZ5m5ZUPaanyNbH0
Ff20HxU+DcLScUFiApueBAKn0Cf5Bje0peEKfNYRNtJBJGwd2hfTv8Uf3T20atxxbzHqXQ3wainc
BEStH5Y8D8wWXbSkm8wBxOklDx0HwVEowJLOctTg+aq8rcKYZAncjhjw+M6UIPrNhffTwxLD9/fx
CLWwiTTF+enOmSHpaZLWgB2Z0IF7Qb/x+mpz31YaqHEzhYLs43P0zeNHyRVelybDTEp4/GHMOLgo
2N4H9SIh6oHbeJ/aL4TGycJCsH5FLR3jL0CPtuHSsEi3/O1JDpKgD9CvaZtKUbgkI/PYXWUppEis
bXycLco7wfWuMR4JhNDU8FSYNcwOxsODs04zhl/u2KTyUgAFFd8J2zul/awDXsu5N5ytE/oQPPJ1
K2V0BUvu+PRyIEgkOfRDgI41fyPKOrpInrGewg3Y2t1t4ox8kLlG+BqvkRqfuswX/KyQfZ3siQ3L
KDATDvHgZ0q5wW1Doukm0jUiMUIWtpDForxUYKXljGu1lqOcNZWTQzJO3Sa+QPADS3zBuThWMNe2
claGOqzxU0OfutmgGFx4UpIdjA4TV/eYHHYxJNfbV9ZR8uk/vWfr1F7y1KLb+7fBMdlcHnhpjNQr
JSA7rMnuNpWLYEjhhHAfSFa9qXZPjp7iLRXt1vLS8gQND7pcdTasSvwUXoXe8rkf+8zHWUNkHHEo
f/cWVrSbru0xL39RveWqxEW/Xoxm1hHY4XHC9snE2h8h9dESeswZQWV+hjOPwEVlogMAFy/8togW
r0f5swTMp2iC5IE6JNYhNMEYJMkBIymOCjXgBbzmeX+i0wsfpQfZhTml7SFaQZ1ItZgX2HddWc3h
UU+oSdplugDhfL47o86L2zORWZANonYvCSN9cq0vbLk6mC23sWjFEK7xDSES138EOzw77NHT6G75
z0UpNDn3CETytko7+6e2eSRFLH35uo562h0fyVyOqQ93BuF8hAs9R/2ETok4LiW2Vo2SYup+CIFn
pKCNQqNZpH9hyxbwEOfxg0ILpnNL2mfTMSCUXpKG9PKss5tcXd+OMu1G3UtQGi+d6nBgb6z/Pn6H
w4t+eQYIaXVWZbytao2He68/ZU1XZJY7oa275FR2WYxiUpLR3nhfyNqDPulgaR+XhJ4H4z3XCxze
LWCSxkZ4xFtOPkcSmZmKBVPNAtBDkTfHrnNI2CYjgfxb8eCXnDwenmKjDqn68uhBugwKrj3XwDGr
Iez9S7U0oMDuUux/AQA3CJiNvtWqdnelatq5ZZ0N+NoGCvKjUh4vjFQgOavyEZZ3ORTlV/EnKQz0
r316AgHHXJFURS5xHfl0fN7anGTX22VzuxWYenV/5eSuWrIRBRewNZzskzPbSxkVhNXkE5nHexuM
wovJYp62ntebh8vqhlOa1Z/Xz5RNu8HqoEjcKCg4nQ67vpXocTAlMnc/ngXhPbG8y9aGfNLufC3N
M2nnyrIYavgFzFK06miTfEkgECOANiLYd45IhguAs3CjmXTrcAw2TqK1s/d1WyjRxqRSb/8IdBVl
ybFPePKzPvCEGzI/uikNctaXRHt3nlTakR2p8/gzTannzz+Ctpme7Nx5+orXClkRUhbtQCdItMIq
hHq7jMxzKaeXUkNWypQVCjGQhQBrdseb/csB2kNDhSW6332TOqxDo907Zh7sNRPNpCX2dufhbyqO
XckdP5IWYykkAZ0UmV73GzKzS6Gt9TaaMOCJDxOtkcgI2T87wdkpvHlJm3K/9SHms1fz8JQeVPLr
S1u8KaKqqxvZshLmZtsENI4740rk3b0oEhefleTuDKl+CljQ9nOrEUXNibsw1EjxBJvUO1rrK044
4LW3R00VsnO70CtXUj9XWJABke8aFsaR2KfVN2YXQ6rrt20Ours4ZGjn5L48U7NgWOrsnD2IdBUY
XMmrtSWwFVNFvIXJ7d0snnoCRGfj5a5M1RORgfNhTb9vCLl2JtzteItR16YvzHYUhB7HIxbt97nG
WZH8IuHq0YjTe5d4LEFJXR2p5mbR7rFu79EYwO9+FINGVcc7wHzFwnSJ5uoH7/WBGwvlZ+A+UstX
bEcu3HT+LdM/masolxjtfA+o6D9tae2lN71ReYVeeryZdRn9Y8ps5b8GBQmn8MV+h9zsYDe11StY
sVMXhmnBt5ielfMGimZ0qwJeCW/sV1CYOEL94mnVnYWxNFkZtDTYWJiakpVJvxOE3CJB53+J4xZs
BUUkKXkWRv/lYm3nq9uHOQ7XjVNdsA6iqy1NMRonpdC1mJ0cc+sxbIpxU6fV+HnRcBxGOfXvmEqe
jKgSZmO26h0YHF2fIg70jS7vlCO9+5f4j+5ji3phjOzYVsk0KEzj0AebndzBNTYKOQCYkTHCQig7
O8Vv7gJmOWY2Kcsd1GH6GTHbgLwsjKWic1UHHde5ipOpN68yetlvPi+X4R/l9rn+oUh0J/gcc5ff
n8opd/Zq4m7NYKgBGR/tOsW4v+Z7mRDN4n3t9rfK+PMzJknizE6BoKew/RhWUYm2KSasR/9X4Rfw
dfJ9vx5S1YoLRt7jeMwsUHXrJGY219PqE3opFVFcMZLGFVNVE5TbIVOKsJ0OM6aV1WGUHXZhrfaJ
mIMbFgHUBOgY/yHEZ7l9uPHLLNKw1R06kONsdK6s6mCYBAtH4dnjsu1gWifQtQKwzu6WVK0KoxIi
sSbWCPLCMow8jo2zckPtQcQHUsClkmAY4GgNbBfNfrZgvGP1kbjWLgYSM3e49kspBoen/2CjwDpb
zpFoJXZxw/F5bjs6zES3jjt+N+FW8LEEoabLZUsy1wKndNX22tjaRUwvCsG/AVFAveq5mOYtCUZg
v4WVEmgpq+43DxnWanRr4mTUKuPEz43WUL2xlbmjEMQF47BtSxUdbKq1Uf3eFe2qVKjax+lYeht6
9HWoEBpRBMDXS+qvma1P5y6jrt1r+aELYrdMJLGbkJfqY+M/4nf04YIkzDiN90ATFsgPPcPVeqyH
LJoIQbFyaxbiX87XRngUALxgETo7+8j4AzKa1fqecfibaCh2ks78ThiNYHW9Bd8sJKr6/zqKVADQ
EAO1jB/EZALFKnBTPF8R5y5VHQO1AmU9ZylIvZejigEvgRVkDxBK6fcJQAqepXEu/1m4ZY/c+L1A
jT97Fv5iwAJMZVxyAVVawbapsep2Eif96Otjk6ZeTfwGXswPBGhf8grTVOv1y2F9+JoSagnUrJ74
DGcB/diTwK7rWjGXK1lbf8na8f8mGlqbV66O5d6F7sf50I0bG9qeCyyrJqOL/a/ST1R9ZLh/GXTr
u6Nv89j99EE8tKb6FmV6tiu3LutAXPxGW8eEMqD8FlrXkdvMY/b3OLMzOSv2I2uguNWclR/dGRug
34n95GmHhONiazCMARLKQji1JWcfV1XP3wY348s6zfxXKUhnHjcO1q2RSEi6PfT8nTU7LDvNLSwu
7Y4vQdU1CVr9Ztjgm9uwNAL7oLcs/P0RSLgjrEQBFTk99a/DtvCoeRFybpCYrjRa/V6pReuNgMaI
0OrJ/A+m3RHyO0wkOECm9K6pXbmBho8n9f67lf5LfMbYp469nzztVJkZf+P5cKC0W0JwKkcp+8/T
jVh8foH6/qsGamVXwmCOYTI/15rD94WGzEYC7GsoKT/QPMqgZMEO9R3hWeXmBJCroFnhZX0KnWbI
RO0QQbFVJ4awPVcZNS8auCFmN2+bzTq9UJHVUMRYFJ0LHCZpCmOeXS+L+EGL+jrS2thgG7rDqCCR
xh+KIdIWHKV4WSSsdIfuGzrrqx3FqxHZy1/gCRid0nWjxLxgFQUDQlRnhHS9/H/AildJb+ceexOs
kBzrYJ9pD1nworh42lY4bwyb6pSu5/dqnqRaCDdOlHpAzD1iY5ot7zKCg/vb6/c8E5Ch1Ldzy9e7
LNp0iGjlzGjaoyaICdy+rHu9kurkemgfJgZaDan7Y/DtFFwo4hS53VtJwHo4EINVJvq2N2Uyk8hQ
21BX6ZT8YzH5XycBo+YoFBvQc6gRY3ZrXy3UVcbKlfHcZnGjwHcP0FSLWc4UAlM5mCr0laZSnkJv
tH4SN4oE2htk9FD1L6aErfSWyn0jcTgGIfzaoEC7wkeBF0/Qk7HU3gF/rvNf6cMEz2LbpXeTYvs7
UEEtK/C26FLPw4wfRMngra1E3Ms0UZD9O8hGwiwequyxx10eHgRcuQ5XiFsGSKZHapeqLaJ/XtMI
ltvhBEiMY21oDvRsgcMBqLeNACX/NQXYGse+crvbJx8pJ9gcu9UGnEWCDpZB7AHEVAXuKz5E+OQo
R6DISTy+PVMyHVzlNmzQWuQo6ArvhoGQluCzrC/eDEKDLVSFT5I9Ql0iKkgSKb2wVbQ+tOqabb92
PlYKlnPgRylCoeVfssWVKvZ2U+cyz8yJ3DT4EVjLklA84f6KTDCYTLUbs8M4uWLUyHxU9zyRU0MT
33INL2hI/bUXkuuUKFHiT9j+jfWGnVyP+j/9u8h6kd+4Bx1tRq+HGQXwjkLcHRTHftjgNLzwYLKW
GCKcxitUsdXJVD6a5+f34AwjnDnIykLVDyGI5GjL09ZGss85199joSAtlrW7JlBcYwnklBO5E2jT
PV/W9qLL7FGwB17drnFJ+6CxJaT9bGfeziuoofWc7E1ieNDwHpG1nqwtHGc1cjEO94BA+/+POVwV
qeGkR4Zxz/s2NgpNjUSJwfq708udhm3maVUfSB5by2gO+AdopeOWU/pjgbFH7xOunhT8MpPQRgYL
HqXS61EnLzBmzflvMmElZoXC3nymPhO6I398DuPgMAjQITrEi5ZpEa1I2zFF6I8BY2HLUy6wMXMM
k5GdFDXa+dS7rcnyuH0X2PSytXv8OS/dB6A8oyqdz1CMepOgLAjVx1C89vU9Nu1S0FjXOk+5vB95
WFZUszCo/kZ1/JO/ep9TP+SURcOdmZZSI6wOF74+f5br4XvsOBKjI8+uzzBOs2dM7jpBlbvg8n33
nVuuWSip+9Jche4qUIOlKccqfrTjQ/yRZHntm9zvmUFHItzKjvZ34N9BsXuPsDYnL0LGW2bBJx7b
kxjV2XEWI27FVFjkHF9emsNzsV0BmgMpAsfn1Wwm+mOTHLk9T2R4sORqxnPKBX8W9wMxiirjt2Ro
zWms1evrp5WxPBweHHmcsIq1bFn9H6ywNbiPADFFEWNcWU3/4KCaEIihwBRBuHTUuEmcaJUdJdVG
TSi994bAo+qewXtFd5icFpRPRqI6bQirI0g6eyntDI9d3PK/wjapjFXC1GiwGw/Jp1n3q4HLfa0T
dzVr3UEN71//KTSbFwSEoBiQuvOSnlJU/Ng62sWXPssnz6qXEoiWIi8w165dQXetC1qVPZYb+Ah1
6Vejpb+KFWmgBb3YNPGKAT0G6Io/kwa8x1qWJudpTOvUzAy5NREvqztYavYEWk4G2lqtOq+JRjNJ
qP7XWTB2GNIpoYh7bH9kMIrYiCOLD28rmwWN93QGNXxQ+pk/FuHNATzR8CbJBUHwJUK8EiBUkRaj
fAm9VPDe81iAB/u6cHQbLixbb8qGMEkC7vXK1+I7MCGgRezewOF2+dJR/VCul+OnzPVhn8JCuvmT
T8oA/hVTUFPP9AFgUmHwUln4q8WDvFAU9hEIpC/PpQ83v1kRuEB5Fl7vJZcz/aqa2L2jFmZF6ER7
Cdd5A6fLuLmr74g8ZBl2sDsXgn8gk3E85zpDR5NjQ1JOvflqumZgQmmxRAG8FO26NGoSywfAJ/dy
jpvEKb1Ums8LaiFCUqxvgUyuJh+soExMw6WacYixU0IZe2Dll0+BjUTB96zoLT8WCvBCn2h7vcsi
B8wscEMpr49pp7et6bxJEOscQ4mWK7wNygLWTvwI//GylkWVfqD3+6Mf7xnRDYSEjiDdLuNpJQhd
BIIOlg9adhacwlKwLcKwwleH6zloSqPNq1NIfKx3NYfTe9zFOj9tZJdncBW7q24I7vgUgZts1qoe
/YkaJgS/oSYwZ3oJFZhEen9i90n7MZTc/ms0KFs/XilHuYaC/3bXf8eXgUi1fKovI/CCbut4X8n9
ZMQY6kcjTy/em+IUOukyz/WAR9pUf8ZiYbRpTGUIZRrsqsHVe4sDTiNLOvdyD1qDTzU/QrB4UXYX
U6NHjhyOm7M3LNE05ToyGGeCs5uLCZfzWVF5orYW0STZmWBef+WArpSEfYQq29HYD0QqRk+sXKya
zdyAPw0sC/w0ZODlYeWh3pWqYb+DmR9kRrS3TFYLhlZSuBcy5+Ei1WkaKZH/bufXOoDpA7ENVkKL
jayZxHWlkNQhFWqTbOA8dJE09bqHEY7Mms1mU1GaypwL+8nMdQ3EyNsFYoIB3H/6LR10R/FX/7wi
8QQ4bbduHKsDUDcazYrI32cjiXjWC86VpbQwHT80XlOxynq+LvI8mxvSgEPb1Pr3Mn2kbbJbmGqa
sH6B+HAsWE2eD5eB2cWpoyEIH6M3yiwcCpE0sjIPVIaPyxyOlOXK6HSh3LAVEG4J1HkfonMdXQUT
J/36vneu9JBxjnqvdWb0A358HSBBuZ+2A5Vu29GV22FyexT7rPOgbY76hXuplnWQw54op4/zHd8s
i/tnnOPirkVtTn6dssrRJOh6vDa17dt2hDDNFjasUZTSC5SnyVumfvzpIun2KixliW/LUvZAtSre
SHuuiBD4pftYK8ofRR3IfzaIY2OmbXKyHRZ8Lvh3eW8NPL0vkXN7cqEjCtPimqZ01SWzIbmWGMQx
eavjKr6nC3ctPDrinaYmgF2zGjjTLeyH7mWzNsSEUv2vVJorQfj2OIULkFPWwnrO5L6Mf5x68mxW
EtAeVeES1nfe9Y4OgquMR3Rmme6NoleENgcuaacf8Xxev+Z9zNrVPHvT3ixUN1sQH+eSPE4dDozF
h8cP2iw4dXnRsv4eSp6A+6kF/p/+6Z3ciPv1/wG9uiTtxSbfvrgY+TaY/vfeKDM+YHF+JE+PNW1g
3KrQ77e5KcY5I6WrQ1E5sCUNFCQFFDOA8T9SFB2sO1KjtTpYVTrPX5Ny/B0+BBJZP/5sMR5ZcVTA
2LKxgDjHxueh7d9nqjGq5Acyd6r/4ODyFf3GVfmhfoYAEqeRYV3d8zmE93S7prUgU37GwJNfHLB/
a3wWAfmPSUff5bpkM2MQIaxbKFaU5RhkyhPDS/myhXEmHnSZ2KkiWQfaqD1sSHhryoCaopX3fj7X
1ZMEFPlGDGHpae2380JjML+BhgKXMXmLCkYg12flKNZMJd9R69kdgmQlP0nYQEqYDRG5vMTcDtBh
p5UwkkmZVt91cMx2G2mCLr7f3KuFKQuyy3+6Z0V4ZQ4O6H2rBeOqaxSS73t5eNXgOESrMbSzVh+W
cFv+a9UH8C/PT78fDfxT7NZkgO9OVOlD2wMQFidXeRuRuU/KiG8NNahhKCoP3bMNvNPyr3C7Wc8n
uezrvK3qlVXhQCsDVQJ2rKm0N5+/oT5raT53YzYycWcb60o6uxg4V/9BiqpAsvCXG9U9pjwoxlvO
dpokHAUK9VhH/Zsn5iM93KGVOZt+kDvRWg5TI8DB3cDPTeCJZ2SfQbs6XfERY9Jug8aIwOgHjSn6
l6Z9vplWojKTrIgcGXSw1qb3Lv2GtqzhnQpqtjtAUWU/UrjqcvNaEKZYUanzjZmBWDAvTWkJLbnr
z3XNsI7unrd1wer+AaTTOQ3UHXJUnq2Ml+X9RJRIEvUK34xSNQe+B4xbjzKraqYzdcx1smqYKYk4
GcnDSPedbubBu35sb+glDCnKj46UonxX3Dsy6aZvfQAG1bjKtwTc5qka/XclVzW4IrkK6Livu25e
u1YJMORn4AAm5PMhbOBdqkQSenGhx8DzohBuTl590bTdt6kkQ7BZVemXf4FVT5cU2TTnSFqXH+sz
k9RXRT/p80RoIie6xuiojMFIfnieoGjOLzvQqVHvrpioGqCMd270l+y88iMN8KUJU4YBiSE6J3E4
y5nVhCCLc2okl8ii6B0JYXhS9LUzwW04fmxYG4vJHxz3jehLz6AzVfe+ZYALDvH+0A8rQzkxuzOp
x9jzkt52z4peqsuNQ3jIVr2lZo0/IINlcndeFvE/FktvDziZEwHb5ika7apIN8ascqLSKMGTnUVD
HdXHLqqGncAGIBhCux3gh9420Gebx249rUZHrr/Mx6zlUkSns6sUaWbxDMNqpvA5Vnwn3ocW1IRv
pCxpOjjZut6kq3nO6qj+jB89bpJi12EFTsrCR0bLEDViK0gA+RQm1eQ7JtJ2CX4eGyQD4wpQ0szf
fbWUPbl7AmzBIxpCjOzO+sRZPPcg0VLPUyCLBQvgSmg4pTQ653fq+6ZypRdRoylMkIzS5kRl9wcF
qE5OElyx+gIe3gTN/YMLdBVbu4gmlQSFUhZALHWKGVC3aekmvOecicSjjAxOBMgs2HdhVt/ZPAGk
3jhRYLbjoEWIWMA1HCOFdbh55PUa0BYqyhPWgOsMpX6Mdr/PtMmxnRHfPIwBzyIV+gZZnxK4IxuV
zshL4UyBM+x09yboBd9ENAj6HGDppodpK6X4lFNSpsNjN2xF3lm/+RIZn5E8n239QWS2JoKo4WqA
Oqp6BC/SDMnDG+9cMkvhzIoX+Lz2O0KW6615Zs5WPtSa8g6j74Wv13y3pesvxkz6RL5u+onpxDVp
VvfZrxaG6tVyCv9qcJGmNcMNtn6LtCKJDaeSlrxuW2Np40N2DPuO955TbFAM5ido1Ws/NynoHmK+
1NInCfYptY8QiMtI4S+ovhKwJpNcsu6n8w9zrUDBQ/L7Uum2uEjC+bI5Jfc7USxWuMO+NvelCAmm
seiujlRhxLmLOl6A8G7bXfQFDL3dYzPP93fNdTc43egxfMA+YKEFHlMZqXJ/bgfqG0Gm2l1ATIag
FpIjVEE0ok/EusvBvSIbCoEDqNMGlkHLdnPWGBgSaCexVJW3hn0YPiJVkXpOnf8lKYIWx6OVDbA2
aWgWp6CwYEPiydPqSxORRNXHnSUss8DWgO9nrRIOLhp4EZO6jLsagezBcrmYzyIgxuK6UjT+/Gt7
CppJ8qiZgP4A78GulvZQx/GFr3H9QDBpCLeitaqoYQDev3VPUu9tBMkvKbxIdVDKDRhpmnVhBx2b
Gv80K7FqaBeTvguJ3mo1ViqbS3dM+LepZIf2YI3nN3zUVyZ4Pn0HVFlQlWTsFbc2zcAy1844tbmZ
fMFsZfv37/ynR8Ol0PlsLeLFj2hFltX92oY3v1pZsSK7+7jdXD2IWq4cVYql+V46uPYbz4rIJQmW
WaAgE1KhiSWnzz9x3DzVrsUUS9ZzFsIdV7GHEo5xxVYzcxXvQQeA0Zz7+G1V9zU9Is24mxb3ghpY
3M5VkyrdfCtKU2XNSHbW0HzqmLJRlZbOVhDdTem9jyQqYGDqXKUZ6ur9VDVMSHTAGbfUn2+VvseA
JHrecD8CNO+oJK0/pqabau4SGiwPC6G/I+12hH8NOvTeh0NlBlfoHDzH+p9LBHUFhooRo7zhnT8O
OSU4iQPE0riyOU3ycGz5dGEzVLMGBpbGpchcSP2uULS4atDyhRd5LBURANkuNSQqzBqrwfhWMQvT
KsjlV9YD7ewtNT3tuTrzxfXqp9defQzosrVqrVEIHe9jB4XVQ9E7SIJwMLFmo7OtQFYs5TmNZ4x2
cZHGbeOo4oaIcp6HHmEocXWlwqVu4rgszNp1RT41W8CmMsUNvNPmnaYzLJPDZIO94h6wbKUpes5E
miqQ403EtkcU6nz3aOOuHsuhl10Y7sPcdP7U2HhCAsPK1iI+ExKZ+t1zRiCc0lgooxsfuM1axZom
cY7KyMiCgfnXe317b6LeL++22goFlYbeQToDORj1vZEq/6fRO+tbRCBTFufrKDlfmX0NDDIjuZId
wwn+93OM4JRFJBpHbReq6bHHM1WyWPfIPeTXUe9KwvZZaaDVgEF7Hjmzv0NdWgUGgDzDxKoVnYkP
ejeRe/o4qtB9h8A7GlUYL0A0a5c8kPWq5NLww0BMhIwq/XgeO3XONp2KAi/4GaEdXbYc6Ju+vv3N
+ePRUAFcuz2dL9iFi0H1VFvG7d4+oAZkrjasQz0JxM6ci/UOET7USCiT3lVDx1a15CLGd5piE0lj
ykBIIEy610sM+FNgSOyTllmmWPd8w0UrlKqS3FAeHJFIlvnpQo90fKTzG6+vk0gkrAy7HUuuDyvG
PUStWL3pT1SlkJyvR59L8bV7N0Ku2Lu50uqhSRipKxIlYwoEAqZFE9UM+IfPWUiqRdbacstfEI4o
p8qdA0D+/NP39OhQVm0feFGGOjOuOElE4xWVFh+kfdoEfOK1BLi4iVBwMbbpMDrXFBGNU89HBr6E
KmZcSfxPKbESXS0CK2mN/fpnX1ASrVWBH5W7WFWfgKXd6tNkw2PJuulhIMK6+QbwNLmOC8vvIExv
ejsrH2lmzEiQdFTzgoIXYlOChnLtaymwNClR3yyuToINCrfvxjgHA6dY34hEMw1HNe+XfhtCiXxQ
iJdY0pAOZ8OAKdihTS4eleuwhPevAQlIYN8HkwvI/VXBxX6qJKowsN3YXT69WTeKyDpLh7d2pJRw
l4fUzdyZ3YNKHzb2RDYscNmLHahrp/+VrKz3sWqwzVM9raMtJE+jlMD7rKg+V++pEXHS+U8b3S93
KimBPn/VAxIm70MOolnFdjc6YcU51nFr11xvHpxrbEcXzfYYrfEL0c1zMo6d2TNRt7ogqGXNTjoQ
WglFUL58WZUavvzurCp7InTmuyTkeAUtQ48/P/Z3Cwo3P4dFH+GtOP/s2X7D6fkTWW14LCtZFy1Z
b4XQdcjDRZYZ0IC/0UNIBsDOksDKxshMVhYLRnqpTAFZUh5FGnW7ZgrcDB7TWXWFa13m9I0Zn+Oa
N8Qwy+DFinKnBSSBI7oJv5UdEjx6zAt1pLTq0avcTK3Om7BkB6LBL/gdxAFF7tvMPs8a9YFN6ois
uEQ47O28JE3y3N7GTXkNVVeReXysRvS1m9fPCpIFGHQYSzOtlGx70ceEbyADL9VnZ0PR2vBoS6h2
PqsFpcRHI6/7r6CB1cMJFCbryXRCP0BJlU7kIWIFQ5bcNgcUoOShdeOXz33z4Vdcko0w5NskrShu
ygbR/n1zNjZ3lFyXbHtH899D9QXmkQoamq1AnjiH+eTrSLOzh/dOLsN+tsGBhYqJlxugIHPtANWH
W9w38J7949/Mfl1diozy+Oiix83ojNigKiK3YcRn+pysrBxer+8D9kUl7qqYRG7qHUvy7Dw1Xrrf
1KThbvf6TMSDG4OKrz7HQSx8mGXp3IAc46TqtIpBkcZg1Mmb0BiN8LUReCY6uU1WJ2TP6oXTAuyC
iijl2oZh02Tqp5NyZjQnFT05n9WlWqwD1xsjghaqX0k/gK4ArLWU18oRhmNO8EFkoDDlHrmF6wGL
0ENLHvL+82xo7Zn5AJbSfx+YngxiJkVLTEUZCBGH6lIW4FBsnoOpZXq/mFKHXp8L3tfmz48y8G79
XNy2WtRgst1MCLRVWNWHB30Yh1AtiUQ/UV9zoltibH4bUdTyZwxlJa96sOTYVFiZ0bxGgJeU2IFj
Ss4sCQaq/5m4aLFVmfM4UB9aiNOPYOzzoBBjgZ/1LiwBvXNmzeCa+VOzaaLHGzSBSPOkO+TBfeBv
UgXa5NMNlLzaGrP72qO6c8K11CoDZoFfZUpj48pehKY4wLyhzaSKwzSCvidDDuuGMifn76oFW1TW
nYD26QfP1ObMyjCNE+VhYLgKg223l/TOKpsgfizLFr0IDIcsllZ34WBV7YjkY46yXnn1HY90Q+TX
xQAgHpUQo7AOQXANFNE62YScuVj/C704n5FU8nnLHFOFMvTSfOWQnl1wyDkiYHhYHdKwfTJDK4G/
8hftZ/argROeiuBya/5colU2ymaeXxxk2qSm/RiVksKSS2cXjgcN+4YCA/aYhCDJDe60QWuKaCmt
Tb1rlvff6MuzPRbVHsn9PQJN0B4DOFU8isRchnAg1/U9ZYAaVqLJVR32xukiJQDGRo2cPs6WEkz7
8K+3FFWPXMbI7GUIIeblJtY+VY1cDkLJk6QhFkYESOrItM8Sjle6e33wLYd0vBVOUBjQwb+ozCBj
VugC7wkvDf9hDs6opzhOwFRpRKghr1yyj2Hb7//tcOaKbuYH4w3c4pjR6tk65tbh3kIo4hqU54pv
iR5U8SBEVMayscddOsgCLsg7bfy37p5Uqg+Dt0IYRZ+XBo/tjcgI982tspDBSsToMLlituhuYKBO
Bx37a/qsGESOQOcrXqHdh0D8S8pijik5DfP8DANjXohjyd5rTArS2/N0HbVcubiPmfHj99/SnKml
M4pRMD3p2aa5TkhTYi19s7lRLeMoy423cww4On3rV0v8+khBMTohgOYTNF+5KO+Pu46Pwxp0wRnz
ZrXxgEDBzL+QQZsD3mCxoOz4Cd7HLJ4sk7hbyjS+SOKBrD03oTTHmKQ2Oqw/3fmjiNGf7eiMRfn+
d1yOrq9hk/i7wn1KQKZYgFEZLDUrfmcVXN2GaLBgN16AUUf+QAhON5/7g+SYi2kOdSRGn0YUl4yk
1AtXDXw10FwBa1HmGD1W8fpeOjoHj7RAls+7xu/ORcb/RqR1b8FG4XKCXZlyPLYx/ZbkocOzdV23
brsjLalJf/lDNJKVPAw3bFrdjr4gHHekPm8+0Y6/dgJGGX1E8ftSmYKMEJbdzu/gVke6x9G9Fkvu
306mRtQcmwrQRafs1xBscyoIphpwSGz5ZYZ1KXBhUNntASZZ7tbqxpBkr7lSoaIPhUWvsFNbbfnz
cxbs21laLmJ2h7Bf/X624Xa/Q9QI50LzJdReLoOizK/KBNpj54eCp+bA4/JMJKrE3g1Ls+SM95pB
p9JdSJvvcQQyfw99V6aOw7WrOMI0Hjx+EdkP9eXC+ezcz7WCOOFxgzx7pdre13pK0mV0aAPdc5BJ
RmRb7Yjw18dOMH+/ejTfph1Xr2XbAGL4UElPaJ5eA8aaJDR+YXCnM70NV2HUQkEfDK6460oUsyjD
pU151O2EjFpKziF4Hn3PCNLny8WX+lZs9FKlJZwodOgGAB861mARsVQ1ZNVC7OqxwHoUfzTXma8Y
MTC6jf7Jim3vK9PU2v6PncsP3ylFz9/ErDkWo/ChC/MTV0evqNVhkcv767RK4+5j0NEsIhMkQ8W7
J/XqnZtepKM2l2igPBOmvhXzr/KM6AtSWyZ2ycYGGgiIM4xUa0Fk8T7SO014rE83QSC/4uCLTmMh
a7SmWyCf+WdMw/7g+F6gODCe833HzPRHRjpsSckqdbiXezEkI8bHgRxZxtbAOW3PXPZ49Ug9kTB8
hNhs5K3wawoYGI+p6PbawWHdNM/Lv27ws1Wb4yP2phpTAm0VQXpjdGrAUnwVms2CUkMu6JEUsyrs
RXeL8UFJUax+s3fXFUsySLeIWwS9T9Tl7MYx5RpA+TOeanCDKiBGeQIaPwylz6VWrjmjsLc57pe2
tou95RkRgDI5hgFeL7KzSvEfijHeXd/ZTFf2/9vuuPPsFT8eITlpXTuSuRNxpStSWqJNO/4AiVVx
sUJscW7wKsabxxKcUS+iu4yTprCHXi5zIKAZLe5v8u8B1QgMm5/o10rgNV7KKn9bSgk7ZesE9Z36
qEFiQhstW80TRf2oJt2qQRdVYErIUZmaL6IdS1s+6mrVbjTE5cIEJeWTKDOAc2KBAhZpqL8gpo7y
BkuUqxRyeBVkYcCEyZGxA9eTZWnHQFoaNdICIeudyI9F8qSRkf+8ZnGcfbPV0wewkxtPjaHHhDWt
QADqmmDjT3qgAyQL6a0B1eTmihHfY3oH1+t5Pj/ctygZsjTGtvAsmHEClhtLi0bqsx7AfOqPmisM
tdhyCi48rmhidovzQ60EP0CkDicoKiP/P1UkAN87v7tRIMi7KUqnZSMwOT+rWGCoerCFlWZw9Qdt
KybfwnRnjLfTy9NJkH/ek3VgD8vNnvOnVO+0nY7HN68mDT0RnMOMqQX6xyCwsATWqewbcLoJEkKP
uNB77mNZTufw4HdlkQW709sIITezuxkWBom0ucJBFHq+wovPBsHdwxu9RRVm5K+bwtmWTE3IrqK+
53KU5z2tT1JXN6HoRSvJ3sxogKMVA3RX4XrRNrZJYcYr9GgTBf3BT4YEeBI/y7IPopdMoiyc4oq1
NoBIpviTC9t6Rbwu1TwPZDYidC2Vui86+KQRMZQgv9shp8tOWgTF0q1RKDQMrhBp5F6gdCDeGn1k
fKbWpJ+ZGtc5FnJvJA+ao30HN32sngPpUXMcJakBGy9vKQu7eL//ktTRUot0SHZ4mRXLCVdVjKnl
JYu21M1rIr1143keT5q0Te9wrHfxfyHZXraa8Aqlueh9UmT7BNlXRBtBk85QYCqOvAxn8ZacY68s
mPRBExH83kJv3GLAxf72ftP6tnYpsuPxZ9aVEcXd1YpyfNVDBQpWgZMBGgYQvMJsCu9KgAJiBpO8
FUfGyFef//8yK5c29NQk5051DdFhbcckcGEtYIv6LEBRK9kNLAfAbGix37VQtNHuWgtiCu6s02tS
dxullUaLzwImtzfi7QtfSVJOHsUROiUnoj5cckNgbSyYBXM7AkzLq8zkHluCV2Gnfo4Kt0TtgD3h
zHiXOVjsUcIH21V7JktojK0rFMD8UMJUD9gM3J0enTqKXU9e1BKeo2XhSXd+OjTrv8VzTkQD98Ir
FD85RxTKdtdD0k0vPXqINuMisvb+pWtYhA3Wx9k98O+TQbsUnPJW+nGh0rg3/7NTz0cn+eCwiCJ9
naZaWnpKfSpAEt4A4OnoOemSIluv1TclompO5ga5fNWh/qIMP5Q2YDBy9pKhwUDcmPTZ3G9Y4Jzp
KhTpkzOarXlYPSGms5sNOjVV6eE180L0gsmuvVH/KnH7pfiF7UAY2oT070557RJbgLsKHdEHbjkh
Z62y2wM5IzXgIvAzI069NLRwVmyStsrapvPa96Ug88vg8SuVaAL4rZeFUeEdq8me30EdvLb5mkfL
Ul1wMpuirl/mTDVNsy9G6QMBd0H0JTw1FiwuuWqiKfJX0fcqWGarU/kyAca+4XGCVkWN2Np7U7x8
/R4lqnTIPntsDACtJ8pCc/7kh1GdmWqZ5MBMeLvD01KHY+S1aOF/uW+aUsaR0xtStKzkkj81Lsdi
c0GcFHkKPbkcbsEmLn3E3xKZPdGNshhaCHqK0der+3d2DK58KMrQTIhOQkaW7jhoWWyVDtPhaD7v
S8YOdbPdez+UPt5TbsfQb1kJ3fnobFWniSpmMKXEsXAQoZtk3DpfXv/aNTXKg0jqQsxGUuYIbdZg
nmR9tVErCxGYdFsfSuCBL6X/7lpXVcBavTrtAd/HTcJ2tDoYGEH2guwFSgigwsLWq0CXYvWXvDJT
jxCkvr+sqdqIMc5UA57m+UpwWWJFpcsT4l9tak2TQ35UHzuEwC09FYMVIa8Ezmes/1lk3VQIFgzd
Oe/8sRbJ6UsMvlBPoC9tG6j2cJwO6oL+7T0OxFk0hLTcDonKfxiHMr6oqRX/ULZhuYoX7ZeRYyw+
hTmR76OpDx425Du9hAbiiv0GxlAMBEla8ikKxEUeZ+zO4MVLdPLWhQ0kYjbh99Pscsw33vb5uCY/
LXjb4H6a1UtdCCwz9BRRkZTZa9ndPWDX9fdmKxHcG1Z7JJPYdDGhZJn8RPlaJtswiswq2tt+jWdb
U5K6EiUtpUin9lf76RoQKL7uMYTjVonbNnLRFmwY9fCKrn+bDOTDJ24I5ffY5FLXQKgMup+W8Nrb
Xkbi5sWTzeJTlVJF8ihgVVK1bP4E7Gogtv4a3qSz9ESgU5DF9WQ00BRNGQACzLFlJybhfyZ3I6xf
IEb0vxVL+PfdazVLHzngpG010Qwg0NeG9AAI/d16qCBjgZdEAZs/Ing7RqjsSlWuy1XbWXHp+xhs
t9CFwf3kelobnZjT/1zUonI3qhSP8OMgIeOdTK1Zv+7UyF6WLLcpPu99MddHxy6ViqFl+fM8K+J7
ugc0I8uzqy+f5qMWaTciQk3kBE89riv0IX2UlcX6X+HvN0FJctIXCfIkr8rtZxELZJRWgfUuzYbk
lpp/0DpgKNh/ZJ4tdDV6jSb9Ya1TFkXJ36P5fL0+4y5Sw5ebv+uRKysxtA5lzRq/biTA3zgsx1Uv
KF8FSeM4REmibG0XAsu0J3CHdQSd2UXGwi5t2JXM9ehQs1b6gB7JgaVxdGRcvoxDPk5K2+Gg5ED0
oF/IwcKCGR9qKlxlGhe89BnAJ+iuE5iXQMnHTRR+9XCjnsGJoTz0iE0M3WLIRR1A6ft57KfiwpA7
2XqqVig32vVFm/ydvs0mwjgctiRf+kLI7obPADVSoAzIG5zwYubLy8zwCotRAZHUvHUwMlG857dW
N5bucQY+1t4mQs18dNUHFF8HItB4p7dzrNVLcuxhVwksURrR54GLofItWrpW9/Nj+vuDqHa4SAWy
X7On4i4p5MwMC84mr+tC1MJdxiKs5dOwVcANuFkJx2nF/QJy7fDfsBubyrNFHhBzvSF+ZXTiBSPo
psRMOYEjO58aWc/ZLJcutDoleQVk0bLHOA3ncm6qczmVz1TelmoKodF7gQOxWwLqcnGR7PINA87v
qB9F/BEAQXD7ou0H/KAHGKZjF+gH2J623JDGLmr4LCvs3I/e0/S2eTZKq4TRNfvVrWKXYVE+1MNt
V75hdPnrBDOzbUdcUbugR1sFS4uQXKhyCaSaDIEPoR7y1JERk5G83NDKVSAz9IjAhfdC2FoXOO/Q
L3xSwzyI1Id+LstmtbNx2hNK/VBg3MSUX9puMnDJ2auSl9XU/mTGspMc2NMVvx0oPWpGhPLDpjeW
jcq2FsgfwGtyZokP5vuRe2CmDh7F/z61nd+0zIg573mOWF4KIU6KgMxRtMdTh4LQjltM4snmcHEH
uwA7iPbCyASy3M/kaPJRicFRe1OCRpMzt0VHjxzUsmmPnyT6ibgEX9McTcklfSUiQIG4A9LGNSLt
SfXzvTobEfpauknzvnTrgijenZZAM/507M8BdYbPapdOB0ix+NwpbBMIh37p7UsNHUIsIZgnZCYz
HW+/C23nbQeqltzxeu1MUJBMdD71W988yhYoPytI+rePFcUM4b4qdm0zE2sJp+ppwAohQRMp6eYY
nmTIJSs3xpZ7JrnVPnxyDNfmxaLvj8HbEYAfGfQfaKB+nyotsKlxtXiQmFaFLHUOZ6Waw25u1DM9
FqQ9z/tkLsChVDDvTJQp6IUKvb1ENRhJEaVPmyRHPWIHZ1zgBypkkRbV/K2qkfVAAJXOx5SZzlJL
hE+TMLsN2WKwnP4cvH0ie5OJ0zcn4otSe3/XJvf6rn1eMEOgwzRzEtALz4qoG7q1rhhDpyITHKnB
QNll8gJTA9mqCRygkQnwL4xX7LlNIZ4tMlAzP2sv873EtZkbAmcNqCdVj6irL7T3+vx/LtUyB53f
31/6O8QgGX9XbtolVGLvpn+3nh8X7nKB5nJcrx5DgyR66gp8L+TzssiVqYcKC/lYLI+C9jH68cOR
Hsg+0/ilq/hBBFFt4y3WW9C8gRrNAonaMRCIJDOPpOF5p/DnQXB4cJSeHBPfMqYNVvFrlEJzGTfL
5jx4FrHelJBhL6LXOwOodI9zv6+RrR1Z8kwkduUSNeME+wBMnDt0AnoiBcu3VIwQn8aS9UMu9LK+
y6j+f2rI+TzsK7RzqlLVKKYvjOTxT6e9zXTFmL0x49k7UEivgkdeA/UWVs9Qnwc61K4fyY7MtDhz
X0iBjZKqyfbUaY0C50q7G9r8i5nGZcwEEPF1p75ntVoqro/W/r2PicStL4M+1vAmaU/WFLLnputJ
vDJntmBYrvaOOp5+6vl0/IW3VAnTw0IHko/sem8XFJVGFE3Vr6F8KYYMpfoIni2hSmaWk096w3SH
CsXPVUclgxQ8FgnMaqi/gX21uTHq8IKK/2EhCOB3YJ2pH6+rvqp8QwIu+U22llJ9W1XdyePEsPBm
wo4quQ2HoQEzwsvn+59AxtvoxUamwvXv58QSfE8O3yJedQLT3dWeZNP4n9ebVaPIcEekZ3699Tp/
GBI8kbl+e5KVj/zUifAMgtqoyXZmxiEy/AxUeiVSv0GQMSQOdc0xE0VusO48yO8GUiKIYFOyv/GE
aOTuf9jhVb6k1TRA44NM2SE4o0DpEipD7HU3UVT9ZGk4N+2U8r0S/AKIwu4jtytCZ1StzjesaQq5
j1cytEcCFX7ctqAL+FsBQThCcEDymHUF/nHaEHL4zDhj4KXHGcnS3sciwVDr21LD9YHBMdun21lM
ydZ4VcnJ08R4JARkERlQEs9+Nt/9HHAqhf9QVf+JVb2XtU4T7F3j36E0MVQM/4D751Q24TlJ4fnb
tPzoGiZ/O/IUDE524Es7Cy5PBJsbGUyBj2C8iNGocwa5hg2f2XPDdhRt2NGUCKtJ9UsNsQ4eRPUC
+QH801VmfyNMm0xjD2+DzYjKaRTyYPCuiOxdeAka+cgvq2puB1WcEV0K0H94zn/981spAwFgokya
S07Noajg0rdIWddNZzAm+Qj2VUHomofvjNVRi4dqAgYLQfe+TRoRehupnCSyBpdOHbFvy/+ugb5D
vdzUxkGtbbQz9Qd3OoNxgn8LkQl9eGJZSOh3x1eT/IFX8VvfLb5tgoD7ihXGWBiaETatGw1NjTWg
XD82VQ5UfPy9uWSu/q5uDnKds7HvmFuxD8NoL7BQgoRf8fLbOuJpRbUnLpTQoEd66Aqhg8K8qVP7
FRmncBFZktBVL9aIprxxCYIpoouIAYbGr1WO+rYOwN4uCDZi+Mq5axIUMsWeiI7rKUy3TSmRFWkZ
xDZDQnX5bMkxsbOCCHeZ2OokgdxcZesPKQ9qWFpPZM3rJDj4wcm5udsTcLEfUef+df1oOYK5Dh6U
6rAWMcK7ZaFJ9E1fwzyMWOvy1c/UvLmTXxXlgvT904Mh3JvIYC/C1BhDRovOhoyH4hGBz4OK2YiV
LPOZdMOYwO/TxsHo9r0gqAUAWXpR/Kv3wHRkX0ioWdGotpFhrwe+IpYkuI7WwBXAtiwdvNFtNly1
qBM6k23nl5MNCYYEB9mAh09/xn3f+GmM+9jLD998nvSWOF2TnkDQw0L0BHKauHCoa0gDQyu00tWr
7Czi2qOUgI+ORHVxWdOggvPn71Azm6Q3cGSDT5PamoNqNC13y1OUtSmo+DDPbT4PZOrESnmeq/b+
bdUMChfuJgZl74oZAsiR1xT68WySIm1wjrm2TW0A3qqav6Fu3XCudIP8MF5W2QQW5p40WEParQ56
G6nsClkeD7rY+t9YgfuBKEeQnIXiEgrw41AY/JUxGQJjHfI0jwqSOnRqP+v8A5+pI8KrQk4leEL5
eZpKaBVelCnLJufZAf2dBTM/wHChSwYkk7XYhFuFcnLlWTYFK1GL/3XSreDaJ4xdZlLdMChSYEEq
YrX8DOT3A++syUNbkIozTJZHvDar3qqkJ9U2MU8jRfIMNTys5NNuH/4s+nbc//tWeL0dEIVftGVv
AR6HMSWubQUbt1g1UUr9Oxeu+cVlU7/WPz7OK+ckVpPjmA4EyxTbnARmW1rx18k4EMbqJShtT1Dy
H94PweWH6nOOD3XdQ/UaCTGREpH37eOZIHjlejy8TxhnmzJHQiFbcpr8yAjZYEEVbc7u3YKYj6Sg
7PGZx/977ZJF5ZI5Vcz6YzK4cf9wAotnVg2boJ3CMR+YTh0zBhvfjeE8ctWdkhO3wl2VdSvLb56G
QFHVemqjQ+g3R6/Ix2V/eXC+yyDJKBuZJOEUXpw2qlRJtiVMXV2HzsjULovNIrh+r9hCo9S3sAn8
5+JvFmKxKdlC6MPAVIv3BAsBe7KRph64CRK0wm9ZMPlhUQNQC+rwl8gMInG+ah8bjP+TfMUSQjXK
SKwv5IkNCv7venQSMwazIeR0pb8YsKNns93npGK1vfPIubhX7zDU/u4kNs9787LyF/Ux4lUkx0c3
NXOfXYqBiNRCtMStoYe4EWOyJ+3gpgJsZYpNGVOVt9GY41dT8Yka6FsAQXaMX5c7mq8cqh49oVA1
DQJ0dnC0xw+pLldSiXO8DNKV8n/ImCfCbyXPL3L8AMfQ9rnQWP+518OqsTDJsnH9NhY64ANnbrkO
eHsHPzXDBZx7TnMdEQKslNbMKkR+Tma27iUo0KxZ0hQiswDnc7a+aIaZQuhIKV8JoOQq42wG3taq
Ar9UP0/rFIEu5DUjrbT4bB/l2VWT7ZHGJRlWP1MKrC8AaK+6L3Qkd3u54AznXbsix5qDi9wMh/0K
cq9QlR65BBTcwndSa640LJ5vSd8UWpKBs77yfLSkx894t+XoXzQvb6eHXKF1hUPIrJ2rmDu7Z1Nn
9XDfJX/BM16H+0VEpojFAr2Ow+R1yR4ivuGKoS6DMnS398k5Si3cPesqis3tcwIzzCAOv6KVfqTZ
JgDv/M7tB7n/6jN57uwIZKerQg5kJ4fSgeEC1rFEc/5mCma2eAQyaHGdgpfRpc6+YkbnSZcCj11/
A0z436dq4AM7Ou+DYp9hwkII8zg0CR/ifvvNlv2judp10+ubUH4rMKSLgQK9dHcVMscRmWJep9QC
NpUtw0+Nx7SHP8CLLQ0J4LOPz+5KJ31iF8Puns7Ji0zVk8LrA6Pg//N5CmMGPW/NZ/wlkD2vKPd1
vyPX+GgzGWMiaun+6k0API6FZ+R/blWwS8Bzpb8p7iGM5AoJmWrRF9fm4VTdp7Q6sPNfDSBM42NI
5kPp4P5tqI63N+yXt6ZDfruCjyZPl8snrGTwgP4QYizS7r7XUKcJ8j7urtdh5dv+Df4H3HI5A829
82j0nA57McOFTaYTQ+PFqqTBirLl/n9X+sRh5X76F49+AArsc+9tHBJ/vbmvGoh/6n0BCd3SSAch
XbBQURdREPwOoiW54wHAvTJ8ZSSWy7D1dba0A/+9fd427ppPiuMhupZBNWGPtvytoKkoDsF7+tpM
qaAmZ2tVa5i2TV3WCks5OsbCe/LQgCMIbv7VFpl7NC3IT7Z/UDkYlNVqSTaveqCFw5d9TiIlZsr7
AkeAq9CGJfpNxZPhs2uHW1Wk8Wh/y4aUhS0uDwo3ZdJD4zLJY3QT/fqlD9NI6cV68dFumOyxT2e+
L5UZOof+diC44+VfdrYSV64KKtxhSvsvot2KkX24ZqV+EDmj8qa1kSNfTsFCBqUCRIamTNl5eOrG
CuiOIwXP32rZGYXLrjywTHXdE9WcLadqmxtiWYAXtC2+hsuS+gqqoYiNdRQsh/WlRsL7sN+GpY4H
3mkm+UVyUWsWKqsGZImVtmxFlxZHU90e9Q/yu4NBv6zmoN+BGXdGr+hp+Gyx9QdaeqGGwuEQ0/77
lL4vIORANd2/GHXzau4W0iX3Vi2Z/9Q8PM6B1ubvYST3GF2xRRxZAI0Xxvjb2gxzODUBg0k6Ubr5
fydAAC3ABD/a6M8XhkDPG6iIhSs/KyUc6zIAUqvyXHUb/slFpxtqksyZv1livpaCGYboyY+Y4Kbn
smIQJaPY++NvS9CeF7CX+oieI/c9HUPmfz/xk3HpjAjRvcTLNkgupo22GDOyevYPJ2EVTp/hRPka
fdPvjKY3YtcpikQp4Slj4uHpMArjfFYq/JOPDLUID8iwZKK1KFZfVN/+6bINnc8mc+oyHfLWvxkq
caoGbbcsVswy6o1jDXmmzLPcNh88t8qgLSkwILHTkCPVG+BbOtIzUDdxBxe9peaF9zk+u/WsNg9U
+ixwUCiYXkd6RBppSEXfBSafOvO3renKm/pI5ITtrnY9yKogiZf5Uo/JHQ84zI6sSYWXGpJno5xK
rHr+I8IrLPxymMrNZQGiB4JuTHATC+XjBcATOS3pJ++JWHbrh9yzOgUAxGknzcmyVgNmKm6GcQZk
scUT66y5TdJfU67KjTofHQjep3/MsAjVtj4Q/1RaVLFxXuhRIgenhEYvdfJq7pf2cV2E2RVm/6gZ
NmKt57TPotsLYe3uNtcF9Hryb1nMEiXS6Q8kd9VwoZFnBsgqHQhTRpjYJTCNUbyH0gAq3VkmiHXX
mjDrASlc4p2Ol8waU2KQbwSIJoQIezMh3rDP+E7eEZ+ZWKLQtKUorvh4W1ITqaMOTOH3LClI6HT5
9nFEqg4nu+nu/KUJFBbdvGS4BPmlBx/mIORS9PV4JgQmIN8nMMzhoyZW0JTdnexBUyntsmdjDyVY
OLZGFveVlPbLaEAEGZcPPofUdD7ODvnC29JJ2HFI+XyFDo0TsKQCS4eiVlWh+EpGILuCv2l4xjyT
5JosymdwWH4xp91g7zDDSRTPp5MJHlHW2oXEaThqvmNsyN/BnTaRZ6e5EUThjpSO85+ZXYR5eh+T
8AxWiZoIfO5F/LqfYOBuV+Wnxec38Q5zcBYfK/9tf+EJDv1TzmYaWLIXanGTJp7/zVN3FEjrKqJ+
9AcmOqGGqWuifzk9Avw62JPxor5jIGiMi+ksBU3ame9MkmEI0uovHumCoisTSZ7LuM9H/gJb/4UP
hCevIlEte/XCqsmAzIs9r6JNP4BMWXc0c2QOMIpJZymI52hpZtyc7csa6lugyNd8Qv4U0Gf3Dttt
gCpMKQzsDG+MJBpsVmFTLOCpD4KEM+0xqr57WGoy3bHaG+3GTGSMtKbDEkcJybnu3VwS2CIw6rYl
DPGZUeX0p6fDqixshr4aqXRdz1hblUvuqpoFQrZilBeNKDXCBXUAbbnIIf792hdv28jBaNEVu4nd
nAwLtMxpq/cquK/j5UEmEuuC55UCQLmAuFBFbIGuGndFEFMdRfrvyIKxi+ouRWR3vuIZFC1cX70l
NzUB9mouk8L4EUbG7L8D8F++DGbn94eXe25AbWxsnrSxhXqmH4kLUZ14tmrsv01oJ/klImJhwj6R
J4txYTLnXKR69FNL3N1HJ8oMg+Pmvg5T+RLh0MM1Wm3rADPnvEMkC6ev7iuUdnChAZaM4igYpflz
9lKMbmBsXzOF55IqwPLa3YVbUYhlYm4cA8oKN7gRgyFhC5g2pcOYE/1AmwMaZOnGIYDXzKaghtnS
em70nbFgWyvrIfADv/esowlN0m0MTEZrkrW/yVLv68GmZHZngmN3FhZBJY1rGwd/uRoig2gbJ3yN
+0A0nQ5jCoWKK9XLcViP+qLfVK1Y67xL03/7LfVMI46afOVkpf5O9Exs1M5ENicKTFa6EF8vEqc5
aaD9UvCAudL9myPvso9f+ZYwTQArAaIzwS47oxjjZE4iVm8LgiAAYwd8+2TU8crnZW1cMm/QLIv5
sJkroRNdRJJzfR2NdDER54TuVmhCfN+pRnSczozSG42HTQTPjKWbLetaBE88/hWrmtQByK8KUONI
aYSMT6M5WgoqGoiLfMjgcw+eaDj8yQkGzwmU+cihh69grycfugbae0KKVUE7Xvp28GFIsN8HL9/O
ZvankksSbkgpGMLcLCa0I+OkyqGKOJYK4PLeheS2jnmUi0b/dLF8mpBLziou+UGCLDtLa4ufC3Z7
iISYXYKYdx7NHhy3EkbgQFEn5JweVRC8e+FlxyraYKH8bB5czL66marIIIaXb/iaPinTAs1HLueN
s0WJtpbUzxl/Zh50pOoTMSWbpJAj2WeaLILtIoXnS0735JEcQXtmv/UPH3wV5uAkze0njMTyGPW1
6NYcoEb9Xz9OjcXjZa7yKwEjQPkFK26Y3Tq+Erv6O+oLmeMreLi8KWYH4N0aqE+44iX/xZ8PYMH3
cKR8OuuTWnAFBLMPZiWU4e/YbRP4pKpUcVUoBjdlG6PdbTZ+slXmfGVRbQsvb115S0hpKjw3N1YR
izJDzMOWXUiitcL/qaQsBp0r5ACCYCAlz4O6IKDKhtnVCdNZyIu87/caLDD4QrAsRUs0LjN0cAwE
6OYk3oYnJpBSwA3FnnalsvieBkSqpkilORY8qqkZY6u7vzryCWIN75SPwXdiYZldrihEli6Rx09C
cXjmg80z1BDs4JU8C2pIhHfHKiu8YaxWoh98BxgvGfYDBgw6No495z4whik9BWKynBScsaE3gETP
27LtD73ExMgfTCeOQNULbz6aKrScGOucTWu6VcZsw9a8mWn8Dzt0rZnFY8hufiHPiWBTSSOT2HBP
o2zpHefuxQLRvB5LiOHVABwpExkLpGZ01GxYFmyaURv1t0EXogPLN13aTdDkacU/ir9QEJm7bOVF
xebpTutxNaFNQ8PcyyD7FrVrFWxLlut9RipipMnVSHqHNa22StEp1uSwJjn6k6Rkikyc9YUJxZMx
VC6xpS/cbdLBYxMre2DEwLVM3iIFI6ruE+XXjXk9nfc2PzD+8+91AS4nuJdm56uJo86zbsBme23l
7s8A4jJSxv9jOk9QtNr8cVBt+CHuaU2dwcIlsDlFwHQM7mDwB7sy3YCeMyDrMVRPd7VhGExq/5Ut
EIPjbHYiKF7ng+a1fGVBC20KpIgocp1h1Gp//ap8ESp1OV84mVoazDSieNV/1PGm7ax5fEhUEMBy
zWmLvojAixK+beaH/JDhzFKc7x903aMDj9xj23AXS8xSTQmtGviJsXAxGCZggdMziVy9OQ7Ely0f
PcVGyOgVe3Y+k+E+Y5/Zu9Q/b+ulQ8GFhZYtKUqxNyBShwqR9mNoycuN/Gqqwky0mx4WdpYAT+EL
4aCRC7rODZ3QnC95cSPyN9wBygDNo2Ljrcdi8omIw8RMD+6LphmULIGmlCelmf/QUm7SHgqHJHFa
OUUACn1OstVBkd0jH67soKUFB86s3MTQgyeMQFbkrZlo8aKnDoVh5tqGfHbmTgNx3NCM5QTFnHYY
VDz4F6H0zjnGBrPftFiEfP9wMrlJjmTcF7xUE2A3wGBn0U1ZfEAmb7UsqpYudKszMx3KbHwjLdfh
sebkG56DIIQL6NMQTkXHUbnJu6PHPIMTobkcayOfyP/3faCxdO+n8V19MQzGfUGoIW4FTM0o3if9
bccTN1g0qOhGn/+ep1otq4WJGztw6ZorQ/iT/Gxd0fvFxFIThtcaJyUJUY/78DkcJ03SdN9mt1G/
X0cSSJxJqsENX4JWZV3VnBve7PvlhYk6fQBG/au36H8swsMQIxnRoOBrmf+F+oz6Ts0CPV9YkbRe
MtSWZejau/X1n4WlDrlZ8JAsMlb1VNOiaQEs+Ngq6QJBVVZaGRpAfbD2dJ3G0wtEMqxRhb4v/yzC
VwveKExsZZjHOtCmM2Zo3UPalG7UMNG8HWYWGytgb/Q3JOZ6P5inAwJjkz0jUlTq6DhTIJP6+CQc
DmDillJTsnuDcYq56xS+3MeSTLHbRt6HPurvnjpGLQj6p8B3lHuX/XA2BypaxQ5Oqc6ODS0GBeEZ
rdifXmiv53iXVHmug4Kljf1hNW9huSQw70ggsOyXHZSZLBqmoZQh5xL9+qiGnc9uAaP6uDgkVKEF
XRkSC+ng+nPMnj+/dpxltGzSlG6pCqZwX30GLoYR5bD47kd1sQiws/Sy3NfXZdMxM7k4OZuRHXNg
FsTGXZxbXyCC39x9kzSxzPfFMSO+XSlYUKK/FZKdH+/rk5dvj00UvAd49PErEKknp0RMJ8NoI/OB
vbmI/QOTmgg1I4tAEThuK5xMPwjQYvuJjYOsNJkC7ZEiJ+sy9QpfPU/Uqjgb99XxhhkLNGyV5pHY
uQWcLY0a2+aU0JQvSKaFtQ92HqxFKNxaY1oNq880I6DWn9A62wuBltJPl9lWFgVAE9gUDGJfWHhP
//8hw7auXHzWLhhdA/XuLt6DE53aT9bL2gVTAE/Hi0ICjZq4NxQMJ0Lqp56B8C6WR12uMxbnt1PS
VvNFa8frzqWImHahpkInNAXcgAVz1BkY/U8HMjl2PsNw065KR/Y5JW/nD/hWKG8Ey9LebFv1cP+c
CtlBdo8ZQez1qJPi6LrAY0LQHI5bBmAhD864Au6QMENBzIiiyd9IjQlLfllbJGSzp7XQInU4rvRj
5If8T0CSCw9CcybGSfNqGH4lg652jcFQtO2GTp5uSBUNVzChtqTZQKTIKuq2iE5bU2RukluSpsKd
/nBtF0hRy32grvXFO8zjkRiplAuuQhrPru4TAc57Eki+a73p8cVsMXpRfwPb8lk1i3x1Gy8FVLp+
Ny7EM9SXJ+1aZmOrZdNWI2yDBRBChOSNmaoEbD0H3l/9G1xx4iqY4tPSMMKMAI/7x1HgK7tAnWOB
sC1ty0vn8bJbPDnyg/KmoQUWH52hLvqxiSM3cSRaBIA/1dOukX0z8Sw6jxo5m59ZxpEm/Ofs2GQE
H1WB/7vVPvNr7FuK8Ae7CLTMtYu9Soz6eLc4FdR0x9SqKMWf+pPMbHZkvxaG6LRPlH8RK72kHPI3
aTouI2gwnZqDr6zXnqxlOJ3n0RVBMbYb9CF4FjJpq9wopf9yv1IlF1K5V2vS+SuI6zss+OvFnY/A
ks/RZrv/bufoghtkk7eGDaeNT/LUmNCePJxzjvPXKLeLcVG/6a9jnYJT/YSEEHxd0TTNlQCjBOsU
e39GNkx1lNsk6QIAoROmIh0oNVDU4l8jCjThNBrh/IOPVcuqcQNhbXYqYBqYbc5+J8tn3MOhvz5y
Ygw3A7Nhqk6mYSATeMcquBfZ/4Vj+2WPh6E0O7cy8+jH+Mn9TgLYT8BoK/eKLNSI1yU6Syslqqd+
lLpaqXsLh2CoT6pZLHOGGFb2Z+LgDMfwV+MmrZkLpaLwUa2djO57tUfm8lvWEW1pF4pKTMN3/eV5
kW3XfzApVQMXO3JVxO7QzOhqSHX+GL80yMaPmhQ1SaynomQEyCD8fiYvYjd5pbcMfz+erQiJHQmI
19lXGO8eTWVu3giIruw/f+IH+GAQi4Gf+4SBZq8hWbS47KyW+EuHJ8uL8F96iqqU2h2sGIve7UzZ
LukeKgUsag0Tes0x7Zpj3XSWZYVEJriUdaAThski3WV8B6TPlKjXGHmeV306fmGlQi3AG76idqFA
jwRr/xo9hRvtfo5WarcJKe/hsgm/Te1rytuNemzOyTLojTFh0G6J5Q/WIQFGfHEJApGuCwiU1HFL
is1e4Kl2by6a+uUwfTpWJFPOWzxEWXRbudsjKswjcsrHUFQEYffChP095pFt6wZZEGX/ItNr7iF2
e9QTO/+ogl980Ig4VGedzwdN5LE5nRuNGKrC7D1cxbHOJ+0d3Ed9WBHzl1O5sYioInJgVXjmqUFB
TYmeQTWmlOroHth/SLVpC49iSNGjsiOOYYaSaUC1s5z5Bdr+Z9arpFO9m2GIqS1B07j01cxN4J6Y
SbQ3AwFr1LHYdblBJkDRPa68UDy4N7D09mbcfPJ/pWVvy1M6zpYxBS5kkjBu66THn83Kf7+Pgz2F
NNIpwrgfOaM7ko9maAAtF2OQ6to0LxzUPPNJc/HkVjT5fMhtlr7O15mlovgRMJKrUUYd/jEgpbb3
skUCgXJ9d6IDSokEg5sXwOd6hm6iYN5SjNH3lSaQAFexV0Ws21pc1aKB1O2Y+8llAKtQeZtkO9Ib
2vU3x1o72bcHK5wFNaTo2QK6PLYuRiC2lzcHw4NxiQKIVRy3saMeqjJufh12Ng3jSMfas0E7cRPn
NWPDW8tH1btczQ4kc2sd6m0EeF/8iDhYZMCgiHwKUeGsB8g8eYvd64BRvAUqUfLVazqgpYT+Iru4
eKXl4WuKnT/bLFBm1W/+UyytbHxVIJ6nNoxVpWMrUrqrj9sq5xQ16TzWTZhfqDXjQ2cm9GuRlj5q
MHZHbFp0ZbgPVs8SrgVlbRcq3BXcoJ/YiNZHrcNDh6juLpqR73SIPfeAel6HSkgL2nOGdZz3z3RD
6+YXtmQ8tJZd+dblnp47vWsCHX1hEjqXgpxvBocosgTyxaV4ROjeV4jh6PQCXun8z0b9am9EaII8
nTw5w2QdKQfdv06rfzbu97W+GGO6/RB/f6WJZh3ZkWUouTkQkWZ2TOtmtbluJM+uVt2pjrXbqcrq
JOngSgKjwWxud/rcsprDA08v2H/nrococBZtpMzaeBlNJZUpOthMjK4p7AvkOmK28IJi+OjXSkZZ
TS7kKJn9t92/khr8ODOQ0p6vEMFxlCDG11cY9eTE2MGnvZRWxQ3IHbzq/9j6RJGP5cWM7/09PiDV
U811cZzR+fdx3M92gPnVdvFXbtW4Yr767uJBx+UL9tB0PJudXCDOwyoEMQrQtoollMyszluaDol0
3VdNsv01D0+XNCe2EsrWtGwjDJF+kP9J3yceFFQPhsmYdhnIkgX5ruZ64F5OB9PjAL2YM6giEbE6
9xa14mZL89XpFYhSNobhI+j/SO3eGqj94rOsj2LcoGHCNfoOMfJrGuSUV/zJo2HqZSZD2iVFGclV
PfLksKabNr1Y7/J71PwrpW2kYzdjbpaBVqng2BPn1AQmzvXYy08PqV3t2qpDTgzteEQ8K3NUO2QF
KA/L8f/kOFTuEeuk1BdAqYuRhYwVsP3K4fh/vyLPusmnkLxG6eLbCw+33oh2EVUlTnPOQaXJbhtt
UPwzUz1tGkT4XIEyqDilqlRCuEysEAdHDP4+EAPIzYoIXNhYim/oVke1Tz1wQSqBWKdxAd50MpFI
397wmlctnJ/HmWBIe+Jem0Jw3bPfu5Ck/EoVArT6CzKmc8GSqMp2sK1fgH9e0bTZci/HPIKBSyWY
wFLRRmm/W0EBRGHQ1Q0Opa34y4gugmAvVPQ8JJQBd7uNPocefpNoHHa9lB4u2ZoWSvWYJkEuIK2F
cFTldCrHyYEatYwVHg44ZRR7B1q0m9lRCOEIF73uotBpNKEQIH4KwK8/QiRyx0QbrlqYbRYI4hnS
IjREqHjDJSe3tUpJSCU9fNM1lhcLaNYpwstYz086delpa9jGRvBxMaZCBTTGsBAvMHBwmFazq0GC
CmW6hMjw2lRRsXWCRBkcWWW3QCkmtA6HX/q2o7BG54ASY0MfYMbGG5b5hQze0CGc6W2TZNpwHYOl
8oXHbuo25S5JQDBouM+KkdcuOkCeNtZw7Ww0fcAx3qOD1yucJlQ4MAbrCV7RKDfaqyQW/DpWDiNP
MVlVoYtHeJgEpluZGYaOurXIhNXhnagJtqj/4657pwyez6UfZutuKV9WYNkeEvxiC55Nmp3P2SM/
hsTYcE8XRI5pfY5pb9sdVtzdbw83xzQbydgF18UsK45wlkb6AFqwGBh57bzBpP5ONDkjXTbeBqzQ
DibD8QpN5hpgfmWCkY/6frOk1tF3ZFRHgAzHh8r+Zuvjd1k8gpWukgJIVgIiLJQ4cPJn40ZFX8ei
OLrKH0ywoPNzrCzyKHjnppaFpeC+rJmrPi6o2XrGp02s5vlMlhaB8VRLLOwInWtNFdzdPr2rdIPC
JaWiWEnR2Up8uUISLYTd7wZLkg095lCoX7GlOylpILsjwIZmhYRgNLqL9x0hOFI/f361LfwGyZlG
2jIC24ywh/W4ohWqvKNZ0zFGW3B7i+cjMO+41bNNfW1b9xZPRaIEb3/KZB5ykA65jFBYYBWw5ZOq
TirXhuYGjEpX/mbJlXQtmIBHEYEtydj2GjB+EWUWkdmviU6JQPjdCwNlXoA2ay8JBw4HWFo7nfpI
8JkSDaWWCm2UB0yQMWgJei34oYw+UJgs3rRqvKCaML8yjxgRyZqoFdY7J6ErTwxSlKk8/70h285b
5yk7BnxW94g1OAemYCx2D+a2ZHhIBndIbaox6e9vPLDAXjt2JnmZu8HbizJfUULwaAz5bRqMNG4w
uLQvNrrR0JB0fn9W6Z3v67+9QMvdZyQ6k7KtcQ6+lyJbxM5eJ+5KsXmw/xlOPETnt+EV63/94whf
WsEki02OlEfs7BLBL2Pl5pVzzL8TBRAA+gmiGTlAp05Qi0v6PoXh8hTvRNGETPiuHcjSnaUUUP/Q
LHsc16OP0ccpMNIqlj2F+s+fF49fSvaH71x9c5/wW1WpMNmy4Xaqbrw1Rs1oAZSypYKTyHyU+uTM
Ux+gulISlkT/TJutSc3QOAbGP5fWzNI81UoRXZEBbdeNpDYbITZ/Fih20ytuNJVre0ah++tvP0e9
hwixvacuU5ScbnymUyXzdNo37Uf3/CL9KgFvHQHktUvnGu5/0hg7dU1FyP7jlPal6u5rpM7oNBEJ
zCwXZ26efm4sAWUSMA8l1hEsGcwS1a9RMQFMjLNBfsvG/02wmsztaDG1aIbUjFH0xXGaWvTx13kg
P78uIVf140gzV7I+HqVg3yxbghoGqmSi5aZsJwGHapk9eLiVlgODTcOTR3ziKwyuqyAbkkpZrdkX
IuLEm2YQAzt+V/wkcKgaTLyUCXfuVW4HkLczSVZO9nreGevqc/GEQBF8OAmAstNz6Mz5mh3wZ0xA
VP/Ue/6OLDQPeJXTDmtk4vj0qXxJl1h4/I4eINeiBy/TFp+fJpMgxP4uvKG7qE5rED1Qkq+1FgLN
QDvROcI/ecs95U6tLmxBJ6RPJuTHJcTjW/7giXwx4thyY21anrYukSu9F8PvfhhK/5HwHCEOaHAH
jQFkt2tD7CUe15YH55CbitoN8lZBQawwocZp0F+uOmeMSv3BpRsVcev0zwrvIi29cbxzFCRGBP4V
iaYBp9Yvqtf1A4h7s64zrXVqOvZ334Tfiw9VralkffgwFH2cmyzK9GA02PLS8YAltH3/B/lkBURV
zjOiDKR0yQLxcAtAHomcum/iX24hOdZlp6kP3rrhIgNt21LxweAgxHCZzLDHGIZgC4wgqw2SkrLm
XtoeGIjEuvJ+pxMEEjmGNmt/HGFnJIPlPSpXGOg3WF/VLNarp/AVVeAZCxRuGoiOQscZEaed9C1U
HQ2NY9uH11ogtCvpVcAVl5vzgxztdG/ivJNGSWfeKEWrkT6IhYzCnDhZgBoDjByE/WBPPkcGCo21
5o7pbiT5XyaacgLn1q7c1yXG6iRVbDBwMgrZn5C/BQv1gzAVSmKL/HqrYLjwOUcKa/ZSswFvyCNp
vVvWIJigPFT1fezmI5Yc+4OD3vFfyS3X1EgHiT8tHeKEyem60FCrUJh/s9AM5c4EBxp0rTOi7O23
lydrMfSN8mh6MN5HHGuLgLhOKfk+RD6UE5h/Z2QXGvhn1cWnSnme7VJD0fxNyZWDyS3IdMsf6ab6
NrExpMCrUYEhNPxnaWntV/vZHYATJrRMhIclYCiiMmRdX1rHkFIHEpwUaLgTv2GyyqJZzJPao8e6
5xcQkE//LW1nxGPkDfGH2plAf1QuqcRlv0ZW1QoI7wj/T6yzDC6CDlGmgUWkA2qXLp12KRHG0Vbo
XrfjmnoV3Znv2TAPv8cB8olZ3Ybjf+jUPGxhyPnBzzebOutQXOAWX2gTh03s5zVhmWeZ06oxF+dK
sMzJqYMnxNVJLi13xmKYO6R3k6bi5kdXRBtSlSkSdurKQ1zma40q3aoF0dd7r+ZnRdgwn89r/lHY
sS0hFCy/K2dmlo0A8anXICBFIC0S8n7imtL/8NCb/JydY0U3drHLO5MgGfpDgMJYNvl1UBmT910a
niHyNLpYy+tDh+B9QAUT1XSnGK4NcHFqeuiWROXxBlEKmtl3hyPzt1/LlJvpF6MMllPAPrxtkL7n
8NeiBfh8omAqEnaumZze5hulksq+juCiOxfwr+fo5IO1zkL9/OCriVDUghjU6yaHXz16dPxA4bOQ
pNbfAw2OJxv7U6eRPzjmjlVPVaGU4XG/M7g2QPeqaSMSMzmjYnlswBtocRroRYw9W9K7+q1l2k/c
uz70Ml2bqwkfsNqdAYxz6l7muWvyXasWFUW6etEwMRmr5T0Jsrfng1e5FZi3zwulOLrirmFs6q1d
af+tJq0CCbxgs9QmED0pLLzrvO9ICjT1e48km2ejZ2PBkFM3zEcYGrtpVMjOumGzKnYSU8TbTGaq
Ph5zxym5bHEgRaNp3eay/91hVHG8cJ6n/4S3tB+NfYyxS7Xxx2azCnFVaLsf0hlpBbEC2DM+wGDd
D22xZk8qia8wSCvJFCoaV0oDBTJ9cN8GkGbpLCaS0eX0uRv7EM+OOPGMsjFZuuFlxcYPhf6h/ZC2
iSQXtX8/AzCEKtZUM1eJj8Ze+V/VlLOLf8VS2b7HzMPF1n3vjCUed9tVdPK+ltRZ7d1Yibz1TLTk
F+LiInkiiCYQT0L2VfHfzVRxSp4NDvQ8n7Z3+GqQd3Xx2qn6IU7uDIWaxFgWziHxAbZBo+lvTtgQ
eivdiKIo56evPmuHtVkpoWouFm1SJFBLwNvGaXGF0umnjQmXE0QNknv9j/WrdnzkUtqIBh8LuLpp
7cp3xsC/oAz18WNpVXs9ZSsB3ULxRQBdZgmaSLfyG2cxSLCxUSlZ63K3w72/FW+1dBaupXr67NkX
eyLIeWT9WdKbzYretGm4ARg1wzlVMGSRFAumkOEdKp/DvG3+vLn9uM4N3dNWhRVvqeYe+/IqScW5
rXJ1mY1gOsP8Q14OZ7s2OgX6svSmMyeGCExn4gQLxwrokFAZ3lV1F9Nz0Y8lbbjClWSbmTjVXli8
ItcDxuJlDJpXpZdTPMdrvL4iUiI1XAFCY9kXlAYzAPP4NycagoYgUJ8uhxUXJ+hHbpYWILQYqpWv
5avSjDLCYzGHhOSRym2SYMHq7kDeRxCmB2sLGmeeG/D6S8kqKWK7PKbkv+V0J7IEO1hzDvzQ0CiJ
Cjr3aIqSy25YqaJvoIjIqwKemk2FOekhEK6cXSTRtL3rNw4R+IieiZyZ61Bu1V2hLGq6cGcLVxXl
J1idp6bhY1Fi6a17uoKg6h5W54CuJ0L+IT22AME9qPAkezuivfaNME+zEW8l33DQWzoDMM8NxqMw
XWWHGy/23NEGUm63uCEkl2RvE76g9MDWufCK62FqqTPqxPJ4NvxBTq009EPtMv4TSyeDP0ErhnFW
oBSh34l7nH4IQ7lHCyj0+9KjilzUup2lUgUn7bBOPZKgw+6c0zfBsMa98395RP7so3uby3KNmei+
5sZZzZFPCTxagI2h0iAkQ8Exh0Y+uUO9a+yRXIVuBRbECXP5C/HZPX02Ne5U0af3Aa2oPcfiH2V2
PWir0ggMuszlE7P67dqV6d3CtpIulaxDJCVqRNWFXOokVdadmSqQMLZkxDPB2V2/Ez93j8IKBN5F
FDjqaZpTDh7y6hRaOMfZv02ThWgq8hZbQSmF5svSQ2s8Zas1YiG64Rp5MGJQymMW8OUYwDRBncaS
UzsBqjOj5qzLE1X4N9ytYBoSYhToCWtsvgjoKYuSVo4zYNEh+e9tf0TNtByualjLhxO0CBnWRHom
n8xosJNd7kVopDg0Uc7THVAnpunNrsabU/88rCLKZHp1ziG9g/X37+Gfht0Adj1Y8ZI+C2WAALeF
2iCNA1pcEErX5k36NlaScArCE+IgDCGqLOLENCjjoIjzBHeWQzVhIOU0s5shgTdlKN0lyraXHiUh
MHTxIj2U2JvYNKzEhTdoqpCI8PESSsLXfbvCr//6UFfxwCVwJgdVg1nvKc6Z+YzF1y6UbtsPTor7
dUukB6wGSWQgyPe5CYFEzcSb27oddN7S19zy0LT0xi9WTaWfnTntjXQoi96SORMl8cH+RMmncRkA
36pANQDgs1SRFIh1V59GuxLtWpDCfVkRMHLs4K5LcQGTrBjmR+r4rS1UfOWpz8O8TOppiql0jJky
+5zrfRNPTlC7ML/AKsZZHDyQugm2DK6F++tcdE/e6A26/ROgQTP2mvOyVchc7UuAQgUTzBucRW1+
EIcuMJakxQ3Fps90riaS7+o0o5799NykD6+ogjtKnd7l5uIag/9CG8PUfNvcLX3YQVC24FHhEPme
odz6Fg9NyPyTNFmEZqWrQL9UWkdNYTWWTwpEZa5SsujxUFpLMK6AozIlEbVNdG+lVAbMp6FfAXSM
90/x3AlQbOnQRNG2v3zQP5Qof5hSHLTZ/GBRW6J2c118ZHaIPonuMTPEfA2YiFJMYIoZafXbolh1
L9vsCCVXmOr7q+BS3fsIkKwL7gdFDAX5R8UlYblNqIV9+j+cv9BAJADNF/vahY1CQ6+fqzYHTCOJ
SKqtJSeam5vRvbpvhkAdGi3wN4A6DdeWpagr0aU3aSC9Wb+oV9bicSatNXn783v+ONrqINuzniAK
evnv3XhhPFiD3pVjRts9IPynI21yGi/SJynYNuaZPvP2pptF8Jc2HxVTYebOFM6jyqCshXsj+chv
L0V7DgEAVgnWMupK++Qgm2KyAwTalnL20IXCe8HvBsLMq5BZ+pmHUfXWr7SiK1GZZUdtTDvWA7yM
jGpBFVktlw0WGXviZTE02MrL0LzYi8BiI7MnEGdCMtNC+KYz8RtEYO8RbVdy9WVyvv89mLmSv7Pq
GkjiGr/Z0UnhcAE45WvqLDhdDW/lwG3cISS8pAVMzSVVdakTIViEGc9liD1RtyxB2XH4CjkiYSkg
WIM2C+HDJ8yAgXduMg6NherZcErFNAZwF4vbtx+KiZ/1gYKLO4dBVl3WbIaPKtWC7VAgef2dgTyF
dQA06YXJ6dxAk6oZw80Nb1LtvpUnrhUu5P3tAlk/4oqhlGJ0rMuKO3O027ptN2uRqf8VnPS2Ai44
Rm1zy9o3kzD1L30gWrpYC+QL8kdB3iXN2mNQPqVtX5BPPc5t2fzRKkWNggMJYnrnRz92pYeVKPpZ
aemjDydUcO1oBuj7lLln4PIefzycaJbQd6klRVxu9FiIK/TQJ5tHmEI3DtKAFAnBArZkElRh6fYz
NG9EGjSwPCGsNBZE3mGeOY9J9B4roTFEKwfB2PjvDvFRO9/r+TLtK1ncRVBcXBiM7S9d9AxmPwwV
THyu2JqoybKVHXkIeTEg9OGgjEDbekg2iJ5EFJPjLkOjLzTz9wbysZQV5eLRhaADOHqtKKPnrICl
E9FwHPl9vTv0lRk72FcexlYFWJ45zggfwNcwkJleRLcELep8tsSDvVMH6Y6XuhSLPDQBr+nMlL91
KHLfGt6+1LXP/ynLMiSvzhEErQJxxqlnkRggs2phXKae1WdUgT7x8Kh53CqbqGDX+xvuYYWv6ldM
EB456YZ2FOKEKe5/8szPtclVPZJhf5OO5hd3ekNVS+aBLaNPjoZeCL/cpZI+JwAwKZc354kmJV/3
SdptMrpQ864HxAWwtlnDUyZxuQkvDcRrkMs+cHCZeEvH4RxkOYhvOBtAVlhBJjM9aTQW9v+Tang7
AmWMe02ZqRrX/HdzVyQ2tz5pNWfAYCoYi1CzlNFoznfVivRnJO8ouCOvn141xKJbRBOxfAUp/aX5
ga7TcjJczpFXdCk+T+D6urUTjxxmcE7yu94VQWc5+mr4gz2pFdRoiygheYDD8pFwmbYuhAI9uCnZ
JZsUZ37Czc4VtyjjfWhscZ2iyPXYpLEmqZpnVnnUXpfDIvg9wOP+7ytAOLPe1AbwQUz0LRJJ0nzT
wV1dxV0vmbdaE+ucaRwU1r+ULGrmG7ziHCI5vywJ2vFEZ+3LH1ngugwWoCHLurnIxUPw7RTSEkqO
yhXycAZh0x9SRfaDgJYYStGcnInmz9t0H8+V8dOvdL3SHGGs/t0MxxRktMD92nFG3t9/H8bNELDW
jPLDPLrgDMIe0ObfRKUte4pURfYfIbPOuD9Zei8A2aUbsj/mO57mQ5eXmAeMVOnCaDjSOPU4m2ro
ZV4VKjCRyOfeqvNw41FjbLaQgSxAFbffWXpSLOkgucweAsWKGFBcKMX5Fg3V+VUwlsviIxgkEXw4
eG4FOmIOS7yM5lqGdHQl2qkWQJ1Sc/Qlgw0ht9RbbFgZI0CsDSjnWnT/Oehs25xHjXMQ3aZtyFKR
jF/gMi7u5yKJfE0JHZ9x04fc19XIBqEF1ldo26BwqQ8/rE2KJ3aBhmpmjUvSAPRM81Bhssa5CZm3
hwLL1a5lQsjzlYPGpEdsPYrWa7UXJEracBixzNV8V1IFI0SEFePW/g1DvaP7PtR5Pys47+ldSd2z
sCx+WW4xFCv3tSxJcYbjNBI5bITfdgdo5WkUkB1fKnfYv40cFHGOucvwjuKOw0y0YNnUrQPm/Hr5
DppED99TUTkB1oUB012b2H35b4mw2305e9pw+gLcIuiqWZr5D7KXGNvdVsAPuqWFErvXXBdZkUV5
fb9QEHVkD1C4Juk267MRbfFbah4rsRChA/AUOOuoHEdBFIp22D+NjSMeGUFUB9ej7qam/5W0BQqo
HKVV1izycJPbFrK6zaZ8k5+ZvUqKf6UxgwZzHoRNEIj5fJW5F2z2KUGw5BjSzRy1HYVtDZ+HDTGT
Lvp1x565jkvOaWSzUvhPYpNFVLQld+OgV2yJ3HRDudPcBBst4bYBw1QlB/LYQZc4VdkdOsAAhEoV
wrmxd7gTBpN1+PAJWtY5ur1cLhsk4iqr44JxcFPMD0/AOZ2amFZuf1dF3GlInIB/7S172/XJ2Anq
YVRh6kSg2yciz6ghauo79eksAJUv0evzW9g3GfNGFTpSwyak69K0QbX5jNIssoXfp7X+kpWlrxhy
M5LMU6Mo5it2Diqeh/MgxrlHamVOUBoLUjPfIbUuNvqrOsJDk/9SHZhC9Zox4aMSlz1rfWhPQ7aR
O4Y6vSbMYqAIvnN9BCR83FQMVk/Fa+RWS6/i7OZoB94wdGSUUviVRZ4nho4hppog3+f2n5J/Vh3G
a8lYBOH+tVe5itt+HK6Kx4YS6KZN/aH8bDCosbblDdjkyawp2z7SiJ8Ah8XqdyAxX9hDOIJGxqkH
lCpIPQSmEekhpaQwVqdPzYbMAUDaN8BRZoKH0ZDPBEKOExKmZ0UwoFqP+4rIZR1jZifRRpVdUPD3
dE8UPSKwZ8iagmnFSMbeL4otGtAIyjohbpmIsUwt4mAuKeEDWfb7Zj2hIX8M+3/7ZL3uVdVgPWtl
mpGjfR5EgkVI+gHlGPLLsfVdcuNbqbrpoobOOE6BohBJVrVuPBoPVNyA64hVtrGVyE1hSZWnLh9m
Dz3fF3a+Y+EHk+4ZwSdFiIXc8HNJPK5klCApbqHW2X945I3KMdt2hmUgz5Cef7YwO7UO/nYg/nl9
ZbZXi+SQxmgb4Dg0dkPDQeT87B2fWTM0pUqsEOVUsAe65JjufBG+lbd8Rb+gIHsZ19wp1rZ2hlpk
JykpEoFv1XFAEi7kJzvpaynLEOUosgQHpWpYpww2zbWGKP+kKiqMpLGuHXYf6Xq4ZxnUvzrC1xj0
vaPQTmJC86ehIRtyQrcSzLnz7REyoUKxJwykgCTNIsi5qlmIn8V2ABvNw/cu5IRWChmtRTsDrbrf
vRhBqp6cMf2z34/Ai62CsCaHZye8pVCmNS1d2tPIVL4L6y0B4lArdYtq+mBfBBX/qCa85SpYEmGi
2RfZt4Z3PtTqxEX2I/xg9IlgJ1/ww5a6P1DoQNk3jjZXIz5UGMYPdcQnwDyGNkjg3OAAPMdTIP0X
LYGJSDV4FDb/CF6q0+FnavFTFzR3S1lxKydBeFu/ysSZpUCauKBJP92qgIInhsP782Lw7yIQkdwD
1tRZT1l1sD4q8PvzXgDSLIN5qGZ+/sTHaQuh/gsfGUZpgWhHUf/N7csiL9G08ZUhb4Czv0zjEuRL
d9tcDtKsNAy4Tr0bmdYEMgzn6HDWa1PPmoFlxjxi0/W3Vb1K8bmzOKSS4txFkPys3wu8JePO4gvg
eQd1Oj0O+l1ucW+yHa40qraqB90ChsVT6whxLuYG8LSwDT/4UHscwSyREN7cAcjJspjwZ/35MDDB
C1hTrsm4pLOTlXu6gezN8R6g0gB3PpMbqnvkS7oRdU1f3QdrBJg+z8aY/r83yJrmocpZNzHywbZQ
YKC8OZV3++FcINS2GpuGJxKDH08mDFNsIrWLpCevqUdrVigX4NgmIWVa/0JCvRTBx07r5IOLjcN2
HeJWyDGVBCmD6qOqieBusvTCfloa7f6XGnwp6zAgoSLtkr8Bg6dLZQ49/houCPIFAEFEmrEapqlk
UH+X15jNP0vIkv94BHO5C7kblP49P6W4KKNwH/7wUKa/7hvvFigXG89iUVxjugIe55UT/0BwzdGe
di2l6RzawUIkWaYCXHvXDg998egQ9DusXwMNVk0wd5z7DbuszhpWI4nnH3cfoUe1c2TrujNE5/AL
af0wz2dcHzAg64mckaYNE8Kb9+Z5w+NaOexEXpsvSo8+DDpHAIel/VE3DOj7IcSsbdRS2TNf16Fa
K9GDFhZ5JTfpWpaYTd/qUIw18LW0iyeoROFgLORqCEAogfxEcQtxrouXLIsdexFFImee7pVIZAQ2
k7aN7nheF7HNqjTnDAls8f6VuknUVjXYEdz+fKod+mBleuzr48nw1ofuMSMlSj86uU+waYrKRo3D
9Ur/UKSKOtlZU7+yx21e6CkZYa2SPJBlXOerrBWI224mZylw6omaZki8JCzH8RNkJO7VaXUJgXvQ
qWSfxRsTDupuDNFxHmRVuTQsYEpgFrEUVl9gWiFBGcV03dVHSbBdk9+I+QlXHMa51HsX8O6dH7HV
tQT8lR68AFbPkun1LCh/HcFfPwJkNTtW3zLS2QqGF9dgJ12PbALB9KdjF5kiYnUQcAs2a/ClWSU6
s2EDpmwjeXEFJb/sSI2rK681O/q7aLBGXXBCfgsJ9gU8cieBZUvduwCw7aVOqKkLRmKbto+IBWlZ
N5rz3LYOWMc9ETjaGtYrIqWA60puCbiJ6234TiNB75K0KDwyloQwHFxrxgjE8WBziESYbwPt1GC0
J/4nv6mWZJA+mYbEcWQpJrmlNgZU1UvPU+GvaUSuNacWwZjukRne4d0NvpCGVkHhRWHMVG6oF98k
zMyfirf6s4dOLBr6LANEKnEbjB84p5FgwzA2p62kOXDSCw3CuZUIAeMt+9SzSSa/EPAz5klorMaV
M2Cejd0fWyxQ/YjQZrqsjST6JDltAzHyUE6E20h3yoOYktm/Q2M31yeHlUi7+XS3xyqI+ieMvaRX
LFomtbZY6R1MwcjjKbpO7pYq4owVBdAspgUL2hE34Ti2Em5+eCEPf1NHJLFWm6KgP3i6eamMz1gh
V0KfiLZAU8cRTWUKL9VRzBvvVmp7Nu5qURI8NC1qY1a+UHacHGyWp7QHXfqvJB8AKY6Yr35wEDE3
3wSmruTIzo3yRlw2As60OLRH56+2n9bWx/v8OAlWmTcRrXJsi4pUNWZyX+8dWKXUMI1ejXOuEOeG
azhR4smAuHuoxQEot2drX0AFE4tzOKDQgU5AXlkDYxv8d0l/bVKgJ6sJTt/jFeSmTabLIhJ1FvRE
bugxC7bSt+lmH5Mbm9Rw6i03LvWz8KgYeJRNcN1pBiUDEcyIP5PHB/EcDP8/isPe6L6YvSYbx4Vz
Z45dFgv79vMjry28TdZuf91dLWukDnPCY/h4Q6zRSZ3X1xL1By/XyGHWcpf/vhNcdlM6r8iAqSSD
0WwljIpcULaCVWSX+CSInr1YpnRpWWU2dbXtNoLS6BArTSdbxSsJZMPW+YZZmIdyDhl5Wp0a3vSG
0r7D7xcMNffy18NYqxLvb2z6BmgCs7+YBqEU6mbi8MGeg4QsaS+ON9h0bjtNtOsEUmr2Ar8U7/T0
YBgZEBcXom2J73zZ1CggM92907sazN3qrrCdNwqw5t2qYMNaPT+Y2TImsaWOUfVw8AJpyxe+B80r
eh8FKfEhneGUd2oAL6QSqYIutPHEcBtztGDb7bcQ2FSn+RAQG8s8IUkgSrX5Il9IOEmQyZVedWSh
sR3jjK6GqcAR5C8khkYYMwxPU3RMxZWGJ/bFt2tg/QvwBV7tXMg3sM4+XRXAS5Jb7WJ3buCOAFwk
z8uLIaGh/gts59Jbb2izisscvRs/U6VHb3ai4fvz4r9KWGj/bC9exybn347TRLquKKGreCWbvI5u
5/m1nvuUC+TfSEuj3irQt7wwQUVdFcrTFogBcC6fc33UNckDMMY190wA8g7ZY/O+IfKRApzicun3
DcAseHwMD9wUhX51DR1jQBP0NxEfvrdHEeX76kpW/g1J+q/ZR+pFL+v8PukNzgPnllJVfRZj92/A
WuNEZiflNmGP/DhtztoJl6pXflU9Aj+PTrhwZnon4JaQ3YJSH+s/63BvC+mvs929E1sOMEZX9vFZ
ynNwlww7aZGcDYXPS1lVhO3W1NPZaO29QdQ0xd+LwH0Bq+AhP6e3LEhrhoKUGYoUyXtir7zp5+h4
TyGZecZlnoF3hJTV6no/+5I1+pN1S0tkJCxSoRdYDBLkIQM40/DxIPJ1KKKeKcF51C4y63J3DD4I
Vxo1bq2a8tWmEgE3fsvk23om/2zqZXFHZ7RTykEnxn0NmzEsNXMxdGLRP9/b3BRjzjKrtaNoLmQr
7mC7rG0zilNdlCiiJHmV3qW/fQUhNCGXH/pFiFQPK2HhP4zAey7FaNvtNP9ZFh2CfesyENuY4Nie
fcY2JrTiDnhfmSgR+M64XIVIPVd1++JMaUQ/fcyAZpm77AO8BUC6TklFXz7+zvNxUZ8fFPNAJ/Aa
vTIlWKgNHJzcdfvDMcC/30AoA9rhAsoFPxBlTrQN7iwQtK3kmldvdcflsj9gCespVnFPLDp3ukmJ
3EKk5vrXpIcOzeGF//9Qib9/LMvB/pgsSPh4ioS69V62UpmVpUD64AcG4r3RMncImhbYUri9KoOa
jhpUVAtU12ck0sktYgLrs4lMByY1YRnhJasUm0mgrZpNic/xZRLBN1tHcB/FyzpxlzZzC4p8uvDR
68ZOVaR2ta+N1UfTUY4ginezLVhJMqC1sc4z8mVRHbbyf9Pnt90pkwd4xbQAW3B/I+Lsqomd09Ez
vH7RzC0V6D7fokFFVw9dlWPLpn5P5WMnkdjgHsS5o2TJ8nigFcXIfSTrD+x5+vlkdHGfXJZmczea
m5MmAP2slJvx41PiycYLkP33YWTDzDq/WJNbTViGK4t2sXcOODPnwy4rWdtvxYBO0IG8n1qk12g/
7n2zHJlffRbilqOpk+M9YFq2vVVNMb5YjGwrHFDVDJRYynT5MTypadrnlLQWK5F/+0lwtUNK/FEu
J38AhRdXM0oezn/n4Npb77b5E7WoRq4/IT7/BNIerCRxy/aOU3Y30JpeEeMWglWcDDLpNyF2tfio
ZXWpw23TsSDgf9ADRPPwDbWq2wyVrA44o89NsvIJ7M0Evn6p1UFetGp/PsgxjnIuM6Eu0a57Ozpn
F9wNTkkO5k4gZ3lndnFlsxCalffjnZSVljv83+9cbnyeDjQIltPpAvUWdLNo6s4cBkp36XWyt152
nr+Wzu50tgCB2UqlFBkndICpPzUPXbYSFcAkRFxa9UvmutvKBfWJCzxU6XUgeAxFYo0rNUtDKAER
3E4AxMAmF1C4d+xGRuC424Zft/L7cjZafGgkSeGANpu2gb2aF73UVd0QEa7xbMsVKMKtb8KcuAWO
cCHlLghgWoSq4q1MHXwAc7FS0lfWEIOKd8arDqJiYBD5+XmCYUlc8SYWKbMSjoi0P/d7pRdtQ09g
ndioqOxqIp5Xp/3R8Ebp/V7GLH97jSeMVHo434bhw2f+AXj2TIlRabhISB11NaimJDXlYtriMr4x
M1FB0xMud5amscfoxOVn57fmFdnMVqK5TDSGrYFMFaJI//eBQdv0NZxKVDyamd5zdvueIIyfxqNu
Lf/xsZen/kUOEe+9PdYAZrP3IRfhaTe73aCzTQRWQaR3WhgoXoFf9vqfRtiTt+TZ8IiGc6Pwlsp0
yu8Ac79rUjyMFh4cJSeavXFPdnvMt6JFtRpBLNYaWQG9TxDkEtlL9dpAXXl/lhuQ0WsyOoJGEXVS
uZuimgUEwsobSL/RTeDuWKpR5EwO6Ps06+2o7jfeBKWZ+b88l5vd46xaaRCo+mZcWZu36oDrB8j9
KCkQBAUn6GayDBetTN/6KpKTl/x3EybPF6P4VzsmAGZZKwz3+7+ksdeBxxRe87KQ4wOhcpZ0r5D0
khhF2DqX14MZn4RX+ZBFwUyZiSqbqD+D2CzzytSlO3AvXsuQGxGZs/45tC3QgM9AVLjaBvqJRQoT
Gtq/Iu5+AC/8/WsOG8bOwcVKw8HYjD0Tx6GHhUDR8xPvtHbErqH76YsjpZbVEBJs2ICBGyVqBxQE
cW2L7vQyFHO/Yfbi+O+AYjIWgx3xeFgh+S1fNzQmSUVTOy22JUyUkAAp4bpan2xVO+TkNTi4tGsY
/Ag5nEdGDEOj2f4Cz7FEzI4z2VIRs/9pWN9U53o8+uaPUYA73MbVmpyM+uKRSU3U1tAw0KCHyp2v
F5M+7pBpCTsUwY6f+KMjhbo0xwt9osq6UafZEui0vX4ZyveAaX33638BlinjvDcVta7RgM1E7y0Y
oGEr52P3lue+TI6/D+A1llXWbYhml+nOokNv4Xvgo2wgG2odJzyCH+vtg8JPaaBfY44MqxvpB9m4
YdkrrPOm2g9J6YW24r/nuYFGYGU99nWmehE0BKuQcXK6tu3KOaPqDG/fAIztEOBem4tC0J7omn1v
82Dx5iDfh2FOMeF55dOTrrrAwP2YlIPAhVVDeqSU3df+BugZlkOJuVl29TNzGvKqVzj4strW+7Md
qrUCl7zGU0lKiX+qdm0pk6m7+utNMlhrysSpiYRla8eM19zVSZG4xVArzvqvo5OUaiUILgijDiHF
CKW7hJcNsKuWv1wJIqeeaY/dELscw4mF3Iwu+93PY3QG28nxyV7bSeOte64vwku974rLYG4dQ/zy
f8j1Rtbr92XJPDwvaUCF7CHeNPPpxJ3x5qYAUpN681qxs8CkJdZt7z86CwJ/wplc993ryL+DypTT
a/LVZfguq10RjD137mGit/c5xsRQFFFOv/mmYJtMHxC3g5B/y1D9NP2LH9h+9Q3ipq7NqyGlhNCA
Wxzm+kHyVpZvGlXWujd9oGe0XzJyzNowB+/fY7+3TPxKrc+ktTU4ODOsVHANlJ+1+Vw/ryO8oS7/
89D+ltpaOnpbzsjXq+X9slN0XKwVq4tz9jvxRqJX0hg+zy54LtFURKqC2NTvR5MiSqUsl8YBo5rQ
IPn2au5SVVz3uI3Nk7bYxGtt5yRQgz+JWFRDkHCF52yO+lpOJYuhuzQAcDALuzzoYHloor7/1kbf
bScxS0qwT6ROUVGHF55Yyv4zfGBVH2MvH82gAUOgXhr3IGDVgpF83y0bQcbhntFAZRLqmgXyyTuf
a79LzDDk5cmLXFZ59r2HS9i8l5P8MAhk9UbPJtpGsiI2yUOuRtFAPsUz00CKeCqitw6G/S0D39ls
D/TOziPIjqBymUykzQhDuUPV9jKq7mTCif2DSz7sBY6i9Uhg+PXirtiFzq4QdGQTurnowRnkYaJd
rQOzPUqcinsGzigw1hlIpM7zy3fKh4qLFBU/mnwzZMtVOHFmF4T2hJNmehqq7jCQIUVkKKhRhlfn
HktL7qN+kGL/cTn6cRtgR2sRJdzfVCzKcSn5LW7AzgF3vhaN3XXk1+8m85qQPwFAj9EPmoxVb4R1
a6achXDmKblle+tHWxXGbQjckAX2YFSrqVLhyPNkPMvYlxafpIqqHsVrmvg1V35doBcBmvMBBTZF
EDK3a2l3zhTb0egULAMsB14wABFOh8gNR6HFhYCQTjqS9qt9GUlH0sPjAxZJVzUGZo5VD5qEW3Ab
lGS7gFBu2EziJYFj+p2zEYC22Shg7aD/br+VvNWhaKR5p9N7q9moAVVojVQyTeuMZt2P5Mrx0qqB
/h4CDDnZHAXPhH9p0GtHCkCMHzfBut+NE18StMMApN4u7SaG/OCnPx1a71pQX+l4LIiTPEJRg2PG
bOpKXd/QvYHllipo4+iTf8fBOWyB6JCxtIy1Wxlb8ynR09FPaBV6+gj2ETPM7uLO0VKK4je5SOCN
BEfohT2YYsbrnxKx9dSYgrWMCV7QIBKrRUzhCZXhfEuk3fUCjcHzASdRcAqFvTOub/QuYe20P5IX
CfrzaTYh3PBjnpzBTEZesvJtesreZ1v+EbUVbusQfRBEX+VbK0zWInJhAC9uGntbl0xzxej+HX1u
H+8acEOpdV8u2o0zzUS/BigW5imwVS3g7ZiL1U10zczrRdYHvj7H5FERmQMWaG8JQlLqCtGHFXme
4F1UzMsET2WYfbUEHcDPpZ0mn/7H54bNS/u8kvs2oSptP9dwnK40rvjHPJFJfpxWHX6LtKsdJHCC
Co9m/smYWO12PfU9DKRevPTL5+zcW9Mtybq7AQ46GwrGElb9lQbYZZpXFKXO9CQuv+rjFKLQ+kne
RyvtOvS1ymnScB3g/SFlswde01oY2v+GHgYoJNVvtitfbZ9kLOEm448b38XjeilkNxyh/xXDY/ao
Z51h6muACvQjbdRCB0BsqiFY1RKat/Qlpkc/d0Ky/UiTdP/Q0F8YJpIvPJ1tIKDvka4bcXoRL6mS
nRLUH3dKLKgnC4NTwZ2f8YBZ1GQ9z7S7HPfGP8tTPkmPBCkeYWgoD/9MSwKsiBUkczn3fYHs73Hp
vqDhFVP0eBvto+TR1che9oXyfPiTopgSsHTUcWFs3KysRl3LEpIbRtIoJGOlZ1xp3GP/HyuVTI5q
Qji06pMvb6yPZKWLRTi3ohDd6N5fUcH2uMSBoUqaRMAiBfytAs+UPnG1f7gOdsM131aNgje3TB7d
M08ITwMqEwXIXMg7Pk3C/k/D9GPzlOLFqjjl5y/Rj919+neLvnRSq6wVgM2NZ89kozg42btG7e7g
sni3VSLd/u6+LYPiIGjCrFrcCZ5hbjWG9iu7B3BDFIXtCcUTtW79+JI58Dq3xv/Isa7ttWlH7ZN1
nNXWFP3epm48UrO3fEJeuVoRZWL+j5NCb6/iPeXr0G4aS7rHQE/aWTyCIFLkJpiran6wNIlwWRDi
vZ8V4ie136CHKatpJ3WZ97GnCTIK4NeZEPkP2cEGZdJDBt+qYQCIGfNzVHaSyhsVulX7eg5p1lU9
7ICVhZyNlEBr+feE+7h+c3n6hDkcbR31dDA4sbP4tVw3qFhbHkuN7cSZ0cavyIMoHuklL9d0gRZ5
6ywftt0B/IqmAJ/10VxqnCWX6ZkgZepYUYv0ssM2WZydddpkqBVLk3uqW4Kw8qvjJUIYk36AA7bv
Yn+OCRAr4xkSu52GTcLtxortgNOgYLqB14mVI8BU7e4R/aPRqgWJtjt2X+RLevlcQy5ovDdMVZFc
3dWM4B/QhOsh77bRe2L+49ROyUQkLv0fAETkNnzswcwN63AbTz9gBmZTf6Ee54MwDKb9cCE+4GV3
PljnlY/uqhRSw2QqvK41r3zTduvmYzyfZKGNekl5YtCtvXjjqGAgqaEa+84Wstrl+7vUyO4LxLHD
N/IAlJBTvM7xYMLIfII0PGxhcLnOF1Cmwze/tVgiiXRyc4KlJw3Mj18K5sxBfIus+2ZhQ097LW3+
/r46KUSDw0w5jstDYl+IzgGfNJxK5w4LP3/wNyJz+PDP+a09maRn8apNacmhQSO4q1iIk9nCc7TJ
nntHzxyP2LQoRitvheiPkD/mZIM6Q+dGGCMWeWuZSvN6nDZRK/jlN8OE7zWG7SyOceWHxHdEIb56
AmmaqsLd6c6fyc6xRy150rABKsRz3HFmL5MPHpOyASFEb93zA5GLfeq+gDt0LuLz2czD+OLXR1MJ
5aJxV7tnEqlBB0uP2S2C8o2hJLS6HgXTcmo0md3H/yvRoplKAPwikC+hbis8y/itlPm4Zf6T4N/s
pxCGRslFrzMxFvi/qonwu/HX+AINmJk/DnZi/dyAz1FbajbHof5DGRb/nd5CCJo/tRaeOdJn9S86
r+7CEH8IKiTez+5njQb7X0Yt9Pdm8BRG/rQ7IYrAH+fzPfDJ0ZWNeafkSgUBipJb4yYvaPBh9e5F
rQ23Kbrz3LqqF0q7c1L5KLdqqwRrXqoKj/d2df7DTUveaUMn+FxXyrkElE/Ocy9W563g4YworZiW
m9p8Fz9/8x+15Ix7mvzkzHumlOsPwZOz7xiCo1iEzmQY00mocSm6ba4P3AUwqbpqcbTEVlS1DLTt
pVdXVES45ZQ59Kh9QuJywDo0d4htuJwxcpKq1MtlVgVPFlh61zw+Q0uJAatftLlIbr1GgFP13Qw/
JvOU2Xw/5hB/RNO28vx+Ji7x05ezILfAyTS5BWeyIuuAx6l/2xSDeA6S6ahFd8VLcFuTQ3qLHEqe
W5he81jUQAq081KBi9/79pCH5djfniZqfHc+dOzG5g2BmLzjiOuUDm+Q3YPUQAHXWvHi/H/FFkcW
l5jx6b8vDlPrm2NCG7CwoRy3t+zs8NWSwRRawoZG5czPVtFEse+58Ii3nleAw5Pa8YXqkZD4EGVZ
GbApCjHdiBred3SYGeenxd5cFLYI9EtIsuqhs+AWbb8iFhKEnmjxS9mg+6TZuC4kRZBSYmw6EcGL
SMWmulIvi6FRrZa7suOpv37wM+WZugVl5LJBq8+5MbmQXzTWY4d0Q2zN5hJ/Ue6cHrAsF7YYqZxX
IJfYyZcmoN77c4QkiAms9w79bvyK5lQAjdqW0RKMDPJpgAselLRaCCF/AXpZfRp+D2dBXHBYIkMg
1yfwQ7eIHN5xNSurliBq3pKHpXx4dzfC92Ae5lEJ6hePGMHIda71ZecNxcaAEpgd994sBioC1Wk0
EAKxhSK9S9YhDbBMndsC4YOAothLnwDp1nAEgHr4x/PF3KgX9JWhtYLs8rn1Wy6HY6NRSn4ABhaF
63AiYzuIw4ByQiBBywwR9X1ay+28Z6GqZH9YKUS72GeIdmXKPyuLZyKJiDtE7lZzqfKdTayJdNCQ
lwcJf457oY5SwT7JBgV2WXWc3qPJV3czEAswBeKp2ARewwmboWC84yCx7Fn+2AMSjiNGJuNqKOKD
jaPBGLpK8Co5YSU3i6k/onJnHV5kmKnVYeNJJgenOlavG3XgsNnOf3mONKqtDOGjP9HaxC/vmicX
i53NsafHaleIQOlh1N8m4ZvrIUwU8/dC7xUcaBJ2aGd4OgChfiS5NE2ONkInrknpWeZ1F+cLT8KZ
9Yet2g6H6vCPTFj9mulLwoqOaJ1d7kx9QL54s7UOjIftz6Y54Xdm9V3R/ur4pxOeraTnqHYZr+qr
RpPUB7qeppj/hY9CKVK2XrFq9MEbr05V9Mxrv8axodv//YbDjLGuw08CN+vJrdYENrj14Eh+4FhC
sKv4vvCxYO2TKEUoamw3xyUHsfpbzAXpYvZFw1yzCfe7hFzWWT4jviINfJ4U56vu6NVKp1lTdv/Y
r7jVirLr2CabGoitTuXNmfROdpNSqjEDcXNfgRCwzeyE1+adEWnfviplu7OJDcQCutsmkfYX9OT0
E7Xu+GNiLscDeawVn9iusgpMRYT+9xd60qEsfBoRUkGTN7zpyAQsXX16JjbFH5XJNmh2q/hdjmYT
G9DhPjtbfNnnZlZUaeHOKd08pr4IdAUNs+zX69srwNQpZh76V29GMZ6ycItYr05z7HXID3M+uafR
sk2RAMTrI79k11rBjG5VZqOf+Ve8DeRiBdLnpp7TlgJeXiEmKCN8yYxfJrlAAUoSW3qzFRHKZCb+
JCiT9rF+7rFDReWvFSFV2/VelEKWIzIjz+lFb0mIsjedGJ7HFMcDFCoufEF5we9Q2ciXVrJSZyWi
GJxSmuU96s78Et+BzxoPJyigxfIAT4Z33WnboGW58yCor31kJM/gegCojqPvVqsjJ+GmyAkZT7r/
9F7DhKvl0WYCjKnJVj1TImbtmSb8EpTR6koQJzEevOII28uDWUAfJXRzOUW6rnVNSXzZdYH3No1I
rfpagRNprh0IsM1w70TRT/MHkGhkXLWlHShhsThX4enqtafsqiXt78pK0/uBSQqCjqhpxFXhb0q8
VgDPACEe0ZkWvaNXxa2XUaW745+ZYHGutohxtVQ/NiaOum1a90vNM2yEMxDDj9bRed4BCAM0upDh
OfrCoV+z4inyf+XLYX6/9tgjXXvPhYKUAtuIyCWWNZd5VMwkCyT4ymC9laC8F6mXDiQK4jgrjnae
14Ssib/UlYJCEtbe1BkhTFNZ0c3jZXuviyLVYalMP+IfGIIh5bxEnJNt7JlraHTdpwvBnFIxezXx
/yv0d3owIXv8MRdsEZJlhZN1awlTQ55HOcrkGcpE21XOa4i2IDR79xSvT5mSaHzYY1sJO7DlHVzJ
C9QZHuj3eKRPEY82P9HB7YqoSdLusEd/eZ0sqMd5sle7UubXiiTxNQNiAXxv8/4sFcRPhcAbLzkv
/cqefHnR0ke9DkQd8iCHk4SniT3Zf7oNY16kROrnasqDVNJ8qzON3O+QksSrf7wfiqk0Wl4e1CV4
1GmBfXszyPCUvCd3JdHuYItfTdtKKN3V1yv14wsTz77GCx5msW1ARSUwAHHk6+Yj/y8XqI+VuZEu
lH6eyU9Jr4ZO1HW0Apm969ETDGtXthUQ3AKv0b1k2i39oXbBIPfzCeXRWtYndXuWcYaKArsa1cyN
S0m8G76YUF/sE3wq+OpC2rxQixu+aZUJwnbzMSv2ZLMRl4mm+w5L2YUmdf7Ko+x6X6qhPVU3l/MU
M/TJ4TqZQ0AOi605THXf7pomJxd8EdcBEJaN8il7AS0ho6g5aXksdsEFWV0Wx3PrRbAQN6K3uynA
d/GYBwco//7xDf1GjKLlLXlVuVy/nZb9urmLpYGyADFnNuigx29RdbbWaNn/+NwB7n2FxQtK800V
xDP/qBaqjBpjP1srXosIvOlx5mCuZqs6+60PiNS7a12ezaUUtOJjWBTO5I56X6bAZbwUpskFHX0U
lRiURBPIgUA5S4aXP4mbOeGuIVyhSt8VuDKfLcZtipoeHnMimOtBwvRT7UrrtJBRduGA+xsejFCv
hr8LTW0uoruqX7e9+ADZqNPSkdM1lotSqMKJnJx56e1Q3XiQZdmZvVBNo5kjOgfZ9i1beB4nPXHJ
0InaWNmZMamNXGOebydb7PpQarI4+MwJuGqMiiN2NOKfGs17k+23LlAzIIQrWb9hola6Gu0S6dAZ
p1S6yuTosEPhTiirsOcI8Stgfxj6K8sKBR+VclFHpIP9w4l+5WcKAqQhU52ySmeVRdiyXplVG1UR
uuyRPTBMdkN0sCPOT4EdFTZ5aYgPHOrBncoCOEI7dJ5afMIEcoyFlYVzZyCX4OwWOaiB2kVf5ZSe
YySX+ONsIbyQmyQcIe6q0hkoV/+3xIBxfal3pim/fOyUkPxDsPrakjFByBTQNhIObvVGPl/Rh/fe
No8VyXB1sCZweiLS5zf8hZ2N+oTPw1FjF4w9PGry0UQXC7aY8RjDmYJ64fysLm1sW9eBu+pA6e29
BcJtu53J/tp3MwSg9hY84OirLxzc9p/w1IB5ryO/nWSoF4Q/emzSTpHYQr8QjLE9e3uhzzW5S57T
SyXXEPFNe9/p5acNCGbPePDDcNyrfYR07D0V38hG6uuOlrPl5z97xPZNnQs6qDVAsQjLOlEmqkyz
AfZcjsdPqY2SAK0J+zlj/ptpluJ8IBiRbdbxrWwV5O91gUEcAtCcfq9QKvURaM4jvBeauu//MLaJ
FsHrdhUJQq+zjgYK9KBf3e3P9NZt7jg9l+U50emYxW8dF7cEGdk5UfBS9LhtXuFSlVIT165tiaC8
sQ7MXLwWFJnOqaeF7PXawgWLS0ndcIcVv9UPeC8zV9tpRDPkhhf4+KikMOgbYTK4z2uf5b7E8hdx
r5GY3aDxH0CHGqY1gQwgQGngqrr5liCqITyqdZzcTV2HOwzBbiZ5qoxAmlvCNVfKVVXAdgThKqZ/
tCtqklQf1d8vIJPNrchxYwRpa57WJylIfgtkBFG4ikNus74p8EkCTPcu83pE4aCVt+o/4nODJI2y
AenYyXWqk878CdkRUvc0wkCO6d38X1Ks4n2Ug2KgGLVAcMVzNfdTVtw1cJLyy0T8dRL6RkTnB07t
HKc+NBA7hB5zzIpCOl16giffCZPeFkthfwGn4gpMQZtb1fNlmU04Nvr9b9zxjPIWhLkNL5ZJcPSN
Q1BDckOeyBaonLNpcqrtveZMAhII9CjrmEU5IB3GN/daIAp05pJN/PM2JZArqFMmW2l/w9MpRP1p
JgBEHnLJfKxUDJgqszix4FUQeEG5S2X0tKh8Ty9TbE8AKNGIMaxlVpqE6fpUf95nSm7LJaRFk2KZ
6FmWTuSm3qekRJKYmR9dSaspHDjeko65YAylV5ZejoxU2hm1WZJ8WhiOAYSApBRvqMAtJ36tVvx6
Eynft6e3lrSllyMewlASTiNNXaDSqAiCtkwLkjpWqOpeM6joMaG/sNRBvw4Dwr5w9l6KCWUuicn0
aMgSJNm+KH74Y+aFFwqgX/ZEQeFJ2Ll8xSJ+2fTRi7vh0ays1wwAvNKtHrQSzTtgMEkzooEx/COj
jrKEBEZqQsvTClHAPlr7mw2xFDBN6li1BaBTec68Yc+QeoM/hZ7Wu16ecccC++lMaD0QAnTosgoL
pVUe1I8W3mE3gyKBjogq37Q8m58fjvXEdugys5ahE0/XaZvlChel0TKcP6aRLqHrSCs2iec9c71X
OcK/q86YuLS7S2hsWbWAjp1z6PdfIWhK695oHBkDeaDYWrQSDsevx0VpmQb2jqseF9s8wGkoboeD
WFVVc9i58eR7xriziltemwO9KDQaWKj5XLDwKbhTHHCKqWpCIwTj8GiUyXrnQ1Jaw7f+ojQAG9iy
aq2Xc+8Zh/chkx4akoJpyZuDMql9uDDuao4nd+7recbB14bjLZW7k7//3gto5+wmHmcSabMWRmMa
ikyITc4tvKye0iXVFsMO1rgNmKPIxwUj2hvav6QM/fZyKG8boU/YxMgBERf0haFWIYpJWWpzIn0i
pjUl/GkteZE4umOgdnmF5MWtAqMR49dc6A9LnJk/HV0OnFbuAjcVJ7UKbk9gaz2LAxOOepfNoB8J
dDmnHCpR5ilL3XwcjxiNgqJHLlp2VsLf/f3B9uE4FXpkPY3+M8Watii44Btn6NNnPwKzv8h5LQdC
oDkNoJFGZuaiWk9hNxJE851wWb8a4l2fAgacn60vNdv91nIzb13up/OMAE4I3I44RSgxnVjqs/hw
w5zdVbjT4d5wLzkNuT2QezXuNgj5Tn0+rl5LDww04A6ZDaqPKUzWaYiXazg3fIXKCaEimeEo6xC3
jDznttCHCSYzW7YsqdFym6dE2FuOE8K4QpJaaJqZsgeB0aEgg0/xz6gypPKbEHg34sXzJ3SQ4Xco
c4DbnbP/7S2m97IdN7lrU8dShc2fsuebA0b55RMPADM9r3SCg2g+5p35rlRBmADnpDG1FDCsU4tH
bCouWXZgXNfKfrq4ieMe2SzBOiWAsNysqRtSWHY4HYnmymSt8iEp3D+imx+056aFrCYQ/aaanYXZ
qUTI+5dsMZ0BI+eto+kz8U6ojdXXOfv2s1tGKUY4vzlHtDRO5dbi4xWyqcaZR/qZwMll5lBLnH7P
pczUKs8HfNztuZw088wkKl6oKCR8htEJ8wdnEvpa9z647JhZNWPBES5DZEyvNniNMNUdFGx+qtac
kqpHGWhh7GKTbfwph83unvVI4IQP45LEeJuQBx7qJDGFg3yZF7somQk6qgZgaAC+rAPE0AMVrXeF
u2shktsrJ+Y06wlA65Gm7rH8cDD95Sey3qrv25FR40IIVWmpyo01iDGyHmTsfDL8xtWb0h8HQqs/
YNLP7teJ5RGn2VOoM4kA6VhFatHlHX8w3YpwOBm2Ep5Bc6Zu9zAy2Bnvg8CppnWXL9YddUSJ2RKC
t/XGBvViwYGlu2ltwQZLt3AgebyxGW6fAVqs3Rr9Eo7Da6CS100cvcqitDS5WrFi1PfS3MQy2l3G
lAabhw4xGGb6qkclGmBOlohMCiuzoFGrGUHTVDtE2q48tVYRo5H2yWLsI8ZhWqfu5ISsiuv/yPT1
hAnlcchN8r1coDXuMWphi9NfLNMSlq4k1Nb0uERAHo/3r0w13xQkyvqRxHUvTPUyorP2FGjCbElf
bCJjz2SKtI3R1GN/w5JflAIlfLygEB4KAhZclBR8cMkv96KuYZhndV3miYmMZYZmjvS3IzIUrmvk
6S5mDe/mrJET5+vn8y/CoLnVp18EaahwoJs2FCaITZx4VK1HtdvpsD1VUFDzUmP5EdTeDnxD0Tff
bzEetK77QuslZdB3Qq2E5n2WcfSoXAo3jDQ/MAM93LEF4KAZ74lleOYdBH3qly9j3dvn4bs9Qsjv
RWdSyttHlH2HrRtmBxecF6kO+qmrxYDSqt2s+9teYkblMaSRDJMgj35LWzSahy4dSUJHoRO49GlX
FclVJvabfQLz70cr47ZD3BURz2fiPJGL+p+w4wIaV7r5suP8La2Z3kj1uELsFjaqjwRzKycsgOke
sdYuZMF9YNCJHkBRo4Aid9f/FjJQIaYuH76Yc3FUlNTr0J1w8I476ZIOdUdNcYbeXStJYXmkdyfW
f2TNcV1iqVrJqXDANtHvXCg9Q3HPaSQnJNcf6RCbU73wvMxBleU+quifX3oh51JDPF2BP+v/qYa8
xL5rMSGecT95DDueEs2FSROlRKDTB2CYCwVolsstPlM1RKvLGnWML5Ih5XRONvwhzs1Y9EpKw4N/
CiyFgBDb5ujF+Us/9yGXTlyGWWqrobU4MY1OnlQ9RG7W0Pdnss8qE4SBvg7dyW+PTzF2Hx+CVEgH
96DM0vCx2pT+3nz5F0pEvbDHuZg/587ouHVVUzDqjhGfAt6ahfjYdhyyVkNKC1m2fT4IeXIo3Gmh
c1Y0cDPDlvdVIKbcl3FY1Wb5+/IuxN1N2MeyJfzmr/eWJR4qlFmhypmHwR8XBAPjofgA4wAPFc7B
B+TYSC7MEL9rdFN+yu0l3IrPYCbep2pWKHokpm1lABJkAMTy7PVqDPtpZspV4lGyC+ap1rLELtT2
7NbEmqLEbV61/49qLJCH4vo6jX2x8WtyWi0OHP0D9LY0/kqxhJNV/TAjTKaXmw2nu+y6XzAYntVz
56rMDuNT+Sz5N/WuIBDFdstOdU9FMCxaQx5G/7IZ67LbNKSo8eHZCWk3ku6Pj5Z6EkQyTSFXZnSK
oVZUSo/+w/I+xPkqt1UeCeM1OU58M0SYq4XZ95KcJIM7IqHLYJoSkW8NdUyb/4k+XDvrv6t57DOB
e53M/Vvvu4PcOjqfmEDzNAVT8BG/1o7LhcjPQOOzdh1QNS9SgnJ7Pwd0FUN5s2XE6oQpNRuNuXVK
qHjaJnAR+kszsS8EF5dmYGMbdqS7gycooW48lqJ2Kpz+R0qU1zLGKFkUyg2KWSIi07HE6IkxqcCu
dmhx1ejthCzJTVuL9x/XoRU2POqndYTFo75V3fcYafinSPy7RTC9sHqczkyOYJo5Cqw2HZZtjTe1
ChI7U9XVsbE2cVDKq+tUvgIwnCZhoBCy7rkjaBh900M+QD9wliGjFNsonjK/C8vHV11Hi7cXoiPF
26vXO5ldqJtSP91t63QL88+bHXGt0x1MUEL430eQ93xLyeHjK0Aj8XqXzuAR9vnmwFP9GbFakkQu
FoZLm4a8iuk8lunDLU0ag5bFwWpZ6jJYsbpU7lLd/T1LZbep6nczLsJE61ngd7VXIcglNC7aNdvi
5u9E0ao+tcN0SGeGsEuRacypuBPO8+FDED4fXoJ9mWIlQ+F8b4o54PnOOPf1kiv5O0TQ2aRUjO47
o7NU7YWqDZSiguyjpnDupLWihzL+RNk37/DqodpqVvQHjhcav8YRCoV7m7slv5zx2qf+38UIn/mL
JTQT88vtrsBfsATA2j12ZkEs4Skz7n6G5TPMxs+swqZGnxFOz4Cjbw/IBkiB3M3NkWTkcTPBMG0R
tK3q2tRW6DbEkaSk0Qh94xD+VDrUoFnbRtQRYnxSQtaPEVZeh+5KwI/RErZ5WXIxYd7aX9OWjxUP
7kaE0oDL4dUvIyjjNMRVUnJUvFODyVL4Dd5F4+mC8ADWYbp3SOibILeDNGGKAnt6Dx5g8kDE/orM
mexdhiKa14dhkHVJouu9WAFbyDRx1TDGKkz4tSF9dKpQf+/+x4/NW2BaH/xPCZAyb0TkylR0Mfut
FJTS8Js+SoBplmxsSlTOHaWPh27Q4MmPhUAZsA11HAoiTE22xG2BYc7Pl2kugHVgY5pxcmBGGz3I
uklazfA92HcawZW10GrrUYgqPF8LT1aS+Y7gSG60Pa/Fd/qqkgBNnQiOkKd5QqXWqjEaXBy52jIC
8V+5QW5AX/ZvibOQ2lwi+5NYpiWN/JZ7H1OGK9aN1XhKEBrqqKSJ5zckcShnvBPpJaYOeLpCjwZU
lwbo7BStkDak+djKVOJ3TaZ446fB1sRDAHWrbvRBQYXjBp9qdMaKxINxJB3i8jsN3G6SWPtu1CXD
XK7zwSzAwIwcE56XAJHSOhb5+sy1VJUVXtWrdQuaYM9gUKuKNNBCv3xaPFEg2jqE40Znkyhcvm9X
dol/5x0XIJMNlnSVfACfn11PfMzgObueJ8uoegULff8ARsC7yJ1WEys9nrrqd0B0Ap0mXpYaodOV
4B3BFgcyeoUmK6D8/lGU561fQeKn2T8XMMwSScgkwQdDH4TK2fIGFU6Ln8MY18ab9blmLgIWRZuM
ZbmcIEDfXMqNDf154Mq5xEMelvdRr8I2UoP3MvDfT4FhCm+69EIJg1AgwoEs0EWTxc90O9MHrvFm
HnfsG9eP9b6fPBUohKEBdRXSpt48Ue+qJ/cP/9kc/CfnpCmeLEfI9P1d+1ybfazDPtf9Z/yEpRDU
97Rw3CS6/EEw2NAjbfXJPHbZVxvDdNy0EJagQjS/XlGpoBNzFPFB0C5VlH1zG+3iACOTHQnGr/yv
KFf5TDVY87CsVfKskzpSAPRSmzQmNpt5lRKZfCzzXk3aJQlUYvepHFBgmbzY9xGsWwVOScfuC61Y
jR0pct8hmkvmZndX1q8YBwdASXD3tobzOOOl0DobgE6mEL0t420QmPE/gHutb7y4SyTFJvrAehrF
zrzz8z7OyifcqLG9qiK9fXDtYmPF7FJ7Pptxk87CUWYSPhvKCYpFnvUu2BDvg2O1tLgQRxBOFaKd
KI8z2WJSKPnvC115jraz85eAghHmNEOyroYUzFfE7l09k/uRi3KHNdUaCrh0cOyi/akhSAMonWHr
2iMYQad+0G6Yz8z7CpY8Gu/UmFuu6Y0S6ZCzlTjqlpCpBteH+C65y9zJS2KsovVEMsOrnk11EUTA
7DkRubbg2cDXL6t/5AQFWrr2y+dqsqpu0oPDvAAanXJlBt+/M6apUtvTUYDHeyjDfzjjsTLbY8MU
nWu9pPMWcwq9In29IdnUi+MwevFhblo0g4R0fiYoj2i7GWV/c0ebPt3jVHxvxrZScRNKvavDAoPl
Wng5RB/YmU6vKY7PurLBf3oX13vSPUsipjxs88LX81l3SmmwkTwvgjmOQ9I88VVI68NFEdmVCVhk
t4bU80wiER5NCTasTO0yk3tpLZ3MdiDcl8yhAanYT7bcj9whpI1CgNlmovk80PXYQwlXsWtJKBqp
vmKsyHgjT91mWEyDyFjwQCBc+msg/fsrx9n2+e3G4BMMaAvyPyFufKUnNFWT0Tqp/CuZ+qsOzht3
hnGpufYIVQP8ms6ag3MLYc8Bw844tQXEe7cbmT0rZ6WsVYsztQK/Xe94sVPTuE1L/uDnQcao+qbi
5WwHTaqw5A1ffJtDxa5seQkWhvhsS8ELOeedjbbbalQX3he/q6FNylgUy5aKEzTu23Vcu7JfSvMB
Nufgoumw7EEu/iiAk7R9LD4ks+byD3zsWTm04OYtVSIzJSdz/G/hJEcYFAouaavvdLpPKAkd9IKM
gzqUph7tGmbe5f8hFuxJzHzWZV4AAFwaaD8DHo0dENJkMKyn5+XAS1s7T9pNXtQ7Z66/dqPFSO0w
ynLBXyqx0otuJk9H/9++6Pdu/ERkSsYi9srKDK0loCXnXjUI0FFsFpg+MPmN3nkiXV3xtQUluAxy
CjEiz2Qemm4NojR3u3+VnqmfxJfcXBaGVgEmVFFQgR8T/tIWNY2AsSabvxlMEi+VfowxGJTr26l9
TGlw1xpy4kA0G22U6cWYr8O9s4UMh9QG8l1W8UwB/SHHxlhNG4R4hClj/44MY0CTjPxExUGIx3pP
71adQHgf5edfOWARiZ0L1IGrgxzM6e1Mu5D7r0o7gfdvuGcIzTnqHjKRqITW/9gZM0AqTvoL4LEa
L2mzRWtEMMCiNQRCUtEFK3mutf7yLmI57oUuCOd0X90iTWUDlo8X9YkpvlQOS48D4p/kV09DmU6G
/iTaoTlGn9TExQcj+ZXvNjCTEJVweyn0QLeGFjZK0NyAF5riAONh0fMiH/LBWqpnKw6M23yd4ey7
BCz+Py2rMDtuozVv05dtE5E7SHMR6noK/aIiF+/yC8JBdX+0BsWCvDF2YchUI4A8jKi0MAMd2Lbn
+dL6RAH1fiNQEDKqbfQaahAOXmLZjvovyfhUfokyDYRxe6csJJ0qx7kCOwcOJnVDEQAcwkxApMJa
DfJemh8BFjwTiLiFZsjPn7n2RLNBSdRC2WDMhMA6FH93WAuYs3yEDYhogdf1IQkIUmhDZrnpz8XR
Ac+AlPAZrwH65u91zltb6TcGAbaNSQS6qoEydvAIjPHy3W0UpAfbh+WjjYktVrUHj8b8+l9gk9EK
+ocYn29c1JV157GyUL/3Q1uleh5xaITafmMKSl6OHaIPsO4A3tM/qVpu4nnU96wc9JxhGdJRmhhe
jyswa0gwU4cmRYVFf/mglK+BGJ7c0wsnXtpWVg0jQBjNo6e38DHgJqcePpdNL/oK0WxQ/Z9KLs6+
rKHC6QFwC/sc1F+7BPFcTCBar4XToyNLX4J1w/HfC5zhSQ4mEPM7X9jfRMMOXKgBiBup/SErnSmI
aBcmLswITLPboRzo37Q+ysQGAYK6fSM2TVrnIq2LA3jRr8nrWlSW6vZJD/ndih5giUx9ZdvXV7eI
muvQikudRiANQuFWpBHLGX6JdlZqalkmIDyw+IAv4V9RCnlUHMdZ8TsWmOruYS83GjBK8PxpEjev
JW58DKp+e/RObEH1yjIBs7Y622Dy37SVcUoRCzGLa2E2ZIQ8czIGfNuxViwXfWEzxAyT1fyxXJyt
PNPUs0pdzUYrF3DtN37DGYfxC4JuG95XCdYmAlWLAKCVWloFXot2ttCkfTQ2/CeCDAw5cAOLlWIX
sEXRAyVg/kgQl2NOPfd4dZ1DwFZWSYZESwFJ2KLbH8AKkvH1b3wa3lAcfhWIPOtOKjE3spTINAGm
xuidG401gqHRZTve94Uu95lPcdeCxFf0MUStRsXETZx7QbxF35ZA4nYqXRhpOnyOkZ/BTRNpFysM
VpBl7dytajnj5745jLpuIn2dSlYQDXMBtSIfQizWAQr1RZ9ykibqNtI7kIDeBDQTuIPC1uSQr6Rx
J87sS+U5SNe9tTFsaGNGYzzmyicFX2phrfTD9eNOnHTkNnIPtF17rvAXqzY0NNXbr3iu3aiagpug
nMdUx3ZNvuenkB1rcN/pc14MIrwwimuCf6obFZ5U1oZiE1+50f2wvvoCAxDLOkMwFRwx+IdGZLqi
hOxpQkS5o9RHtHaqUHUy6yhKs3N4LVq+aU9gjRFBELoZ/9ldIxS67ILDRgUAuqHukco6Moerfnvt
0RMZwuleWHNfbgjScs8AIRxAuvsi/72/vIeifZwRPI65GK+7pJkLuVls1Ucpez3b+v4nIMILNB5m
Q4LS1JiRbBIhKtfqDVYRyOImL61k9YUHS6izqTX9I1g9JWcM1wX/rehicxaxRU3EPbDhhJlzSReP
IYwYUcczfHGik22DeNMMbvIkZjIIhTocKxRdiNi64bjTisS0Wjfdr3svpMAl9xFeDH/nsJzWl+TK
/4KEuelNvo/qrflSalbbMNck9aCLe53AsA4uLtz4eiPzJj3Cp3lMulBIvrEzrtSoI5deO0jKRXDS
8RXWqipPKFkiUeCD67A/5eB3+fe4IudUyqdTsfDVdReRmElcAfVHPb0xpKToZTwcJKo3xMR5ILYR
RabJ7esKsB0Ws0xAsQdlP3a9ka1ltxiwkUqLT3QncuyEnA2xGz07HhM06cSzQD6dJBgZyW6paJKe
lmBr4XiytOHA9S3Hn44uOELn1ABeJpIDFMwNlzKs6caNReWgkMypNszqNeHaxbT+lF92C0Ep+tZ8
ltsvcrKtUEGjUp5w79dG4wmDC9oCZR01NhkaNpCZ+GTfkYrxpLsiXXFTzNNs1dzhJbp5i8gHdowT
02j4LI5kqqGAL5GT7EMD0P3/zGH2F2HhOStS1kz/O6wPEkofKSayPSrcXNAjCKnFTUHkXE15szeE
R68jrny1gbcRUmxy64H3eEIivkUt+zxfA64B5AUmJ1xKpk35AFboku4cOGRdqxe8Gt61eTgSsghS
T9HZ90xWrV/mWqTfzl1U13KF3gRuqk1cuUidJZXZBZX/pTWuAd5/YapHtQk2IwnocxQX2huT8bJK
MAAIASUJzjxIEgKgPa5noeOqKIQC9wACxfpamBednuJeYjVWZsx34Ue+Go5Pz5+fcW/27LNF0rLG
ZrWbwQ5F3ilivVpZDmuE4zQ9qQfb/fXNFpeyasZBFHt7RaTw/0O8HQY14IqKyP1I15uWSVbL4Sbl
xLjE1R4PfZ+O2xlA1BmVtSRlhAGRtz/PMlp6dYkHG1vuW+eMxJY9GsrPv+48pYk1qqwheorOqUIg
QgzLlZJ1q+eXrHOQCUkpc3zD69CThCNqUrnyM9P2nFDHkjLQv/fhPPvlj0kObZmDkhBzSiHmxSir
JbxjNHBAe+RHS7qWWPuUdwjuOe2Qdg7DoPYWK9OM88f50BHe6IHkklUxJM3rOJkzZ7zpqe8nq/Pj
x5YZ0d5vYU863u/D+7f0O7P2Ns4YqYXPKV0gCI+MEbiLEVZ46w1amXMLoVJD+1jDhfRlkkV5uwS/
r3BLfExL0g+FwJtpz/OJmzXJzHVDhhwvSKQCG1xPxcLqrywLy58mUatvn70srFTtOtTh4vI6KdXx
5VTG48ks1akeE2MAYyoeq+A2xQ7sBP1YC0MFGp1phc1RhHXNHAZi8dZlYBgz/sm78uAmxev6keqi
3hKh8YpS/R4JWx3RrQIWF3ijzQv1hHk/hiRtnyti2HD++nPsiNWv4U6rMEWLfn3W0stEdeoqnecR
MHG1g35QKcfSKkoJyBhoX+uu/lFFZvbafV2wjBPIrtegYe69HeUQJNje2689rbpU1XEBeETDcoaI
XamISjKM6ZRRW0P+E1/W//2JcSDjaad2GEn/BACwaIrJRL1gX9R8WANKqarmsrVNjsho2x8UwxNu
RDbzxcjx2i6l07Il6uGHuHkE0ZRD4V54S2FE/jeB945/TK0OAyAKgVFasigtwLWySyWzOixTtKbw
3dlnnC2C07niX53zQ3+67pnDQTiDKOLUjvLgohX8y0GKYRd9qutRIW8TQ1EcB5lu+mTOFmDpv1ex
lj5rMNDc31Zq9NyIzL5ULxHml2H8BZKwP1Gwtbt3ThiYqe0HnuYILXKwRKOvBN9rGczOVc9aeUg+
tBbXiNPVXW6xda4IBWeBmFfhTHMX/IlGAQLEZVJ3kp8wKqLuNXgMLb61do1+reB98g72r7Hyl99R
ABiJsOub99WBVtEkaVoKIT+8hqRwmgABlsBxV5X7IYbZS60jrLyLd9VaE8RoC04tDjoPKjBaotR4
t5rnZ+Ie7FP2/g0EPEmIA5G1FLHY5UNo84944jxzZQKtoLp1mQBGCjEfwdK+5Ecx7pOfeV2TefbO
j7HonrogkLxDmkcvjQkQKnHU59ihecVKF5ZBEecugNKZA/2oUb3WqqK55rHcjOGKXCqysPMHLm55
pUXylBV4zQ4xN5CISjZkqY0jZVFkHZDzYrHus/q2GNxkJYPnwGDNuiZa8LAvUfdRrcFaTJ8ancE4
xADJmTu5voIvKN/Ny03WbwBr5fOXd9MLkvm4+m4CgDeCuhoCOhYOFKdLROlc2r7JxvamdvESlb15
2fWgK6XsUxGanelHpye/KXCeNkGe1G53e2b5uYcIBgq7+OFB1Eg+mdc+P1ER0BSXZgR744tfF7I3
5TrbyUTCv/2sd/Q80mBPIC40tNKIkfqXEJtYJnqU5NOICOp647l1aG4bBm8csaUTZgSTdDOkwPgU
QZuIQiBFEG4tX2VmaB5dLcQFdiaQtiTKk+TMyA7XQywsVJ7aHVL6ti+vqtkjdlRusd/IIq2Qx7yd
gwJw+HkwnlCYoNSNQZ5nk2sqOiQR92MT7+mKirV3Tg1i8HGZsQT2ASWkg5QDa3auEhG3ANt9uN24
eZuTzhJYD5nsr6WfB/GMX9tnuB3Yl1zEGIqjBnJmewcMvbOwncnFQ8Chf7rQZOKKADQPXlLkgSiK
5vXkdjNnc//KynFRBITm8/IR/nMScAYJ4eWgF5oeuruIpKbQLw+8xfP9pMNqhwmBJa4+SHWpXVos
YCjvjZpdgHHH3h+PQIjd4LUXO9a+F+XwnPEoGMxNv23Jd4Ujf9wcLC/vS6cMtMyp8IEQDPgrKKXD
40ik0KadLx6u15h06gr3a+WRRAKpvNf42F5eqUNCUilvYHhzwiqFiSrB7SzZTM/Lj5SGcXlnfjt3
swHACPF87ZU8WaOF0qIpz+KIJD9YGWS71n1GQl2WHoNPf6clYxZo9nXAI0c/sC2BuYDm2VuAMlk8
yJrV0yFNb+TvNKZtzJ5liJl1beSDsOa7Or6ga928prAD0QCQrNYqkLx1ccK3BedRmOPK8oBwbySy
wmUBLHbEW7RMnz2++NIeiViUG6Lir6Zlxap/fCxlJGq/9quzhdrQrNWXuVvMAWy/vKGUftdH0BL6
v5ngEMCsUCE24X2Vr6N2PGJy+ndKJJOAeHnny/TILBR0uYBktrBdPGouqjCwmZhmf6BS74Mo1tqV
6il0EpBeYBnctINHgkGk2e3dHL++tBgn3a15A4wrF/ezewE2wqniHUMTTZY3/WMiFNJOw3uidWPT
2RibtWsJAbudwVDyEVo+n/OWLNXSq0TOGXAj0KIt6n2fU8a4A0SLnWh/hfeNJet0/8P1RjnR4pRY
/MXTqCkdxItDW1O94aZgNHM+nYL6h/EE2SauiWEA4WsTe4FmAJT5UD0mys8VdSfXsNIFl3r2uIdi
AKWEMcD6+PcFISbh2SX4X6fU71CMujGEV6T3RjqzSu+xhzYQKhKWXYUmnFwTuXLxwCuKSYC+R8Um
XHGf1S63KjM/rqPyNho/BXyBrXvFYL+UV6U+Uam/r2nAcWuk4eX7Wcgz0VaD8vszifMN3iVoICn9
Q95iiksqf2O0YLf3ONjGSOwz/JCzk1UtFtYMBAnpZX/HOGePOayapboGnotJDd9MndHgVqJcsE9D
c0d0TVEhwiA64TRqPc+cWNAcDbKRxZ2s7OEuAGimj/OubA6VrKCe+paUgmof5EPLee3JuvqVHzmG
ziOS5tFbB9QwTLxsraz1W0lyIpTlio7j4Msi+hCh8cHeToCgrljCbRuu0mORvGGGbd2FbGpU/TK+
z+2iO59IuVMZQ08h1AtR3gNYOKhbA1TnulpyV8TKYv+AldSICmlAeDvBNZ5a7e6IeAblXPn83tSX
hm61BgGClXJTg65xmq4O2Fj1KouRxeI3/LCg1z9WsXDWIkbg7/1/d3zOsCEi9Nh0PmiDwvVxqXfw
3Yf8yW+0BJmA1xtOnA69toHQDXTAkMkqqmm230VIiXnuChESc1KXAUq1zm5Zz+ME+H5f6QPWaGYf
M9iPB3h8NIcdWWsw1yruFvXOchA4y80vBtBRA5XtO1nksiDbNsHFp9Uz6T+/rCGFSIPn01grtSr4
JofYRlLim+QdYf9Tds82phehfL/he7G4qT6/4UDQwlw/J3M3jmyD52kw2p6ID/fTn62UPpjNSes8
vFt+/ilpzliR/ZXwvYLVnixj18Fx9KRDo3QrLAOomNpz56Sxt6+IKpOV77Emj1UKo7+deJkokzaQ
WHYkqyFkFDXBUSlEXR3Oe/e3AdUgK8HN3iZDUP6cTiIU+3OgRd8btjkD5yAsMO0IiUlFbFUHiPkt
fVKWtdW5j9lSm8TexXPuGfd84RWSvX9dJAJ8XdlEjoxV9+O/x3PHSmk71YcOp+mMSYLMTayp/Hct
RbmyXtzTXNSxMJRvN6ftvDUV+WatYzzpu6zVNtqWFrZPhcmlY2vZqI068SHk33ZDlTdGNczVE/Fc
lnQs/ASkOrYAMI+E6m8oYF/VYWGnY2J6IphymVF8o/GIbGxqJgeRH6/aQuL5Ooqc5EPbxXuNLQU3
Sl6X262wg9Hck/bKkEn4kRPIcN8vY1wnOaUBOLWdV+laHdFa4ureUlGKEbx0W1kY5Hx4DxUh53WP
jyGkWQGhoZuM0qJbELnm2sXBZ6DIEQzPFfS9jRBuUGN7b/fiSX1Ji2dJfWalvhBtTp/GBidErQ6S
k9wXNE+zL7Z7xIIv/XdyHY2TpfrU72sGQVEzosDgchDLRnFF5lmMmzVNGnJs+KMyNZzdfyEb/7rU
aMg2g8JXoIF8WnS+OD3PsqeMQooTT8do6JNIskzPZOZC7smESUMSSA1x2pHNnsho7YwKwhYfoOsO
GZIagl4Q14h1mGGpjrZzBisce/r3/uaKAEdnJ2ntrXoFsFWkHTjqhzXMeIgiq0lI0DJGOHEvfNVU
gSWQcjt8zeeUx3Vk8H3bARTZk69YKtKU3sJor2vzAZ2GRlDFczKT/ZbbONTeyn9z5cZifTe/Mh7H
1TlnWbc+jhqEfnkKVCyX5k/kgOWxWWqDiTdF0BMc8dBtiT4olyA4bubohOyumI5dbq45zcTpQwa9
+cZ7ILwO8twmt54+8fC377UqKh0AblzZKyrh8Fh6/ueMeYeiALKw7XgMZ75WjK3GKu9PToz9IQzV
VIKTZO980uVOOYwW8jGuFQJz7BT3W7qEYIaf/ZrfHfzRfdB431d/p1Lao3tijiLFb0SWxdcgBEm8
a6c2h/8H6tqj+aR+QvO8CX9Yeo8MjZyDoStf4UFRTZTUD5HZ23qUGNyWmodf02FPGwJcSmCIc89g
DrLFuOrI1qZlguvKa3jhnrnUbsmZ0tj+hgChDt2NVUxQKddaQam6zPlJAIKzMbjHSbBH/zcAC5XF
U9OvQC8qlsDzGtLw7dnxs2hmNkOTY8sitAt8U3igezQYhhHQyPf/Qjydzrok/kzTmnPTCu/WBRQl
zh250H+c8q8d9CyfRa2EckU0tqoHfdamY8d4Nw78pAUM/cG6q1NrRL/Vm1I9jPhkSXGh3WTDfVDD
CuTpAj+vD7wOCNmg95sR8zytgGcUQ1W3xA7rXEO3EV664nr8kPFkmodObJaO0/6POazrXIdhRl43
XUNq0Pu151JJlBuadbt/vIrSJCuLlZ2uVIdbH/VlG+SJy2CYK1DnN761318oQcctI+BV0MRpJXEe
gK76Yle9reFgPx5jeskH1SNkpd/XedoMl5l8OOp1Uc37GNXRMqiF+1uvZSB9dNLDapPnuGArQXU/
V81Zxs5Y19vL7SSTZeYAPmYK6T9E5rbTecEsxNzaQWJRqy7gxl32kcEUzw8ZKMWYM3iP01NRGzMQ
nZkoz+U7wNZKBv+YYqAiAiD3M13zlInsL9hDDRO914xRWfK8Uwbzf4M9FPdeNMcH8j19VvOtJ+6p
Fd3VWT7wQmbCSlGNJlkwRp2xu3xxx8JdfIh+pFJTbOpOC5gn0qIcdkAXOWJsWaxO2GgET1xCgbdC
w3BhHcgHM45giEUdLwfIMHO6dzkfaqyU9ZYJAvxbCatDR9nafny7w1ASH4z4tyfYDZ2QGlvLoSDG
MaA4ROoU7hnLeD9g4mCVEqBwJxGfcqiYLICeKdrZQ84OvfMIJvobR2lYWkQXLJvBiCOW+ck/nN73
bv+oq5AQ84M56yLjJD3GXM2rfCX7sGmx0Qy+wH0KDyd8iUywDo7OORMjiwWskptjYTX/QoOUWgEz
lG7OYH2rzX82i8UI3WdR8IxymWP0oLZdZo3fwPzettKzq9v7dtclUGoQZ7Eq0HBrC51p808Zx1Ir
7RAFx24aQgRER7Et31bt1lW3ZfKzwq2f2lsWfcXomDGzVEONgBCHtpWOQoHoR3jyqG4hUSH7yZFV
Fxx55SGH1iYXZiFnD3a+DvQl53aB/cP691RrC4nnmj+mla5wf/RQQ5CFQsio29saHIDvkDwq59ss
fuh8rTB3VzEMdb4Ne6+vnZOu2aSX9/sARVOCg1eza2PH3yUXSgviVVcn+hh/0Rqb+XX24Eye3kr3
+Ze5FaX9rUjreYMfnzryRngNzS7uHRdGv7sk0x1Sr1hDhjBuBUUVd/DjBKB/VrLF3O745bBw0z8v
3UulZQqg2Zhst5vlP+1qMjr3yn6gg5lCgUVTPMdhfkF3wK7IKw1QjH0NRqdz1xnLCEh1nxvxb4a9
F0zqU701G2X3pBdrt5VXd/qdcWU+6AwMfH/FI4lW6uVLmHRfkjA6YLJQWOGj1CEDMSF+z4q399sj
R/BHPxUPGeNwW9jRpt1GfpEIm/L/wFC7LxvRBu3vrx2AKkHFVxk2s4B5GLaAOHIdjtGLnCNrCBHx
4Yb8uj286Q4PS9DBWSt0kihFkRHzThX4Shje8IyKIvw1rOygCDYHxtUg+dr/vtE9u8UF1aVy9yA8
eHIa5DIfB0vyWLT4i4glBs8PtcCD1JkxgFHYzcJdw0Wwl7w4dxKCeQ6U64RW6NSzZVv52oKeTAF0
BaRJNRSMJL1Thruk/D6+A9a3lvT3BlRq0Y/hM1t4NTia8WdWG4PdLV9fD04L/31uB9jo9ka/yBBH
V8DvBVckkBbGRLnOXDNpNS8WlNdXepGI7fgwCfgpPo41ZFYqk0g9mZnNTE4P1DsfOTvCwHn9SyUm
RUxT8VmXmKmyScKnXnXRZPprpwGk35Oo7aUQSRYTKNGYEmY3h2n+jwkVsfvBNS6tr3MutEJ63nCm
rubL5VtIxdzfaSBzWOwYG8KW7H5pmh2he5Uu6dNt7TyNT360j/ATrDsIIpJBRn68XHxwwBR1Csko
uFyA/z+RAAw5xCOXU32XIaF15IdjQqasp4pnP4O0ZD37MgusUEIYv0nXo7VB8kWUQemLQmEZ+YJg
/B3CMrAKhBDO+ZhJMGoozKfr+AFT/QfHkCNJPUnaawqlN8pOdVoRZLjGHgfrTaaDbQj1KY8FiFNw
uIw3m14oRfq05L7ToE3WpeZcTtMFzdE5lppD/Sdzq7TFgF2AowMEJKxxaQppdnEYvsrkJSc9u0FF
LOh1SZnqgFHiQ6eXyOpRADKNUXGT+bj3Fk6w6Ji8OLSGlUqvKB+TpH3W56aNA6uvfXkgKDr92QAy
MdUHsnsdOgvXohs8qqYD5xhAk7dpBRQko9MFuHy5t758CFNS8aCRs0bNWobAismShDEeCMLiHEc/
7KRuBmAej4wWZoVUaNDzLzqP65PbmOopJdC0ldv5WVILPP3JyRRbqPTbvqW4WjACid0zWHhTC+dM
/dGM80vqELiJJNep68q3xmCR4binEdTqkdyZIleoqIrEwtg+MJ7rXVsRocZ+cLMUiciAS+LEZVUO
xHwhF5j0QBCeIn2PaFYypIduGAad9UmbQYROuPL+u2Nvgmurf7MlCx+jb8/G/CS5jJOAT1oro8lz
SAuArBciu+Z+NMGq70R8x3gV7EJynHGJEKoo2nz0WdxDRgp0AqVe9aOI4DEE7w24xVBFDWj31U4h
nJ4DzF5zoBNlqoHD4WlrBWvEafhM9BqNkZE1Me94WemGU35LS2ghnRIBizTIYREDWYfpxel9roPb
XLURs/zSwmF4h7n574k8r7toykyeE+5yADiHt8/yGhbQB6E5KucNHirAJp/kGeRIdeNB6Kxuj6EI
oGX25Ti9Siyrppab5vhaYhIi/opbrOJGg87WF1RzXEGP9Ookn+djr5eO21ctMaVbRkbQ0cR7HlVi
zyIIoQys6JrfwyS3KyzjMmktOOXH9BVg3wJVg8XEDncowbEosqBSqCNTknawqkSl6lwM6pcbGr5y
6/DWm4EPOxCrls5P64eZApndEVEyHy/6AX/quQLm+S+0s7lDjnK9HW+2qAd0+F8Vltwz+m3izLz/
Y3OwOXNpyoaU50392ekUJOmu+aV67lfdCngrKO/Ht3qEghsLTGEWyNQZYwanHlQhxhOA0YO4b0ti
h0bKHfzXdG7+r49fLeRJ75o74ASW4Nw4BpX6W+QpVKuU85wzI+RXMENB7waGnH+wJW6COe8nfeWX
YZ1OFm7oDHl0WEagsCV+mkI0ZMSXdOes2qvDer8Wl9aX25wAGdvbqTHVaI9QS1ev0buSxxCuNaeW
tGNztqhDu/JG2wOMfr5DvJo1CCQuwuauGKKLNHItHoWd/nLe0Hf3G8lj/tChZ2yOEhRURkjaHHMA
F7D9IixlbHfLvYB7ktdFxTjsDZK2z7FmLdNjqffLli52BieCNBiw7S7zXprtiRIrHqpu02akas58
cxnYJjsVyJTbh5Cxh4J0gDD9IYRCSO9kc1FzytW1A5sUQBlWnZ8pTUG0OLpwVncNZU40p6WwrONW
Cx8Dv+ArA7134amvZCMLIQjYbNowfSr7FF/ddraig3Xitj156Bhj/RbOxMvmiPg7trXAPg1jtUEG
6E4AmYL4+bTqiubBB/7rjm2lD27iJkBAI5SJLI/wrHcFDzV5Dxhnjh/t/Rvs+PSFgyU+klD1tPUn
2YCqPTGenG66yt8JyPKVY6MM6/7IVoAaeiDm7GNG8qd1+srYuSwg1SdTL89euRQ2akjlj97M6Ukg
ncCmmfDfnyHfth8absC60ZU4ZV94zrct5/i2YL7KYev8GXVy2AiXi5lSKgqEeTee+19HdvWBZyFt
j61QPllQH0GTXlxRN3c1kB5LRL+U9ZGHF9ID9lmtOzp5HxaipIteep5bqiR5vcaaG/6o4pAkD2kE
9bAC4S/PK5Lx1KuD91ZANFSWvQtXG2j+eSKrtEVxWlna8jQkOnJ2auK6rqouOieTDUplt/vn1Tsl
Ff4OIy9rzeXCplTBNQhSz+2Y04Ml2USQfLf5AwJEVRExloPuXdiT1wimigCvkHyrCbj5OhpGy2Ed
GP/IiwC1h2OZxZMxh6j4i+LSrYCYNZb+TIwRYohJjHxHOd5m2ubYdObMygW2rudmZFa/tujGNI22
2dJibzNx7FGjWCH+Li3++hFh+rMYaWvfAx9jnw0U21nbMBtUDyjUMhfWhF/f5kkW2omE2BDjvCW1
bQvmP0RzqospzpK/jPuOSOISMrcbl0oaKp2kStLTvoowU+VgudeC7x7rPWzjFoL/Z4yjioZEy1/J
BmlvrNzVgQP/HMdNKTTV5igfdZWEnvHBQj317cshSAy2CCTr+afi7pPMwkxVUsga9qQPzC17vWNR
KOBQnqfN58Fk1dNbSBjEs3khUMWe6JcfbbkE2PhDElBWZfL4zwZRDWMb+hCT58FUySJySgPkse6r
qoZriy5tNytSoY2+12E0LcyaNRr97bGRly2RcXCWZOwi6CKgfLBtqW/v4/dDTaaklZKdDa+Gv83g
2hVfTJytWnmFt+i2ed+e/5WIux5q7MNPaMptlHJBkGOWroF8matBaF2FIMImpZqH35XliYtbPbqI
OM9o2vciyQgV7wnXK3oonndO33g5Wm2oAzozP3HPKgK88YPReDQwtjoBVqDbRdt2FGiA+vUr9Hht
tMXoy76oQD2tm6ygETZKmmP3dJUTsAyAfiEOKXq3UUv0uc5jaWojFCG2kNS1Y/qMdIYtwrQWNCMd
Mlo85fkSc1lII/UsYUxt7NIU7X/z6HsUqHtXc/Bb+7WoO6+3JH9L7gdG3D0J6UlkDkXhr2eIH5g4
owjPBCBUNPBmVHHSEOwLMsYz7BOmbtEVSB97fcF/eBWwHYNdah80R+Gh1lPhFsCiBVDSJfLUUHGU
WfTQ7O8d5XoX7kf8zkiAnxFVV70dQI4f64b6OCtc9kXk34o10BcthVXTBSjDaMyhQdqco19927So
FLMZQlRLQWZbG8nfrhLfy9guFPjHdyzOStz3Ldsu2yPTPYH7ZIAVYoeIQjQd89t1BjU8Dm3YCnKi
iOwQO6dzAI6Paq2S6bH9t8Dh6/brdR3Re8p4ZbFsPufMc6us1GM1INw6IZiF0JM4Eyegpb06uQpm
FQd+UZ6HsyYgssBQonNxWLOi8YsgZWTbS9Ou9EKQErOVseQhLp0rb56t7sPUCvRvzyCd/CjnEtdH
0+1H0/zvbq33H55OdNCP7RrR4KhNnRHNRS4M6YOpHrY10crssIcWSwDMDIK35ma9+a92bvnrm0gz
EZvq2vpOF4o+3QwvokOF/soK/+nRPurmTFw9nZqbLvrDfmu+3Tr6Ih1AD/Lahx5pR8XKK9KXeo4u
LRKy2Istro9Ze46M8JPlPgJzN2breD3jtkbXi2teOy/pNy99/XmTc21kdJx7HJDSDz9aR6+t2A8U
Ir+ceOnsjHv1tKURfq3ST4sKHhR37O2VSIEpKnTVhMkHaw+k6+nGuYEAqkOANinG+4LWMY3Z2s3u
rzhtZCzyYoQiZ2fdKzehAdVfJhR9C36LDzVCaDLqlWIzSz4/ykw330n1Rk2PO55PfnODZh1HPKBt
n6Sgf0v/23yS3FiQH+4Lkt6Exqg3mKltJE0D8fw8XIx+R8GDu++A1TUOibbMRgwA2zwKTPeyC3AW
WQXGbPZb8BDavX76ZT6yglsXtGMOKylGcaYWjsCiMFtiGiqO9DYS/iB72V3EyJ11oNhqd3EezyT+
K3990ASz0cnI7MqyhuQq6BMsCQV0tQr3/rRUvasA3sDslNtsXtxD6giNxVGBIlLdUC45occV4sYr
Mck/3PXB21KyxMmURyx5nvjpqr5NTfyP8Zt5leOMlwU2Tzoy+teMh/VAJwS+esA/Kij653TFUDpk
YconQ3VrYlf1Hk8UDu6GE3/rIwKFkwqYj2axNeRQOTxCNUw++D4gXiBZyjs0EKYf/4zZ2geTGGgt
LKgfCa9yLGQxHa5fpKs7rU9w/UjixBrH8R1TsMKwvi+t0/tPwa+Q8dw3iubL0LWQoHE03pD2Bo5n
7lf2S5JLANzNFOSEif9n7lnQ1+eEF7sJCUzgrKX7Hs+B1ikek1IwSnZ0TUT04/Z6xrrTJugGKzoM
06UVhwtnjLFm3jAPrkdNSmS2FlpVTk/411GnELqAWcltI2Bv3ssAuFdQhdMHqvcCnDws4aD0h9I4
u9Rgw+EhMvVhV5+OrLFY9ADL2TGH91pakSHO3NbIDrl+g0NIwzNfcnhgnlI1e5lJu/OgLjp3wLy3
yxsvGS97UG6X/f70ifeRC+OFaYotTUvwWAHekpHP6+Wb1D3qPkNBEsifOyzU7yh1hKCJJrXl7zrN
SfU0zV3hAcCruYW8P6NG7Qe3MyAD33IZTCPbTHmUH54JPUb69q0cTlh6aNL5b9SDQfHyG5QrVAg9
6IvPV5JkyZwbcASehL1fnsGguJ0U9GhTECXjaWSRXa58YqNJXl+6dJNmXZ/XCeqHAqWweLoYFE+r
yE1ioz6Lh/dGNldGA2omDFgJNBe2+3Aas/LrUtOpJFrFjOmcnGMnrTKE1px2D0vhZGAQ6LMbP3wB
+cbQ5CNcksTWBDcXDXrsAz2DR0Pct6U/hLpo97yG1aittmRZkKD2EGp1U7cfKEUMYVrOFduSfhLh
Hs/j13e0W/SOYU2/7YJB8pFq0fkc/sn0ILTu6PchZCEgdRkPtjEoUPA/Q6QEjliLXbNmRT+lnLOa
hWsPAbsl3tYy3QHdTONJbA+ejRRbKaIYnzEo9KDRFori/6vSnHx11Ra1lpVCQd0dZd6TcmPH6YB8
NdHZg9fpqMdG6Pq79dfp7Nm7bTJqn2YSYJe3DmWQ1bcONq62sC6bDB1IKibQItXQ4KPhmj1b3TKH
0GNyot8cYlnRXa5fY9Wrht0d/gxe1Dzxr4tFEUeLMm3BYEluDm958/zxenLcWoX6Z1iwpnPcq/mn
859lHJm9rNUPRGYqgljNjK5rAxO/f3eiQyqUYOjJzovHrSY8A3Pdv6FystLr2EOerl2uVnptmtn2
PdTEvtBqPBOKuthxBfZmr7S4p9fnV55qEn0Q+iVEpmD4qKMQBqR8j1SQmY94VbD6R2i1LUvrzRk6
cvtPcMRbB7b66ctP2ZOjZgkDJ4hJPiSV5RiFyOLTQWGSGHA4FnI4KEkeV8riASB/22BUG5iyETBg
JpRDHWTZOhCVx8tHUzcIDJYfEwAlAVWcClCoWRj8nLZTf9h7Csi1tK9Z/d0ZsjOcVnHV8jpiqS4j
H3xcDfHZ/Q0Z9TTwETyN5EI4noe0lLm7PsAMX+XJ1vvKKvOWaF4aRe7Z0u9+6Lj/7aN/XP0j+dBk
M6VhATZXfk2Px/OtvekTczDpyTpqkK8AdKKa6dnF67MarkTV+Jk1h+JAYvt6DD1+EXLzUU/tQqP6
OQTZVMR4mg4AvuySLrl6J7Y6oYC8gIyIf1y3x5gT6sDr3nJjCuODJk1msfvBbxzJllaskt2weC5M
X4LBsonoC68MH2BHU5xgIxxuKM6VEVDJBTjYcYa2Bzrvu40tNyLmLWwWr2J5NfJ+hwC6NCDsIUVq
R6cuyNG63JMZh5aXdEYahRWPzA1sYgqtM8uPOcY0cz0gGSugtUUOYynYw1oNQwBBCnshQjpvoQ68
4aWtNNH0K9fU3h6WnP2hVU7ikSAOKSx/em2rtMQp5SjBSerZXEy0VtqbGMcM1ssWmlGFK9xYcQ4N
dAsSw38JN9SUCPRm+NZWWwDbSPeEoTG9nfORpkM1PjeiHZtRRx0Z9yWZP6N/rpKpVmZOBo926AQS
P5JNS2oLBS2iIfhm/B50btBQ7dKzOsFr3OKcKDRU3OJf/GxJB1oCVjGOQW2ydIUk7SJJp4vas7th
oVR1E0f9sBdt7TMw3HZNUPoWpEc46DKNboG0FxGhyr58H5DPmC2LN9kR/+UVX23CfmeQbFCHiGhg
Ogp44zKSXRJHq1E8ZXqHQd3/id6vILDtecG35lr5zxcsGM59TE5cRbDT2paOySUxpTUi/j0pUeaw
EQ21m4E6UqSQCMSWXacDlufd3XTHsUU01kpV2vGem/TE0eEEbVJjlJSlMVFI6qSjvzUhxEXrnNHN
WDw3GRS5Kr1T74yTnBD7hw3O7n0p+bIKSGFoDYFgx6WZ8ygEzVfbV5PApGfVMgeBcEhhFnINfTVl
kEZNHyrBO9Puc4rlBKwBc40MSZnvEIVIVZ+W8BGULtX25lrqgVCsqLzXHBBrtz+RNR0pGUyelpxA
s4W12ydqrrZ4wti+GO+vOyBReFiVXL7zL8/Zmf32OLliY4PDpLaT3j/el+iHryM1WxjzpQwJvaA2
vs5hzxpSTzHgfLid90hvg8yQe+zZEf4fTr1CYWw2SeBnX3rvJH/2fY28PiO1PMF98qZ+e19B35An
tthjbh/LscvKJMw9P/IfFWL5XZaGNRz2877TYPU2mqb7LvzSQZEroqyiFKOylHhVKD7tqkYsDKBl
zTBJbv3q4hwtsstaw7agCONemh5WJHD/TK88Y2fFKv2P7KdBaw9djLeghwjixo/z5Gq/8jlGRlU4
QHdthY3Hq8stlqDnFPqZcRQzNh22J55/yZQ92Ar4e5tS9iBRTy1GIIazXV+PGHB2Hb0hNweqcDAu
AHHfH+yOzGXRGLySXoBLeC+gNi5DV7O4aKFMKKhYGMAjnAhr3LpNU71BYtHfVFFvG0W+/KX2R1Ww
w2lVkq7D8uwKBZDGID7GStZls+FlsVZu43sMKQ9CGf2jeoQG0lFoRSNnsds5TCrsygQMVg3zakU4
H6vzVbaIvFwtejsVVglt9lHZkZ4jBRk59j5n6sA6e84Tn1VgPfnTzxMsn5Vzji5QZUctAZDUT8C9
etLixO01zOSnBSDSiQp+ZyHYsDfV+3aX8I5dX77+KDx/cHDvDQ+nV/s1nNCc0Tteszroq5yNmP9N
0gw2BbbDFaus5RmoLSpjXHcad++OZUQfcNcO+BqtCqmUR2aLAIqSej2MkYYH0Vm2ML2UiSRyenRr
iNdI1l1msj3SIIANfaGrHNmJs1fiP+CZTVk/LsAyHtdzwwLS7RNEtA+RsbXTiIULF7+5M0SqNvVD
JlWu2xqhCjADVvSy+x25gda19L58poskIpIvVtRLWdnLFojWfvwtpd6afdRy89y5UHMgkyc3V/is
Z+wFQ9SqO8LcHXYlZHjrQLxTE2klYY1HBjZuDbKrYRXllEPA8pWUMrMnqd+Tw4PhfxU/IiWCoM7z
cu69e5S2bhX8VkJo65UTDuAeX3GG866X6epcV0PZP2tKAr0ko5ZcJXuXbceipezmACpKzsji/wPp
G7eUkia1xsKnbeskGf/u36zXHY6+Jp6Sk8+Oxwx2/M829WOO/RsMLz6w/eooReKhgoLdvuPXijgv
RY9xbxmm2xmoXzi7QuJTWWkU4/1PYjPC8VqBJ9uXNHG3JQHV5hAYl+lML39K6fsY9ixe/fZ+0YuQ
LRLTQyJ8TQN11nj8617RfX/gSM9TwDODKf9255oAgso6ZkrTNljB9G8rI0n2Df57vBIMcs33aMXH
yNRTQ5yr18zlwoR+DmoX4Vd71eMir1jofVvXcpulKBaP/luJRHeuy5JIv3n+kkOA0SBXZKcg9rUd
7ExBdWwscsXOqwYYRSZvztqMopXYgQnWbCPnZvkZEwSmrf0bLgdcY9dB9K3CIab6YMYJOtRVRJv1
CUWbqktM0QSF1j/4uxW6naZy6jcfdMEFe5PAJjvbfOt/Po13zNmlIhaG1Kkr3utIdo9ZaUOIJhVg
bhYeqxmC2Jo3y6E5hLoek0gc0H+xiT4YhbW+GaXI5/6m+G1ACXsRIVfKSyek8EKEQSV/vDmzKWsR
dYatJMSUT8DWLXLaPIFjnGIS3N3m797QkqD+qzAne8oLtqHRgWFiISi7RChzNm/cThkFVpne4qyI
2DxVIZcdYyPF32WOBEf/HT8U3ta6e6VSLzr652MNML7e4aOstOK+veErniSjA8Fxwtx4hqssHRSF
2idk7d48qNZZZW69rgp037r/ckqtQRSZqKJJ7BxLyLcjF8it2oV/lWsv7d1LlXRBos/g1H4Uc06B
ZhQ9wQ069Pu93DPAAqKnIb6fzwT/1hnCWnWKGZMlgBPrlhTVI5wCDqcCm8/4tKK0LUglHTARy2JY
UYBOg1e+GyocG3n+mI6RaCGkeBC8o/bFtWvlYJ7xW5jiGeImLOzx4pfgDtqvpVOA1EwL8yAys6gJ
Qhl4KrEOALGISaULd99idKI2gQrwSVLRLWmfHnr8VEB2nPk2hreUIQoPFaEFLXnaD6HpYmdA0WbK
ai5MJOdaaCoYde4Jvcwegj3bE6iMwycWWxBIVcWU6HkF17Z5lbcRNnkG4vrKUb97+mBCexsF8dRx
BWU+tCtqda/iwUkaAsZxa1s2Isx8yzO6DgHDod3gzXX/S2ng8qWDwHn9V+sys4rqz7CAw4R1RD4F
zlIqOlWfpo9g/I6wn1d2mLTRqKlQxWwQFpL35wYS/V0LvCeFfFy3JcVlLto2opsKC/viGmn7HSCL
0MlfDcVnPexW0sgpz+zO5TP2Cyr2r6tZntwb+X6aJVtZFTeUYLPyw+NcobFXxzeAjpLKoSzfao0W
95nqGH2RLV2eJ0/4cWO3lORdOHS0NPgllSxin+F8lRAwTumaFc4L9v1Mb2/7URlBuK/WKOdwiAgV
23z1wI+4G1djy9E6HOWnV2JxuQDBDEcskjL89byWVbGsGitd0MTTOwN717AXT6QGxYnhpdQQi7Af
xjmro7MMbJ1yi7I1KnyHVclBlEa2FI4HR+EJBSuC/RQbAZKwjB47QFi69NX79wTc82+/wVfcbLZj
0ZzBLwyR9tbKSMNKnk5fiJChdsxSTr3ZOKuM2uyevb53HqZP1oz2LSSrTQ3hv3RVzVdciEuruEUV
0vCczOoMoW63DU9jGZDdAYEFoZ2SptVz6QgxVn+vJxm98ZMF54siYXCKUial7xoorRTMON/jmAMq
vJTIlN4Wvqp0wihWHA+DpXXaeMH22yDJiIjXxNJjoznBgANTJJbT7AjDTgwg/QizAUQJ5zDazaao
vcn8uGUNjd/ekCpvFjcaKEqXwPcgl2LU5E7QIbiFFVgrVcMj2nvzzkaHMI8M1qQW3+TfV0Qzmxba
hqGUtxcImduNzq8szO4uz8K5FOY3Bi4TJhXi1AhtfWEsYov9nLdMpzY5QIujuxVG7Ehuio418Dbo
w+s9CddzUKpgQ2pVAOH4q3AzzpXvM4i+kNOc54TVnSzH7zyOChlHu5W7jrleIusCuxUgBcJ/3Uqp
+PMu7n+LgfaklA7sKFeZp69ugiU6x9kTYpI6AI8lmTK0inNSK6BLkaFk2iUnZPcv7eg3LKxcCWfw
UxOT/m1uZI6pskTPWew5IGUFtyZKktw2D+2IIy836iVkAIruo6VZGvDgSLSYyOAnt8QBUnPmZV2U
RXEgrsatGntyquFa6YCYPTikI0k6YiB3PTA+YPrZnLLxQ+h+LSbHsbUUUs+LOFBN5/JZ/Pc0w4uM
sD0IWH7g/V/JqvI3lrlyiHcYzCI2I2JPh6y4kKObbQ7+gVHCKkHCfCHb6CWm/Sd7J/SUak1CSxuI
lPByHSq6oIJHeCE1rN5vyZfHCtRAghxN4zLTXR8y1sIcNdC1THXe3SASGiYBKW5/lbjjmo6d4BZm
4hTNzcrtTotXX9jMHjpqOb05BTjzpCO9ooR8gU8901DQ9kbNvV33ZWOk1AEqOSd0Xha9jOUdxM1w
0f6jWoyPraeldh6F0LiSRA7+fW3/WA/Vc94CRVZR+qrU2d1dga1qjRbcNakwE4Xqpiw/KkFIWJSQ
vY1r64E2GApL/nXv9xUV6RpOMjqExZbsZeKmZO/IZfUiFfI1JG23SGUG8+FNLA4AUkvGZuVKZUNU
LiKUTgQONn4nyPuk2YrV9HfB9obgaAvfx1iWKs+Jlgqim2aJT6E/Ui829gobVlPv624xCF72VBrJ
+BsfkgDz3DQg8pA4u0pApo2QLueDcDbCaxmeHMFg62pWkGVNO1Scp1yhL9TgIrILSjMGOR7h1ddz
5p2Nu0NoUNEdE0aTJkbOpfBM9+DHSR5B3ZEY9TkfomGHXRGj0QpoJI/Dxfmc51BtjDxUaoCJIZNa
2fCcYpOdUsXJW3K5oNlDU2oiARonRu17pwgLK09+49TOohAqrXb00Oq7Vik+N2JK42FQ8bhNGTeK
Trj9+UOyoG2gHwoBsqjKrtmdQf+f7LdSa+q0u28HdLK7r33iBHbiN8063ykLRFlVvG2HxXxA1r3l
IAhoU1vAGIUyU73MFFDesr7PDXSqJUwjoKL0zIP+g1tJc86FK4nJxuXRjqxiNQ6z8UIzs9TEp/Ky
sj25WcC2vseh90qFicCnWappFbTI/v9EWD1/zh4xf79HJzmrIsS1WEpxMfz1FcfU+CxWvCfAikFp
xiwzsw8aUogB8uOsGO6ll25UhEDL8oyypKVgI9Asyw1ZqHeLlqfYJi9G7oz/w5S+ZPvi6/PIzWNX
1M6L06/wsERhMM5tCftNBe/wYeiXVkcJfmQbT1MNkfNv7Bl8m35EnjhnamlIO+4cBRtupxHNgLJ2
HDz571fIptl0hjjJRaRAoUl/Yy0VbdB1RjE0o8THFEU1ssGkrKkqSvP1aL1FxPHNiwmIl6SFh/jP
H8GjZckk4GjVY6oKFrhX55CrkukrstGJNOyJr+of2E6PLm+ZCtvMuoi4AF8A6QoEz56nrwsTQy0U
Jk9Z0PoSRqBbXduS4zzoMRkvGENQslBcMqa8aKMPWyrNf69FV/W/n85poZO7Bjc6sgxr5/LDXg5g
uuhRAMNFJKLexvj76ezdGkS1pXmnC45VvJNWFXQCpj+HHgrXHrmu2KXtdsrJisCWKYegzF0unKr2
NfSPj1EFIO+Y88mwE8RZprynUoXWD54ixLba3PApj9PT2nAW+yn0E48Sp4wxMEZHLCdXGJsMosw0
ye1iMTdw3phQVNeIkT9/A+q5HWzrxmN5myoY/jeR9L1adaPoAG50Eh29j/YFaHqJqlG5ChyHYc7y
N7/eCq0rDqugNqjTHe2bEAOj5GnA0tMatPE3cRUAOAJkWNBtv4R3p3B4mAlpbjaroKEVnxb144Fk
w3LZRn9Y2l6D6LdNJlOZM09G/hhdywBEDfb/QO56TWrZ3YhJ0X9N5NjzG/LiCCI1FD6Nh7l/PoZa
DNlDgiGGoE3oP4sy3eIG49SZ+SjviHlLp59WcUe2a2XsJmYznhu52T5Ej6Qqa6k/De1VHSnrfXh9
9vK5/RIuhq5tAqydi7IdUQbaRLNGBESpkzpMvEC1ypu+TRSX96mprdOpK0yKhEgWEP3neEPSLLie
sQujWw7ssBrgysfx1d+kIIk1cSda3cND4v7jxV66romIIzafisn7o8QhMq6z8usNwG3sy1hi0OIi
O+LLma5o9lZnFV7nlcHwDwv2laKwnz6LgMUs9K5O8W8IzmbmKFfh8aPvDfYiRIzexLQWnaaEOuIy
5Sfr7PJxrvkERjHLkyyspPRa0qpSw2djQW6y1Uk5+uiDbCZirpeJXXBJaN04OqMVFr3WijhBdUcw
e5AZ0szYmHBUM/jGpT2hQo4E4Pze/dDQZWqBOIjgjg+g55RG4LLh5ZW/j48fJANJB/lzBQjR9k+n
u2Z0cqg57hbZJcXUtxOAKAOJ7O9xK2lMzaSVdMmQrPfNzDjKVoOWHz1xW6ADgi4lgmHMaiuMxMSU
/V9sh2yB0K+KzV1qMVa8OWqiZ0va5p5c5MIKSxb2vp/1T371Lb1TLVZMQFIh4wZr1uC8zIsHTjef
2bBitpLYcfuG41CZYwj0WR4YaoHzArhaSb+pBQlYKZMGFnj+jzJP1lbQ5FYT/BsHXPpZrXUKklNY
whJLKMiKept3sjn6d7MZHuWK0OlwN9DJYhDMf8/SxQ4OG+yF0y2fJ4W1Do6dBq5vukrttnLz1r94
IbHL6qfpQfPjlq81uTf5cVo/cy1kQy0ae0WZ5ejixQfwk1bJm4UR0j1kVIzgrr5KyBb2c5h6OLXm
AAIB6NicuTAVhAfLoXmhkMpqE7nTn8RDRBZQrimuOYG3GzbVJQ9Hf8RaPwVTWwi/6cEGsC13hvFK
3aMZI5O+HHii3BtbGH2iLPC0dCyoWvOenyUIdjLUOijttmIc7ePmWVd0eBNTHsaKnjYCDOcJo2+L
j2Gq0NUlpZWAauJWStouXKlhcWzW0uGEapdL6swp3NtOTxI+Fp+v6TIWu7ATl0Ilggaw93kJulwP
bPw9RF6qtXFCH6IhN1dUltV4XWzdSsSq3HwAzMVla7xi3VvdIWtta6DFo29Ji4UiEMfAlhfC6kbO
xy2Pfr5MuhbN9/58WFb0mOJzGh7+wWHpYLQy39mSgkDhMESRHyLpa/Go4ehGbN7jKJVgALn7zLNk
LBHU39cUnyl3JQw2IoXvXIOOofuKSjox0i9bFFKzHXEi0b1UUYd+nSyOg5OFzVbg1PeQQr11w4zu
YJeRdT5sNIAlHcJeshtNcZuMdNh3W9C+pU8xyBhz7eAVKKZhYsq0+hnr8kcAWh642t8KryWNaPTO
WYs3c76aso44+M3bf19HmvbbNstL2W/2fvnqDm/nwgQ9WdqvW4FKkrmldB00obF3j0n1+cBtkwO7
LZbvGIGcdFlb4ZdR66MRNlKW+XDPkoby1Uym9S1VuFMnoUo3oNBxn7bF2M81sunJ+ox35sA92Z/u
TzHNSHnw5w5X18dRTPcExifd9l4lg46boNOtNgyx94LVZsFP6AlGvn1tOizN5HqREQHWdkbGrB4c
gYy6uk69YdA7HJlWKwQxAZJWeeGVlIbc34p1TrhzB1AAUmzf3QMx6EU3oT+YJiz3/9nIOevfIH4u
Ks0knfBs853Ug+Luf6PUejZi5IKdFLBIrMZqUxzXlaGlzAWuhUEnBzWkEaV8PE+lfdXJ5N4BQKMD
AQ4AwU4/7yFX8emzzxjbmOZvPDFpKjFRRIMVVz6p/x5W9t9gEmurY4Yungzk/jFMLq29AFmUASPI
MPmeBym/ZOUlMuZKxyDQ5m/UZokc2MRVQHH90/TsYZlaXyzcsFWAyzwsDm4isYYKguQwBY4tT2GG
+d/EgsgV61VyTZvSBTXx1tjsXzHmoWeQiAy6fRMshQy/2wLv8x5Ptb+CKBfNE1ajxM+/d4K/2qi8
ZeFy82IIiXS75hT6ffj2b6fCigWi4oZKOYKm+IKcH0X1uv6gSxTtxVxfmNENhUxNmB11WYTW675D
VXPYzGJwNtlZXpN1L0jebe/J3TAtqMGzK34YFZtskWomaqXqlWQrLV+XDvJnU7UwhaR88ejHwHhP
SF75D+nuYSuLP7m2S/P2dv9VfEnIDTYCBsT5I/RtGbwEWmmpI72uk7gXA8V7oGGt8V5F/WELhjAU
WZeZatwwKdGAWQ4800MFtmVInETzLQc5uA/eUvs6rRB3FbyDFKMedwITD9WQjU55H18B1eXGjE8l
qwQ6s9Twz5OglSzwMd/SRDFmrMGIXQ8r/gYFfW3wSNNkvCZVXZg5RlNJGa6S3wa7zrOl8uGhskTZ
aNv6PKSUms+yCN4tkG7fazrwPULvW+IW+qSBVtFpZA4MY1KlZ6flpu7ip6R+3pm7hz9TOsxJkk8x
ieN6vi3SRdbEUvAujSjFlw7w5k+oiokEHFODd+rOyvGGQsI56A+ZOOIF+Fk3CmxqHssg2Oia4k2E
9hHCwAEyRDCvf3DUNjRuD41oq/ocbbfmlXPbFvgvc75rwfup2b3uCuUg6HlwQrkcof+TZSpfCp0A
ZZMWyD2HQRJyj2yW+A/UQYpQCdSSlwzhCg+jSi4JdauP3cwokAA0+2ANRvOLS/2b/yhL9QuvC0vn
2/SOEqji2OxHsElpyjsvMmBP8kzttaVv/mviNBoie7Ig22gUOOvzm3OhnVyM/0ecyAXLUlJDm1Ro
l9L7XsIdv25EbCl9pgtwu3L8Z3/6dQetYoL+Mz2lLjgLijgdT3edD/DyuzRUos5YS7MIbqDaCpHD
SyFiYHt+m6XtteUeRLEmUrnYx9EZ3Enk5aw1Mh1FTUAojKwua4cwHaSmdS6kgDnBcHhGf0Ojbg7c
3LlMBP3h4e34JeRfoIjr7T/Ow8Bu/ZXZFfndPRL6yrBx1eLW4vZqy712nnjRzZ2AaM5Ungr4OEJz
0PwX8H0mPcL9u6v+3y1eaJ41mQTBxWr/mUz4A1UwPHxXV6NtbABNWd+Q5PImdCWS77OiLbKl6gaQ
HT8gDoAQgagU5KCNmIVtTmAgomBFvCzJ6B/e4qsA+uOaQDzhUJ3yy5jgV234BjUuHEU2z3W4QucU
5raKGr/vwEqqDoK5meRxKhwNKSVlTt38ZsI4gLIPcDx2ftmHud4ARZlmW086mt1caCPzTpEG8RfC
sTGnjxMKV2ms4zw5EUgrbDJVrYXpdkpcX8t1N7BWMPbdbY6MdFbLynToA+07oDC2BWVEH0KDmJ5Z
UeayNkfuyMVNikGIB7+WsMkIehPFOC/HhiI8sw5EAqv70VPnClsoB5a6ywq+25PF78ujwXRZguga
0DtadKSTWWV/M6uCPHAER6MyWmtew2x0fvC0jS+mp7Q0mzowzPMhHjeT+WhwwSLT+RiTMzii6ugC
NZLiWd8Yv3r9iHEYj3T0J/9zIAyyrMSULer0WrDsffor/2wyWwlq2tDjdVAV8X+lmECZ+bWs29Lh
5vGvNKYhB6EE2bMoro6qtI/f8fksH5w6zbNVqLEgqrNNQaycKbry27jj+xzXwws47hkQT2N+Gmkb
CyAfqtRHIJxftYy3B39fKGCPgkrgvNHXiAH92I5Jgcf8GX9tN49SEZUbbQmizBDGmt9GcuSsDdBJ
fvsqknPxUPy0tMJAisVvGEBT66Cx8HxD9Efqz2nMg+9tkwsUhm53UyC6zWIVvG6vvrqGK7TyhCXX
jCcEge85V//i4NDXfD9HZo+xajIA/7dEvQ+O3oV4ci2dw9e5Z65T+5ln5o6PdokIDsCPF6IYJih5
tm2BrPAq59v9SKP3gv03hEfKpRhYjplO6CFVXEGhCm8Kv4W7NJzrln15LLvWVyd00XTLDkLk5YSp
r7NFUGkdCHQQF3Dulo8zJwvP60brfdglKXOixutqnSTlRBFnfn4LO3xD+bxXtmUBE/bIfiqkTSTs
u165WNrKztjm1BCymlzHEBfOFwfBxaQc7JBsjMyL8qc7k6kz9o0o/r/ICB3qxz2+0IUGh0Ga3i8Q
TLmYsJyf5jTx1b57ZxPv6XQJgD/GzzxRR1CKRbWY7qDVl38wgtZuvc6BEWAuayys2Pl5ukM7NE3/
SygCsGoPzmaPv2dDvMRSGkLuMCo6OCuU6pz6Pdd8ClZxCg/iWTdi7KF30YYdXIPx4v9Cdq3VDsiA
nDCYyAJ8JFcpXxqHK8haKvBsNb6tajriTW1bQ54eeV901xByAihhiqKFzF1fPiovkbT1ICcN/Zuf
4FDXAoGhiOdgr/YjDSWSWfjtY9ckhRHSK+u56Gz0keZ7Kt3Z+6bnVztlOj0XtirJIu/1soLNuc2u
ECs/Y9NtuCm5jzXT9qlAEAbkWoMsWV87PqY7aA41xGiNXJZczRGUyzLtVYd1AkJhj7HnOzSbTonU
Szqe/b7WnIVe5swoLD1Ly0QdZBYLlV7oKlVUOUHhS25OMd1wNMKiPCnviLNnghDNq7XdONYvD8J4
8Qsg53M/hmUZg+W8j92diAwP58qFhXPBSs3L4djKrKtOuHyCG0Ny7eJyHixdqesJAqN0NdwdkKhw
eno3RIyt3B6PWsAvWKXWGAlOS+VCEtATiLn2o4DO+OaWnuRyat3D/JH/yYHe+tgR9w9tJg3cuwmV
Hv/bSFzUO7EpvN5ZDJpa/+WrD6T89NZ4XR4h2l0GvH+5jUu7BAcaHduR07f2hF0Kyb5jWmUbMV7R
TQxBZpm9a4KQ4mJdGZzSjb1WId0FHPD3G2QJf83C39IlSF+2hMBZXIZFf3jmGTTnd8aMXd9HQGXF
0tJnHimARVZg8zsrE+ix+ibfily5xkTKdJ3VfSsHfB03BcaGy/s2XRnyvZsXrP68xE5Lyl2SNhl0
PAr7sDrwXgUTWWeonmpQuIiBchWC63SBJeGu+P55yuirqjQ1xhbS3NsXz9U2xkGR6PHwcTH+CgIB
BX/o6TSWlbn6y98AktUOX8AP1a2yzOx5OFf/zRJK+/IpemQTU4ftPOjf6Vv+HrSt53m2elyinMXe
eXpMTTwr+NxhU35z0sQhSnnccTzdtnztZOLMgF1C/UIgNzKt7osSvlTCnd+I+dCj6u7rx0B7NYqD
svL2JBF0fWYV46GD97n53S6vq0EBqftyzbmqN8W9zm6ByfgAf3ET8NKBhNuUBhluQrirVMdNp3Fm
yq0BdV6D2lc9wd0yxlfLqEs3hUrkVMlo+8DwNDjIdoRe07pNlkslx+/eEvzH/mLjkK2Jm2Gkloac
YZ9H1MyNMN7+uHDYBhawISCbwPPIGwAsjja7Daopu7FBKOsySteC0uU9kYwZuckTvdKnsAe/KTfN
1t6EocFOlSqgHDEPHNswO0ZvVKETp1A6yHsbTevd6CQb8hfdGRzUjrZNpbwlUH3WaAnLovLJZe6A
gTk16Sdk9ME5VqUQOjkR4+F3fcEZ8a2UYy0j9HDy4U+xWvHMtPICiPw0eeEU0K3KfINVf0ESRFdH
PRc2wPQ/dgZMguKDSFHJYjUwwH7ex1vE5XofRPgsvi/bNPLTI29w3UfSKhyRXnsEdokwHO8jdA+a
FtA37skfnRaCsS8qij+84Umsin9pKFtof/zCzz2a85PuUnoTjqoIcZYm9k/Q+WoH1zTVacZCTfLQ
HeSvxRVmSkjioSdwHNOVAFZstqwh6Dpiq7ijyj5upa+MHoVqtVK+QWcDmIfsA4BRrnbRx/sRAe1W
mr5XWLDjrfZy6rMSDi5u5BeW9V7RV9RmNlmQ7Ms4B8sCZahQG/pPzf9uSt2G61+pdbef5QinkgrU
YR7ut6GNJC/KJw2G0uu50HRmg8uvsTqGTiyHZvMM7BB2UisHJ/8iFdFuA3syKeNr+T6du0Z+HS1j
agSQOM0Q8f+30s2nKMTWNGP1l6YiMXT4QhNRJTKqUyo/5dKxhJ3BsAo08ZDKblm2qK1qOplabD/k
hm5qXVq8p7VxVi1qWxuLujiwlgw4yl7X/qYKzKLuYhF46GxuChmPZ/qfvSIGttyFFAboDJV34y0Q
ZDs0jjLnZbpv5cmQF5CPYMFokL0cDmSrS/IZOaQ9t23+m+Evc856y8gq91FHIZwYH3Jv1DgQkPRB
6HsG4EeVzpVt0n+l8hO3Ywf6e9fvFW1rs1bQm0U7xtEJu4Jar2d2cWmDU8W47QLbwFNImOirdGDq
KvZ5RiksYQiL7CbCcarkSJahr8aQ8zHvKZ/QXBWi+jrLb8I08MTGOkI0ISeQRoO8Zadx/zzk4V3P
yN0Xb0Sjubny+HsGDhwURt3/Ms+rosp5T84zSjVogxM+BqqPU4LMvjzVj4sWxc0fqEEkN8Lw0avR
jBGvyUBHrTVAJX2fX3JA75gopAvuDQpL8apMilcVtcnIlmElJz5xcmX60ku4OySlW0/Nu2MVAQNO
OuaLOlCmTj//9LnnhDzkPUXVCzdnt3qP/WSEeH9eSpBHILXzYrEL2zIWB3OPLZlOrTzeEcqBuu9S
8SAcAUtePEfTUC5YITCmBKcpt8noLG28ALhA/0QXhTwBUQQ1GQkQ/xIekdtZhGGkYKR2K8Uom7Fi
mwe548mDQVowYGhH5hMt0uzhGKGJehCOrOqvAQXEIm4O0XtuMwz9907R2lYbn8xPfi0pquf75pmR
2wEJUN2DVC96tCwj/9uCKN4B4Q5IFXewwmh19tZcm5kwUfXjCUxs0a8LLXUS1f8NLmTIqfcqGksx
GFtpayttj10SHPi5RHPhj9767JBFG2zvvR1K4yshCvycACxZLaZyMTcY5k5jLbsgdY4X1YLeVyiT
nZbKj6BqVOb/Zq+BiZiRJczyH1QSUEfbXHiLv7IYMx61hMn+r0QiyZemWMKNJ4m69q7RwsF1b+d7
AdnNDJkrBCZ6OGFGvCDRLj2U8XDLgQcRz6ibdyXjkvXEWH+1EfCI0TT7fmgJBHj+1PFe2qmS+0Cr
+ocD1eyc8ZvyTt01l88mYMGzeUSfpfguh6ClZj2TkOrdIHFoo/SVnGEBna4KY3VifZ7f65V2z2Zv
9KCDCiaeFFyadPd0AhKFDKyilU0mDbcaJ38ByiEQrlvYWlGHd69JPyhKMxHqvgUY8l4aIcZTrSVu
S3QJGJxCEi59gvDo3dlauwnBWgKZzzv849Cjs322Ch9YeIidP8UxZbmFaHnONYD1AozDvovHrOl9
M6oOw85ZZBFNrfkXJLf/InMjbjMyp5Ca3OIrlPOSndL17sz7/Tx2U0E9SSEiRb4/OWa1DMMfboDH
qcZ4jHTB3RheFFrF+2+Bc+mstsZRHaLhjgRJ08fpASRuxvLXQIMs/h5d2yDq99rJyjIMaW72a3Z1
+tawJ5CbBLQL2EsLfbt7JzrjgNl+zHFInFeRZMJIZ0gFHh3H9Dx6LShgUoOEjYvAHGMFdrzji33Z
okkvSdrnYBrh3gcY8z4W/ywa81FpQLOEHM1JNPxDUSJfrDYWFl9GM234aLS2RyVtMpEg/1zguytA
4hRNyIVngpGyKJjBhviKj0SNGrvwteh4Rm+PxxOIiQtC2dH3Ml4xOQsCsaluEMuMZ8p03KD5Ls46
dZZSlN//RR26bsbXsc9iYgE5EpZA0rKFOhx3Ic1DqZZZpssNYypBfvwLyM9HkHd2k8UPgzofb/Os
jR2Wqf9haVBTbicDHXOUBJIxbltDemEngrLONxqeSRDKxWLNywKOIbAuaFZ16iM1UCSRWMIvorsB
ynn2BCRe+ilF5xd01HgF0+txAUXdGU7wk4hblRJXHaJ6hSkLJlgOlKo4n+GneHsbZIVk13L7mXk7
7X5DMJ6h5q3vAQU3gxspOA/lfuTB1NzUUP+Ym8V962pXyAp23HklKj6Q5tVjYTL707h5xIBl7zYS
ertjlKBv/W7XdjuuptjCoBLsq93PR/VjZnNVByNCLbUoC7bJRD8dcL9YWXyAQXmDB7GdFJycjHx6
5DmNYbFgBYh0k4K8us2ccApbwJdVUFZkk9X+psfseWPa0mGdxVXnadWZGi8GsrRAlUKB7d4KKW8D
t2+7/qpBxxu83V/uroSMzPk0yqWdrtFi2W2WPaoPW3j2MSqrGAJxSTa2rzr8It0slN2bfuBXesIa
hPpuTzBvx+gW19RAlExxcpS8Gg9qvrODSmsP20HMU48lkDvZOv9A1NW7hED3XhRUOo3BbkAhWnXJ
Inxqhs6lGd80UfLKWl9wzXNJiBhBLzlDw/7vqoixV2EDIyqqT98FiS9P7W0TuHh+UzIIGKsphzAK
XpnfJFvFfRa2igQPfPYxMVL+e+bS6tohfuxe6AB2i+22MTgZH2R9cPN1V5s2y/iGS8yJQztojlJZ
rzTPlIZqaDPXfQi9QXLUofC9PHBTjaJvkcQu+YAfxZ63alomRlkIZ2Qxy+y8in5zj/FSDKkK5zDT
jHjlFogSQCiRwB/E/meQrwTLkbAIPwANWVpuboICgEVuK/LhiYiel27cQuHIDelO73cTnJHq4378
Lz4H0gy4EXVhZPy1yd+eO5ucgUSfja6kE5xsrzqr7HWGOWNM4rvurdn10kFpa7C8kdrZkFD/cZTi
lrnGYcLZCGdU+NrzVGXiBHi5R+sqrlwvpDbdfG2EwSuntTad2lgb6xbtjXhCQfJn9MjnBThVxOR1
RZ6H30t+BgsjaKXhx0LdNIX1rE3UHejUlmw/uMTF4cxbQ7jYk0b2CIc64j0nSLDyftnlKIx2qlQu
FQtMC1wUhVRdRpfDsqGdfn6rBOGwxM83KXBY0yzUUhrEv2pJXV2B7Kf5/ja2R1pG4oPoJuklh6AE
Ym4Imb7+7cIb7irwiqNTTURThFWK3mOfJit8R0s56Nwh9TtqyochBmxCA6+RegBym+2aHeCwBGn5
mnzQGbf0XYv8Gwj4zyii5EHNswQyxz751PUv6VfyxFP4FOz1DsZQlOU/deipkfhOA2DzWrIm/BZK
gRYPJ9FJZzkBRTwja6irL7akbxoWeDmFaW+/4d3l5rbOWOApg+F7dC5+IZ5y8R9TjP3JwGxSamHp
HvU7uKk5ZGUiDzExh5fXrlXuBHWasmLuzDg8cLuznpuuPqbx8KtHHsCAzAVbxRUEnKT0psLeeGKY
qIXxwda5mK34CXhDIoGOXBIYwH1QX8/uPNLxpmGAOqvdlN4vgWUFUE5tfxY2eXhq/qIp2EESHFQo
pbYkQmRFXv43mN3lMgWxQEXtjoWjtnxy00jp4mJ7ybvHr8fEN6HmWiURvi7v0dWQ8zMdPeNcd363
2uAv1ejBtoXiihjcqiDonUliVb/nEH+811NU/rSiddnDLw1FvaJ551EpjWzRr+BJnDbSq9bpEQ9O
XU3kT0O1Y2JZgqZK1x+HezraeNz2gDgIMFhpcebL1KJk3Ptdee23IU9fg8wUUNBJkETtlrVToIuk
AXwTt2Pa8QPElhl1bAJ61+t6gTgY9XNImG8DToW4JHQRtfYiIVpggKtD8Eq68d9BdzkQ/OwZEKvZ
I18mwmVcdR/EFBKNRsRsNPg08dB6YN3FfZgtcKFxQccCrafsOw4/RJvUGWoa0Gqfbk0fZGWurDVQ
dHcLl6T8fp5Z1P7MqZodL/oneUZOQLar9IW2a0kSozfM8ZipxoTSYn5iAIA8k/ABlBcp5zDlWszS
Yk5T68Ym/hDuxrjtyYxMO8Dp77ImSBDR/C2n1zDDQqD8W+yToE1iG4DT10mK2xYJ2e7MV8NF9kUS
h8Mf7d7TpLnqo956f5bq0Ygm5znSeiTujutFsmh2mPgGMYIaCg+mnF2wizffwQFLeQxML062Dybu
31R/AdYhxCXAmG6FwrYT2g2EX8HxCWAX6jD0uNXTqJ48dxdaCKeAsIeDywx4ex+u1AgB4qFIAzr8
bZmcsaAPJwQce7cgV7iS0pkocF2bdQOpm39RrGTvHcE1XPje77peY8WhnYbZGtSonEIzgHeUU2qO
7OoeQp6BzyB5ocU7T9ZP4ZBxrjJzKanB3jBFbz1Gj3B0kh/ggXtM2IJjW1yX/IMkbEyXdy8A4SnI
zuTdj6m2prGIlCmrSUbn9bf4xbIitCpp91HamiBOMfxqLb11NUWCCSRlF4N1VBZxiOe/mH8bXqVL
vfON2e/3P3bQkVqhPWocbfI/rigEPNMWu32uQJXzdK8gvaJ0zTnx7HD8mc5gzBoLgTjybjHoHwWv
LhOtwvWE0ijzx94DB6KCIcb996VDY1HiY2GnHg2ofEcGLPI5utZI1V1aWNNIG0xq8oZqoFroIAR8
bRTFDkf2kwWcwSnuZ/92txvvX2j6HnuKGDCPQw+puvD/YrMteTaZdNG64MzoAnyvzeVuFiSDiYtS
wgMe3ggLSgLVM5RwmS8Bwf9QpJI4HJ+2lbmHfvlR39CpQj5RW3WASO5biNiX8MGFY5fq2/31fnqv
LoMVR7MGP4Y0JgXLjVpgPpOMpkqJJ3oW3iIyfX23f3dRvALZPLjkMooUxqeUfddf2M6mofsOn12F
8EElqwik3Md4NdlIpYxHnm4NoDQ3M0/+L+b1Hx0w0id4ATdVyRwtZlcLRRRbOli3/bGUi5KxwGQO
LB8SaemOIOuFZx1oAfShYV9jm+QDFM49QOnYUUsFF9Uhp0LPbvKVXKgOmsp+FFzpZAVSejnzVqFL
nJCHtufTy6Q/PcdGFBP6DZnGZ7uWjXFjxdx186cxsjKXx+oY5o+f4l8+1+SVmnVp6FQT4EsuSGVE
lBEEK2rOnUp3ZJZckJGwFnO7L07751LBwNv2NfWpfDR+LYxfOKuuLarg955jghh4XgZfJHjAxX/R
0vat9SVdHCXV2QlT3T9mVmbJUDLW66sg1m+/JKy3LvxfYsIcydCUp5XFQVRZ7OTWL6ViRQuFTZtg
31aY5nhbuexCwA1t+SbUELFFSQ5SB7qtFT+bk2O51iNlOLujahB/2dxTtK7MjVf237gYoDJPunn+
BbcWOQMsv0pZwT62g4bKQ5tIk7I42T74ETLRvf6bxbt11Mr9I7fhxmvJVrMwLpEj2BFhAbVn24f2
tgaYym6O0ZBAfamfwVe1+hwpCR3mcmBQNGGrIUdG/9O0TY+sTWe4fIQzMb1kH8HfWS5sAVQzc+Hk
B6kcNzFrDlB7yrQa83n+ke+6u91e/xtquxrxRa2ZFzGsNUq1orO6bJ2iGMnXVSAtLiuWhdgnnnIM
WvxsWMGoMrVrFGSRckxszagIMflH9FeoYWP582doeaRLW8TJLB/hwTHUKW+9ZnC152R/BNTvh3U9
eHYXrzVQutxl3NnnN9o2dfSzEdT2z32I5MlA4xVJrs0OT711vEJDxwvtl4z9r/6cWe8cBfqlQ8fX
SsKOhYtxv4EAyDDQObJvAid/W+SlVQzcNudAmvNfTIisnKun+g/VQSHAtjkdhbjXeYL/2CoCe043
SIw36dLUSDwuus9JMhRyhsaNAigQdGCRVazpLtx6SUVpUqGGn0qmEZY8cMiKb1Gx/D42p4GuHOSV
2OPYdbb11kduNLdt2iVugSJLL2LgEhHVMCkppjc7m0qVz0Wqp+0PTYPwHj1ySGsenLaupBes+qBa
naiTwgw6rtGym9VooC3S4Nrq1Iw9DvPEmB0BMPWOQlkrlGn5SnaEUBeQwVCNCW6m+gCsDkmQQXyf
qJ7mAz9Rf8lALSijBwHLUAWvy7QcRpfLCO4jkTGYiUy2CwfjteZAqcqZas0gzM7GX8MeQLAbxYkA
yGj4z3zw1oTRNDA7+HGlSPoooyhsQ42phOh11LvB5L3IW2f4b6U3WNSvbsdzt6nmMZvpSfCN0mnk
EUk+s58VYE3Rm1uO13Su9BUhD8svyKMnkDzLyTEod8ZgmXrnOXzMcsirLANfzJyHpywRcW1uDc5Z
9QwJx8+LeMVAn/eBIgnoXHYPW6yg+lxG+tFjxmlF31qP5JZAb9czTK4OYbpisBaF6uNBr8B+tGHq
p0dFNP1zobnBFwyXLr4IKC0FjqTj0f1v6sVRwr7S5dORhIEvYvL/obVces+sjJoZKbpclDLoEd16
fQOMKR9XJsNwCmmmcD7RlNJFkJlwJgigd1f8WIWTp7kAKzt85U09wwIKURVRIMgBwZnz7u8XuIMT
qrrISkne8Y4B27YufOKsdUB8iKHD9jQSJ1iIhw4bfd+fXFUZ+HcSkEeU3j/mPuSII2Z0fEth58hq
Jf7lSVNzPaz8wWHimBEDn8HULxy7ydcwjVSJcbq2J6Ou3Nn+m6CBh9lpdFAaW+I44wTDl5V3kiaM
uIgQSMYUQeV5YTOzIRAzXyCKh9ZviGjhdN0ViskdxhyL4pV5HXlrAmuMJm/e2lxsPo6YLzUgOAuK
LL+c2+08AM4j4u37Gps9i2DZQI10y31snv4m1JdPxpp6DgPdWuf3CYbxOMabd6cZtNyOD8oNn6ad
Bsf07YzTgaxMicov43sqhDwDK0lacDrtSKq6QWQaTleJcLFgwnuo+VzVNQKeLKWIRrRcEoIxJVWU
WPvU6Syl3eOMcr95HYJEaN+Qq5sN0ojUzEs4HGb86ulUzRfndK98qR0j13i7pMrSDVgMHjFv/CqR
w4p1Zaej0x4LniMc19ce3KbWIBn+X92X0ev1jJySf31UfsmJhvSuWWawib2UxRDy5vYDvLIFcFA2
IFuY/FadUZy7xyrvCNTd+FAuS+DoeFceU61T8tf76edr2OeBQpVioQxcCLoYrbEdn9NxsvXL+XDx
/q8PQAQAi+dckDY6wDAk3Is7uCAhNFoSChMfByeK6xwjNuc97AkE94oiZ0krvzvjUyLVCijgjh0j
/+9dVjZ75zOdpYLfplG4IIkqcHIyMnq7iYBQHufQCUdKQdjkYwODDAfNSxs95djLzRUrJEoFesGF
beFjAESJ5hPY9xK+zd+gPbAJi3slqmvAZvUIJgmkgOvvtG6LBI/ezFW9P18icaWBajrXqsFTg6kt
AmY9MrzVEi7Dh/K/kkpu0p8Qd30WaK5/w6kIPDaY7Ty64LG3lJnThmP7XVVmLQYNBI8sTYGIQrrY
tf5Rp5Fv2Nv1A/FuibYtIoArDgF2p9n2djZJ65GQvKoX3nev7zNPbvgCfCJG5BQ0DZkNs7zlwtXZ
jRAC0sIx40XCqJ5vnbKte2ZvoiYTLP3o6SLQO7JVLEq2S35KxbjvE4JxFvCjqJBNROmaa1CqtFIJ
Cw4UakjTwlZblSJNFsb0wIJ+V0ETFVEi47MmMKQz/+I25FW02iS+SPgm4FKO6BtcTkQPs9w0ALV6
TsMk1m/6RrNm+9xQ1SPmL95kI/hrs0bIyPmxrUu3/2xel7VnovqqqvbqPG3OmhMcjZGN4QKKKic4
ZVM+O2tF0k5xFXjgwFa87gsLtxNz3BJnYPwC8dzJprPHsP8M2YmVvd+tvY8Y4TqrzMDPAkswOT+U
giz6iQ6P+stIf4phxYo024IYj5owu8qQ3O+w3DWvra7PWR6fxPwlVasf1n6LdqFQjWZNzGm3i9Bz
LZBXvssOKB2mRCIyY6YTDam2lo3+w6N5RVM44WlhKpg0f1rZDC1f8G2Ucjxx8Lx3LUe8/8PZ20+s
8j601ZWitTl14TaIolcHZOtwbSfCQszyFDyORe69aF5T5vUrMvxXbsELTc4pVJ2eYndqzI1sUEcR
J3K0a2T1XLMUj6Ft78bviZDCCqh/pgLmf3i2gNZlJt/kFUZQGlD6tBa9d3ueKm16q6yBnoph5/SV
FJVG23SfqAXg0hzYtnS5zEPfPshIJz1v2NwQfeV0bdCoLIQ2TuUMqRkCRWxK+V3MD444p9QwGt79
SmSmNc+yE/x6p1zqfavuEiWPGfEoQnPPQDKMFaeKiCb0U1vTtMKj3WcCgyNTAGRO6jB4o0DJUAdv
IG3OWc9HFYe0vTKMXn+Ly8mEyfjJjFZgWG1uvHPROsni1O6lpfvLBLG5fRywdEbJ1dDctFyUCVLx
3T2jWfgK8fT8DN2hz+jsSd2kA130uray4X2SVoPO6TKAWsZySfujxwWnlgWq01KVenek5XD2ekBZ
iE/feCWyEByLgq/01JK3QcBQzDWxcCLQ4UTTR6K/u7QkLa8VRD5hXIio5pKDPGtRmK5ZXqMdbLGa
JSr5yc3YGRh09CXJ0RB02jsvLtXB/Cb9hkKgQuJI8aQuWvihMGecZsqxr0+MQHDgp+d0nAOSNylg
K2tIMHel/eswZPv0XzTAHZMaUsTx+YdhMWhW6eeX3sDbGLTnzrkBs9/OdVYdAFO32LCNdw5xMcaG
UqLLn5jjLm046mEamdZI9jNcgdZOnjEQ8ycAhEfBkYbJ1ajwsATOm7nLXpkyIlkJsH7TUn1PVrcR
lGH+Mg1FLwAyUUsqHFTgEPq+RmvdAnnaQPNVZ3gBKoRWIa15jngQS6c5j9fL9z9ebtO7sgG0Ha1b
hauY3xv1Pco86ilwWVeOqVTKynWkwpbAwRu4ws1dAEh8L5gsJKwdlY7BmhNoLH8XavGSy0SEaKvT
dUJkPfPUJ7eFNBnZxpssJwlsx//EkX+j4p+s7tSoagexfyOTLXNNQavk++5fLtxTLpT4y78Sljo6
dvcYBcTVwOVSs/oyizR2saejIhUSPlab/iUFvHG1CCVXVRch/9VZfH5JImg4nBd0+ri3o3a6zLNl
3Gud1UYD4wtPW+Bu8+5LVSSXBQUNDSoXk6IjsEq7Mb+7V7RSvmZ9XVyxeRjqXWAdkrRaOs8GDBKk
Q62FSzvH5S3qpRK4WIMR8Nt5xNzwZdVhDzP4E0KbjTKxondRqyol8HBM84i+2pBd2AeXpyMlHI8y
dR0nZRBcQ5AIBaddG7Q+osDGYI/kp2AiH9YkvKyeXtTZdFqbI+pTCYcxOjJ3EUdWaN5SsjkHsO/h
5Bk/oVl4K8/+Hoo9bgSf6ILwB7YmlzWbXI+i8dgTemZfFA/4GrkhYnI2Lw4a91qc/zwcHZTI6Oal
5HEncyXdG2/dPKKqJwONrKkpeqZ+0VjrYyOD7E9PN7viFTrihBMPPYI7uwQpG1RbGl6fVmq5YcXN
9+X6sd0mPjmRRXSx3jLQIen/77nD/wTiCSBjTANKd0gWPXGXpvSpq4PPVYnKRiTo2wk6xEW+O59w
p88VagzNqpFL6KJmXjkx6v4EN9qrwQX3xZ0YAEldOLFeUgLTeHrdV3sRlVFZi0IbxqFMH5OTijQt
E/h+icaRA076d2OftCEhb2yUg2+x0GYkSYyZG6WVbOq1XyQGBHClWvt2ryJ9VeHTrJ7HIUBbRq83
I/MEqyZoz8SAzTmS5vXWYXvBwW/z8ORz4BsLqCNAEtpVGyGNib0V0mQZyHs4EmYxXYURyVLR11IQ
gycH72pCRnq/YsnxFK/sEqu+jomHJSmX6byAz4lrF0gBpZ4wredTQKenP/ftj1P2F8sOePrdXE/w
z14Zc25MWMeSM0dfb2ixc/pAZ2PpA0XjmgPV9TV37NQg8gunBRfGGq4gj+VE3e8dwvYucD3wwubg
RKl0e6ZqixeGRKMwQbRvAudqWrH31vaxK15zQAk4XCdzKZvMCfTsKm+hLO6IaLpw8vQDjKzSRvCw
5YBoZ/3v9o883Dj+HFmNDqWtUQycLPtHqxPEkBQpPqjmNpoFqN8fs9GmWqtk+YnRpWNKxwNlDebz
3WZSyIwekjrLzTHeBX4ms/ZXMRcnPFnFd34c878wys+1QW7MPVIymwCkuI7QSCI6d5JW0/2zt+Po
+0N3bSop9ItAFDXqu8OBmBx39SBrz9/GOLn05EdG5ZCdVu7/fyiUQGtctk57o1Xh24E9qpJ1CGKQ
bEREpMLyqSWmQEhd270ZsM6Jtn0FfUWr+0UUr2VacLlSJJBWz/LkoJ0GLGIi0kh0Op7QHWA4Kl18
LXW/wMdkCkyTbgrVPU8YtEWcMWsvSdRi6uAvDdLMd/eSxasjEjEVCXFiMzZy1KzRdCYBjPCAeYuQ
4VdX8kg0BTq7UiwObymTdEDpfBcf19xMPLWktnYQD1HuTpBeA8zUATtXfWUz6nTpd5AJ4aQyaSxI
7YJ1CHVEeRHVt26aG7VSxNhLGPn6upjrZ4ga3W7Fo9KbUXPAxoF3xiG4hgmfujaAPea6cJIaxm5j
dx2lK9qOT6kx9S/NyedcCKB3zUTYhB6d+JVqU+Kedh8Hd6PSzyfTCK0uGf24ffKL+HJ41vOBVA7p
fPWePZ9eAaGJS8yBRShmllpPKTBLXwAV5CTGiRS/4zmixSTyRKo3JFJBX0KLuxZc3mjnFesnCig+
G6J9Xzqg8JSxlQuwL2KdThrBQIv45T/vZpBNHA9QszeGB0kVKrohw3IzmsMOmAtD0LPOE1FFO4IO
6H465xETHaI+cIFb0Y9KQPw0/A/fCBNN8cKGeOdj9cauXhQYzJgNTdFTAFW+lyJXgb7Vxlrb6X7h
mabLOkceTtB56viGgoOtbAZt/9elKskWI1auG04Sx+udIk2G1Jze1359M+WSRAeDkH/0y/omnknQ
FkXDQaDGEqMpQ9UHxpkV1Abh91pYawkv39w3R3pdBxqI+DSrr8BOBdWisBLPGGHTungEJW1F754o
Fy8gd57ZTjpdV8/XZdzv+w5Eog6BkC+l8XXtHOSuJ/98XJZQ85OQSdaVuFqBsaScPpOuHEGjEzUu
kq75KTYJ99CJX1jSrh/VPTyX1IBtkzc7iiW16jnHf7jn/DAa2o3Yv1GcOCKeUaOfIJdHQEAa2sV/
Tz7w7rDOmSGPS7bLOM1P2J6T9ve/JtkULcFFmH3BmcHery9IZOeB97kKZGKdb9bhFaxSNS/pf1MA
WTrRK2qmUu2Yo4VIoV1ltAa9UMHv6VjOM8gEirWF6wTPMIw7NoFVkP/cPYtc69gc/6SiycwQu0q6
K0CsynhIzQpfCzVp5G/c+VApu562YXKZ57snnX+4rlm4gYE01YYhVLKbIqWgLwB6Kg6fCJdCWXzT
woBFzIvbAMcYDf5/A3phpAm6B7npLMkwSGodDBbamircpaj7FzrrWqbXV/KuVEIxCeOYDS8de018
6HD4oKt+BVBDxF8w39T1letvWE+4efbz+T/fZjtQZpwzQxNcQEqA4RS4F7rBAQgISGxJXlf3tmnp
GnPuEd+EZBL6Dz4iGaH124gfKcK4lLAeDLVDBBl+QyE7j3kQFLk2aK2x3Ml6iFy1psBrQFhUsxv2
kjUx6jLN7c2/zT41hpjxZjsBBfRGHI5mxZIJxigkUmx0T/NAp2MSlZ0pQfRRr/LOpZWE8BaL8NOf
qD+D1caAMDZCYSi6OxusHqwP2IVVAeVb5OxzZ4ISeMCly730Ya9rpTU9uYUOKGUE9x8oDlyVyaAK
F6GXH9LhCIbJy9huuX7trldqA/Sx1PQwq3zXcbyWebW20KpsZDpxlvd3LWaT9EIv7szwVjpe2ayT
eCw9effOFAoxindpq50WtoMj8OVcy3WwMDm6B0BOuzcn8x1lP9ZFEPJbmF3IwAAaPZvvgnXPCofm
BpeI/oaas7+WysWNxjpKns2nXBx7LAR+f8wKFiJNw0IZftHdtJ1VeFWc2sOVXAtbfXS1F44s8atJ
H1tKeRUwRrxmFXQ29dZ5DbcuqbWst4p51hBlIytfvBZJXx2Smjfn1KrBQOcngYmwl9YLT3KPEV9Y
YyliaRwiFEVYq85XFiqqlT9Mnr4OfrXc5JzemwrakjvkNGtXUgx4lYKfovNC5OtgQQ5h1gNrX+6T
v4Viqew0NKUC10gcRRD5Stgtv2yUE5Z7If1LejqlKeE4gm7AGly7dp6m0BGrX+Qgo+0paw8XgA+c
Yr/Q+Wg2aMMqURTVk0cgRG1ZKVFoFGv6vhxKkwC0jh+a02jBzbqg/vgacb0UNDynwK1xGw609nS2
7mzODR4MsjVaL6vSgeCvN4/C+/R3zqrl9V+m3AuIa7OD6RTi8Gs/sb58PIuXV1AfaHVGNQLJidg2
hHaTm4sv3dLAYz/ZyYKZuIUbQAf0SJCC6Azu3lGxcMsGyWYRKuMbWX0bcRBCHK7Kz+hVM97KdMUf
dZ1JBs1quQs6+l07FBJEt0V9LoMEeWUNF/N7Av9SYqr7R5+7yhuRU6iR4YGV7I6RwwVghZo5SA7Z
KoSAnaYBm/0nNVfX23r38mb7yfDB9+IBKeb0zR2FloslJnzdQJB9pINpPlTsEJEOB0pDfEOL1LA6
MhWiF2l7TPHg+N5/HmxugV37xV8si9f4bjWcQ3NDYQrm3BJk+idpZSyHU/YAHK2UtN9Qh+VVl4VX
7DM3rc4ZC1JjUhZNMxR/0PehXkVaAn4MXvLcBZrv5KWBhLaxoXUMb6vMYFcVKTFkwpywKk7/P+oC
LDDX741uXMH/IofW/VqModDLaU3KdBiciRY69l7k7PgrLaZV06uM+HUUsdjH8MPciupBP+86pxZq
JCLDVCnSLiDTN10uJukI3tz7NY8nlVTELPjgEBKCam3UUEMs8fxCRhAO6twLRW7PVVVadftHS94d
km4q/WyMZDehEKSz3G8Bu1vIoCLaJeFY2DudBEPqyFzOOpNDirrJHoXsEMp3gjY8rnhEUfKdls2a
WwtIu+tS59sONWiBhKsnupiyj9H0zMcwZ8BmiBzJt/MXvhWl2S5fjKyHlFza3xyesnkqBliM7uk3
ENi/LrRA5NtYJzeCyVTvhAQyYovN7GtYWGR/ICPknK1wVaTMkBJ0802ZvVGYWrSrlw8Tk1DDQIED
x7u25sgOxP6Akux4vNUCl4R6KnAstLd2BTWxH4WMM2LhlBBdUsma8TnYwHcKPwTxCzQXJ3+r+U1p
tXisIN7Y+O8tzoJ1NF5VfgUtZeVpIK5aTpJFXYHjzZ4aFtz9bGM+6Q7Qg+U+marDc347TmjLHjwb
/UqaUGroUgi0jtNQCLjJ5pAfCBxpHqepL1chLu0yjJtpI5EOnrzsaW5TBNu0AHRrx00O0OQi4144
Z/nfSCUY91JB+jA9D3vTfwbJh1jRu1FExm/Kz68nAr2xnWdCPL+c4ToIW9zOn1f8DpvzMkaX4Zdk
6A6QrWf+tbf1uwX2sSfc0hw5i8ntilTeQmwRIsDGPqHd/aVhhKXYM/5fKjFkB/QUKy6uWETohabo
2MSpKmn3QMrxJ9PtHrXlz5P/DJmJzD3OFhX2MOW1m30iQPvpi2O19VSJ2tiw4N9x55QyYntqExMe
fVFisVwUP0ARi0y7W81zh2z3jTmt6msVXPOw/27Zl+9K/kWDWxYq3Q9wQX9l+CVTl4jEREiYT6h4
IGNBRfV6v+Ixz5upTVDdewgFBeoaNFXU3c3bp0fBQzqZBENTsqlYMLGiuJGVjHLGNSWba0IDxyY8
aGTcu13jcM0qzcmVGRFcLnUTxQsSjJUzwmj4Nk7AUBpIIpj0Cz/IXUALj0zoPZBBW3SAiLTNC7JX
IqYDmBwk43roTo51j1kwSppguUrgTKC/Vr9U5+/epJLk9lYAeT3qG00hFvQz15vgyDQzEqlVf718
C9ICwrE3yaEsgHDWkfaKlk6IJxpfo0Y/aBuShnvnZF1UYp5pDSStcwFyPXzoDFwnCD1KUx5XMkZF
ZcDZA/mGkQ+78gg+yR6AOeyHmK9UuBy2jWWTmJAzGjhYc8fd9djL/5V4uWWmjRVsQhggJaYg8jQw
rWhxUEbyzIBksNVZ2PUPwqFznBfjnn9lRrqWVqQfZNwIjsHLHLxut+I3RjGXMfwroFXLo0oWj1CO
PfJZCNsDqN1aJRQaa///T7GeDavkFZeUMq4RIVAuyfu8VaWhjFteJEIRFY16seEKG95TG0DbvQkD
fPQAbvi8PB412z0gQ1s7BHdRPSy17uJxfBHX/zxNXkWz8xUzFL08+95lTz/qnNCp9QCGAAqGv+Bv
lXcIPdG0Sn3/kNP7LFX82u/sifrhZjZUD7Y9rUa/HjrJi+vdxz+Ob7Owt8fJErpRR3CTaBrxO2wB
SsR6cgC/hCMUxc0xD0nYJCTWZu+OENEV9eRYiud9D6FEh8AGuk71ZypQz1ysZ6hyyncRFhM0vMxY
WfhPFe78tFNZQjolPePOE8vNLfAWcjwKrS13sr8W4AqZf3BMbRoMx29Ehm7WiZ4ze4QZWeZOFVqy
VmeO3O4DKSQsq/FHvnL529pZ2kPzQpOAewwt+fLjws3RvCqGcIQsRX8spOnbsMKMLKU1OqnQbMyP
0wxxneASENhyPu7VIfYZGzXregRna+b77YPdMLObDVsNxXeSoIK/zG+NsGDPpEnB+Cc1yc/pr154
f1e+dfmIHFESgCnE0+oTBXtR+hM6Q75M1NuF04rHw5qp/QMRNbCvbihM48O2i04iVimbDfUD4+Ht
7AL8kUWkzhQXg06a3MhW1T1dnWXh96KhwGGWfecXF4KyHixd7sRUmU+aatkOU9qtaBJ6yZ3yRCvi
fcBQry6DPLaG/0XMlJkJBiCNiZymKONlbB2kQ5dtuxAHBZ2cT4HFPCjMY1pbLenUu0nEVd33iETg
Zgu6cxKc8+I0wJk38UlTdOuB58eIyWqbuGWwvcJrBSKh0xxCRn49vZ8LDwEXSB6t2zETBF331TRx
qb7Y5KjHqmgZDjjMitsTsG5e6QyOE6L2tOrCrAwv5lx5L/cagSKFUgWdfPnFMvELykd8lEGq0UT3
rqmfUy4oOR2tv3ZPriDuQrMyeUB0Tq5nLm3JxzbzmUGB36T7UrhBUAgLYFu8zb2kmKToEiNs1mbP
CVvIW7fRdbT+S6+cwNtuViZlRz6I86y2lnhgEiFHF0URgiOqQUi+kdlNywAusPGBOktzNSHRb8uz
TjMqCochMAaNK+hmeqwKFhRt7Lp3VcsGAq0v+0tVHdPn6P59IkgjEEakIFXC6v2sRTK8dXaBhHXO
12KPwreUIlYiBRRA2OduwSz1msZjYTm3fMQCdoQL+SMGfmBmd2HyxbCLEN+3RDGQgF619wcZ7mhF
tAxooVx/KGTw+pnOIfHNiOvLnkq3A/oVZVa0VHj7XY2MdFs204PShyr7rsoRU6/723CHG7P0hQ5s
UtMa1n0c41rdoMdWP8zRzoIdHo4r9NZhT/thMCW0GY1lmGvtbuLgbaUCrXrctisiNfZGsrzFPMoX
SWvYBl9f3uEW4GXZx9Um9SjjrGMbT7yH+dvYcitWGWxknWJdqMzBL3wZhaaFlK0Zn4ty9V8vR5GX
GIxZNjJPzOB0xzqQH2ObW7I6wqdOnjAwcad2izNS9KPosLcjd+BlaejpvkQiOdQ1GCLLU0LAw9H3
K4RxKvW7U16UndV4NYnUzXM/i9R0VcTIvzOcn0YrB6nwu08ZEKQXuKbQXjgWz5nUgXn1dstoo6CU
Fr2tKJeZ6GwVlmxEiyR8z291Lkmg3jBUjD8okev1/o1TgbBQOx0k7r15ZtY4SIg+WhEJlviWlJf3
KLV476/5D4VCfnl9PC8TFsrws29h4S3O3o4Pn8560a5RFDlk6OMAEIQ2mn4j7EWohT0BW+PVAOSI
6qVUfkaJY8Fys+PrYOuXVc+RrvO9GRJx+E2ARWKQ+J3MYMPy3kbFfuUo5/ulQOxLJgEvShpQ/hdo
oZgZgnz4BE+TzFeqsdO7cTig6DYZTiAYueqbrjkogTmW59m4CE7UR1K8exxyu8MhGHsYt79eB+Q7
e8UletojcxdvvRnJo3r5/b74HfryQXqDlpWxy9vhTNB7ioy13Bz3HBJD6LStY4w6zBa4mfCH1JX2
k93yzcL9smaaod99xdkSJ+MietCWwNdUni55ianHnPzUTOTjfkyL0yDvRTWl6LIFIcG4A3lRrYM/
7lX6y7hvrERfUdmgaFTQvVzYjvV5PLgTorpWFSZ2IxwrFY+LttkOfphOE/SevALE7xw3XviyqXjo
TgBakR6nueQya67rQl1jeJy1+/gfc5DI06YTPLMYMptLBJEs+sw+b58fENq32PwaSD7qHptkuro0
RuHmpLr4F6lvrlZK72JgYLU8x5Q0oBtwGjbw7hCAotTIKfNfCgdgXHMM2yhnC1JMBmLr1/4tAdX/
3a+4Oe/+TAsQcjBXHmFybSqMrNxVhXvobVTa/v+Sf1zPtbA+4uXbj1nbzAUIIyUl0+yaMeSshn0l
qDmxd4cpeFxH4rlzrRLDwSgfz5rHaP43Unc5cjgYM181MUYihdjMPQjQxUEKkb+lYEh7DAS9/5Q8
uCn7/SkMV59iQCIolryIM1E4lk75eo404a6omfjHQf6cO5mANpdGvCG43Jd/QjZ9ULFxF5spHnn4
6oOF0VsqiNAoVE5Ns6bcICLYrMn4W1pH1YEj+BYJeCE138kLEQNkxT9ZwJ6mF24suSwlqcl4Skij
z4h7T1Lht6J6EqevTsPv/rKqTsY6v35m8tlIq9PEhuY1pWbMwqWaFweAJa2gsYjr8JZV4iEniwM9
wC9PRmIdnXF6BGYiRsH2PG+S6jiOj5yQhhlNP8b9VrsM9RmU1WKTvGDcL71fqPkUee9sTpR+ocH5
RiK5zPh7iRwMZt+VJ6i50wY/ZXpSoWvi1T9ORwCTKkvSqa8su1E/kMPUz+5tsIFqqkc3KC6cDVLJ
KLlHlzb/IJGcdha4AvgzkDeDEPyenhOwmdT26NFB0KrxwhV6PdBPfIFAnWGWHTGL5jXQvZIHdAWP
07aQ0j8s6WsleOQkaqzUGZfPsaWzouceTW+pnp+xis4oaTAKAtmrh40oOt3+bRwopz33bWYPhaft
CnD3SZiGcwStpkYUGJ1gR4RgZT3PrBBfHLOv/V7aBZubAmgV5OXnTSs5gD6Q9jNixyn7Aw0l1USV
k5e2JI/yMxpdBarY5PQP+Bku1UFQhblWMx/AbUyw0t2NNxdetMaTXH1WieXYzQLQ+EXXHOzi9vNy
vkWSC7wNKOVzP+++cqDExCkYwY8kyZnglS39cQujSlzg9Wj5nGjOf8/YNrI0/g2zfjm0kXXV0RLY
TFSnz9vWquYGgpJaqtsKF6Yev+TPRj1HX7a0Q8as4Oi3IsLmKywtTQdiSaLwQAdNkt6TzW9uQLFz
E3/Rd+ECEOAFDKq5vx8TzHJ05XmH+irrFBm9TPrxYdzIXdq2NsoV4eALJTJyvp89DUldr6i3d+bZ
gB3TpW2RnEZq/4iq7KaI7RLKqrteEu6IWEKrbsv9tPQgfqUFXU6MoUIa3vHOO4SX/3FgU0Swsdbb
eByWgnfQRP1nhhsE/NXEhZXceGNKYlRXls3QTFHkoN7G0bh1e8r9T1Gn/TMxmHfMyp0uRa7anHAS
QJANfRWQ4b2Zh8q69EftlS5Gm43bVwAHGYYDqH/POxDIKvzKPWUUoF8dEJsXzARD7V4N36HjLtI3
woXugXPhJkPoho9sh7Tvf72dGz89NShyBZ3ZesnEb8p48PzceEdXIAhyyYc6NMnr29AOl0y6YyFM
9/jzN1Nu9qqsuHm1NAK6dLzH1+BrAloer9/toLlNm86e4QOaqKhqIEP0taZ7aMESKFpkPzlO2U65
O5VXbuBFf4Hn0yyp4ONC3ZVRV2o/tzWROfhMxDPOVxOC66wMoGtrAQxj/zu+w9NghodlsO6HW2Oo
m2QbLjug2cqC4VzlylcQitOb+iqjVIc+hiUebRoAtsmiHvd0V04KF7omG/0FJXQnNQe0gzeafZL0
QAEfXMtG0jxHHxkHpYfju6gCEYz7QgFPYhIZY0Beff/570KLWeo362mHx0rDvUCEuHdBSYFCIais
AAKbT/zmPIWpNL2z1Jd2v0zuu/lna+PgT9KeW8+yMCbERiLB9+IHyDYa2g572NwLFyV1k+gaagfL
Iyn6ZKcpfIiRKTbuCEvUx86caGLsKWBw5t8F9JWePfGGAu0Offd2m0q3OsCIEKRkMH1frSSTYieC
HDbGFZeBHSWz1NkmUc7XbglIXRA9n2XEid7GjkmZGJMlyR/jjqpANSQ93VLmKXIYl0PP4HiY2OF8
EtDqigbOrCD7K8Kd2uwWPsKzE6poPN1Y6WjhZ9MscE3O4pU4K/Xi+41sP4egP4hGICklHvqBqfwy
5hMRpk0llCdzHJCLi8qkQFtFb2bDZgB83F5FQc6v8YtMThmCslt43TAjFaLBaLoADO+FQGFHPF5Q
8RYWmjml+K3TmqOj6FNQs8QxtVodr3AlTUvOujiTYOM+0S9+Rgh/z0DAAcVdGxJ2K3uJ6M7wK2+K
cQvdwKIKbg0dwaya00neCl62G4uCXAj+eLGyKgbZmSw6gyQi+VkF2aKqX+O9b4J/CLQHNtgdSSzT
UOG4uSkOnK4STafhRSGwTV1If7/a47tyrHTtNwNCrVO9cEnxgngkAyRcT83J/We4HcyzDdzvqcbb
v0bA5hJcfVvTL7L/IZGMPfMndcUfwXb7qyM5RNpzBkiDbdvJ47B2bijqs6hNH3+mvHBOlU60ysuw
i6ZLpdcaLY+mHrb0o083hyrP35TD5lZ6U0KBqh8s40LHQqAZZwx0zkFwx+2SRbgoy+Kyg0rzN1HM
1t3FpJyaUuLSDqatGW+GbKrOImSFYzwrjA693BRO9xj4HJZxmyoINbqHG2Eozy2AzqPhwK/OwB8x
vB25reb57MCjeQ1BHyl6pxcSeRc+Q8A4ao9/BTJcQu4D+Rs13uDGf3RUSH5GqOc/HJ1KD9JpLzuJ
/YYgl8qLYHzJZ//8jj1tUeK5Svt18TKkFuqVu5LIsBemkY704beIzzau6ulzPwrbKJoqjHacrRVZ
gMkDTkKtfUqFithCTgzJ53fTUi6Qx5lTVtW2emHoiqGYfWy/z63wX5gTpYykLOQxT5YapkbxI2fZ
7+MMf4fFgIhNgduF4CANGh08YMa9k1uqhw951VVxlQXjouG0Y73U09rYLGXEyN+pz+WECwbB38Ig
Nar5lIiqRX3z2KhkYT2sDLnSSZ038FS9OIElI8I/q9Kr878UNLv0Y9f0q7v3D3+D2eoyMpEbc47f
cxikiRxZl+OXm5h71a/bbCeOkqciKA+zYiM+aQ+Ab6rjCd8W3f/vpwsT5wfV3GnKx4ORrOxaIPAh
XOg9LGmx11rwve4ogNLqXVvXxv9j/1IXOw7MSis4jfT3Tk0hzaM8vLyiOglXlsJq0cSzF4brzV1b
pOdsUMT/b5vZAMK5rkIHf/imt3TIbSiXwXrUf0gGgkdkg0GUu5Sw4zczuVHSFjI2FoNopQulwKpy
Pu4P4bt+esWfF00z6X2HuSSBVUkl5hXMGcVWZ8DNhSFA5TM9Qxc+qvdEPEjZvkI9KSRe+NvpSF5J
cOoKqUxwDwFhgCxaB90aqsFaZV/V78/79nICZ7TeCtSV4iDIW1Ggrh8zRExJ6lGVwC0fWJwAWhwz
7bA6L6OQONT/GumcNPYiQjDWeiifv7zHn+U2nzVddb1jEZdh/h+J88JkZveo98o1Zw8t8zFBlGOU
sRsNVLOn2pcDKDD/SRB7zcDseVQVrMhLmyq91qyTdvWxFvfwallCvZPZFm8TWiwvhjJ69KtcxupG
N5jJho3nug1AUeYfbUd46tbjRf77RUDfsh17LTT8N6rRbw72c+epYJl4uGn9+waju/QbtIpSbRE0
Q4Sa4HaU/E3wKkeiuLbBYo4DMgpQMoAU9/xbVB7Uronr1smWkT7jrGAmXFgNys6ho4/gZsW/+o1h
blACoUMofpt/ouke0Ax9JtsFGvloPFBChi+R5kdqQBDKQ2BM/hBJ1MlOHLtU+lcknGemguYRwO1W
ZFjKaGrjTnY8U1duqRYooDAkgavpbbyhsfsSxAzBlAI/nvfEud/h3uhPLBeZlnZiLMWqap9KIBJi
dfy4ooOHOAPXhWFCiWH95k0Z0AttgXFOpHS74ML+c2bmiyYSGaLdnRj+ffEtkGNLxy4iaPx0TBZ9
fj31q6La9mH4JnQokiK8GuzBqoNx111fsE66J2de6QNPqJ5dK/hI4xkpcfRJ/phCoMFUG5XrNxqD
QRNbUb3ohSrtlc2FUAWWGKFixdeyXyVTXTpfRcTJ4R4rtrRuqCNejiT0F39jxrf7Gj+nddssCa+A
8FEgdh+2n7yBlDVtAuoztzu4ieXcV39KeAN80J2oqdIuWFKvY6VgbEU78HbvRYRH8xnjFPR4tEO9
do/0M0zYNKOKQ07MVlCgRTBCQJk/RpjjpwAMYPBCE2b6Fw+VOfOFJoWrNwuQSIldNaLv9xWE/WS/
mug4fBrXZgrI8xjErUF9c6ibdjx1DAOpkUCPJS0RGahe9A9p2zWO8cihPu0usNQQJ42jB/+e8lW9
F6Sc5Wp9xLM7mRsKiXjMM2CE+KXyUXbsaiyMOfFUQeJo9bA71C1Ix625kElqEHbhvrtyXhbHBAf7
EhLfK4KdVHqmol+yscSgbj5qnFscTQAHDf8cmor7YJEtJ4xSeSmIf2Z0SEpDEpLY9ZLF8MJ8Cosx
zJm861h1rQMHycUtkCARVH26897IBcudsdDqN/sySI03aG8WU31JgaEp34XQLFB/M8BH1h59FPSD
m1vas88EvT6GzVbOhr0jVCF2zFuHUcO7BW83ZDpSWkm6cvvS0CMF7dT8rA6t6t2f235amjvrlgeK
HK+SlJ1iMtIhJZVjtr2bSJm5Lztv65ZjT54cw7alLA3xLPdI3LqwCxI2hfWvTQyXu8cuxj1llnCt
+x7CBiO3UhasBEwmCL1x4DxmrNq/pZFwnwiL9Q/y2rQ7caL8Us/EdPMbdgm41Qd33Nk89wI6860B
bd8E05MGDGVdpZEh4iLpFw4RK9RyjmihzVhFdM32LE3iNk5jzGAgOKpbPvxa9AXjXxsO0rheaejh
0ajb6yo4mtHpBDQKgmWhkV5YuPKoM9prnqA/4jSnQ8jyfcBUJl9dniL4GaDr38vSvCidpR2TZKI9
hAcJ0pIDGh/Px9OO24Oji2tNazUzKwZ4bs+eN2LfC5kW5F6PyXJ22LGePIdxpXB24xFrgPPL9KBj
2xScTcH7Le5CYljdy/tgJo+6fimIlJaayicZQ1lc4GAzE5Y5uPYdIIexbUPpLAUWXeX7vK4OZ/NU
iBQtrtD5CrIX+W+pPZKmbjtyVaWO4AdPErfbyR99bElB9M77JMJRiMiammVN/iPuWH37/WVT4Ero
2IKq3wF+BDJrjPjUmjT6bTtHu4pGVsdSUJHevU9tkGVuW9sENiT6GYokxAiXQiSQG8rYP2/wIvoY
U/S+8p6Mn2wRDTpdmq5qsyfq76+sNFyIppp3VTU5UTrEGQdCYkDcCVkg3CzZRxx1lbDO2TXe5KiW
Da6HARCgqVOPTWX0lcOaNbgyHXhjmHJBUpCrVjF2LucBg7FIymacDaLxXTSekqeRgE7aJq5M6wO9
wtmmo4G7otj8gbzstLgRzuK3UZPi4JY7qGpgsnIGFwm0kIMtEtQwi3BiUNF22q/riXvSpDsDZgL7
+DpDt315r+2mKy6WPPtuPczaXY9CUuG3sq5T0ht9u8jchkA4Xj1Iccoap3mVjkvePWgj9n/HZcJ1
5hJh4OuXgWi8dvVV1GNo0d/+DNSWfIkw9ZT6UJbYbEHlqWL5sUKfj1WveVve59mAQ8TblCtfkgxD
01BtOGnwpHihR2BMxYFHnqh9JhUujgch2erqgbD7vSkmCbONBJM0UopFXwN0nA3bPGwCWEql+I8X
qAWmomMTZxzK/pCMlNmkNnPiSjPMyzvA7wagJaqwuoQoxwzUP2OkOW1AODbVxotoJPl4UVgmd8bd
CVgJbrF4vj2lal+3qNzQphAiqFzvTUG/H7xkYdsguuejh1WD60z67tZrrLzKMWr6jbLoO75LZ5nH
sDoQDLiWaLMdqo6KySQjo1mx6nbGCI4JpibsBUB9iIbCT4pLczBF+ZalFjtYEYbpGHLxXncPk8Gw
nmTPd8JdqnzFfkl7EanUuDsLgL06o3CV4ibiu9vk6Oa1fdzmdotkCArNp5oBelPotvdrLdoXR6vW
EL90HBs2aghWFE0TK2JsTadvYoIPEPuPtTepOwUfLI02OsgGgsRhRwsSiX3kvrvUxZ8sYG5gCqRc
hLgiOStS7RqCBoZHFmWc8LVfZIR4AR7YW4rXqGgOG6Q5PUQUlKoLvbthz3+aV3iod7ytrB/LxU76
LrnXj6xnikSjSHGEp4IcU+KBRcRPtOwvmq1brw/HYHUcQo/WpoOX49Ys+roCDwapVEDDKOKaitTY
wQlCbJkuhCQfEmYsUqbjmgEW6NNd8rZ52SiroS1yywrx45HScI14hVkJNQ/VyviSPl2wYQblgFcD
XcugVMIS6qtLR0m+naiKKBHNugcx9nb3lCi2FyqQcjLyKe/SyBD5+yNfQv/pHpmwoxWbndiLthL+
DHzfEBOMoXf8EYys0t0sORDgD+BakGedo3EdzWKYf4Jnbb/YLRz+L051s8LzUsaqst/Ax4bOhZTp
j3705AtFX4khTvLUq4H9iUvG7A/0h2xq+Zz5TNvJw6WXbQAeyZeKRmKxSDHJ2XzC05femOGxAxGF
NiA9opEQx42y+9EZwB+vO20gqqU8QTvKMJ5ybItnxucR8IwOSmiZmAAmVLCwAerJFs1eNhDr6Shy
UPIax65hg+txig31ML0HBhC85GdXUMIM3Jkx6ZUHz7lcLEu6mldXeqwgJHMPEjrak1xPNzMW2SRz
ZM1rjFfAJ9MpfSdxHx8JcrzJOyJWWQGC0CV46IEMmi9SHCVyJ0HryxpZMYnpcOhxPPf8vx7OObj+
nyWHKlCIXrUAtPWN7A6C2/3Y+t3WHRBVCyp+NIJZGHCplbdI7zhSITYFSs/eThCOSVLvRpq24AtD
jX4fqfR8MCwW0h+93wOgUrCQ061zCfAZ9QQBoHDHHl68M7bvgrvwukvgCBoGqN7FdEx8SkiXm6Im
UGmIxSFQ0g0DIg2VTcCn9fpBpRwkAlgKLQzVopQVUnSAr9I46gHdJHnl/MFzx2mUdwvs2HLcXvn+
6pSFszLIjdMiwEWV+Jx6F2hhocg+b3uw3JJEZR2kkqQkimWGZ6WUIfzqVNWGl1+5eFmHD/TLcAmq
5j1c83O+lCcXreE5PYxPn8krebF7gsgQRhOky9phKWNZY79X3lFJU99yY5xkK7J3tsxC93busndk
dhJ/9PuVhncdI7QPZfi9ehc1AcsDZTTrxBR6LChqOL8WsMc11O7vQzncA7U7AGPHKOgpU0iiOQJ7
0KjTqhFM93Bg7TjBWIrWSpyzjnG+WnfVyd6/wiVeHhbN1XMw2SySC2xUMTnNmEbXXpvSnpj1ar+I
t58uXWhWhwan5SqegXIf3IWlUgVzs5lKW5ENoP/SHfsqkH5qB0dvJVjRWpHmhde446QMuLWXzmu1
ysVxQIRb3hC6BH4FIiZa79NbqGqKdbutUXF16yN11Aqw1KuNttdh/4eq0cYufKQ8ZWJ5zwAXkXPs
AIEpmvJcmqIHR5zJAmQNAZI0fAC70L4dmLZ818Vh2+X0rYA9LqQnp170MGC7Fm7Khc4fFl+WXi5G
lEl0hhaoo1hR8XKIvGAnvJ4sgYhDyF6Y3NJO143x4PTs7xLhZwrVfy3IeUox18XhQ0KflEQ+DjID
JLv7Scp4d2TMBdNEhDrGWtQNbIAH5ftDabTRFI41krqDvK8+I5kXIkJYAxXDX+beSOtu6aJHdZ99
gcIRcFqkI5Zlc8qnQKXzPNz9JkcV9Qr8TcKDj3Nz8NFRKZwwFABnslyLj67Pt/56F28eNF3ivr5i
ZvTF9OsRwbO+Nuo90x+0JJhp10Sr73v4oCFxIWgZmqq/QK0NIEYdezQvgwLqpwpjH4gr8JjxKbZQ
mLhz9t5bsYAr36wUTUayKs5d4mbeuOczlMy0M+ksN+yBPylxQuUeVV7RtSw9r8PWfItuKtSTa2pi
LXYbckph4bGuAQoN4POzAOFBvwI+tfDAPGlOKygTXIXi55BTBlFOh86t3QFSJ0+412A08nhSKH3N
F5ZGJoe9zrucE0NMfVKpe05B7v3+BhM1PjzsOwGcWF57BNf+6sBp/7h+VxNegEaacptnMRwh4SVw
fQDmIULS+7xFDrDvDDgFGpJHSvZ7IO+JCX209nW3X/qun8JArVHBz7jjI3qXnjUsgfW3o9EpfI5m
70/hbRKp/0jGRVtk6/8CyvR24B1+IK04NV9qnq6iFx7rlwrXryBqxLcCsFl/tr473JbYGSchFzxQ
/exA25uiHt54kzW/3kRLP0/RvU5He4HPKAROXjyWt3jbcqO4bZC7xdfQO11U2rFzrn5kYIApOJPY
TMh/xQ3d/KPdTqLO+DAmuz0Sw6rKBi3K59HyUB2LoYSt9odwqgCD5uZKFp3kWjKnA4FNjZfG30Dd
jl6UsI2GlU+u6Q2dryWJL/GybbmFr5hmFVol2LBzAdsuNFVx8/zJnfFpw92KA+YZtX2JjXBuKfqh
3XK3jT9kdepB5smBuHl8XiPPiKwp5qmSSUiT2Chct0boG/tCd7wwflz6Ap08yyygioUsvbblIydJ
3SltFCGnB3PU2FdTwQbjGIJurlvzgqk084sqJ1ZYxtL2KC2V15Mak73p0Pf1mjAWEJ4ze5kKjG58
uUwdGJMWPvuYN4/423qcbDPovC03Ey/t0GdvyH2qUJIz5Z2j7uLM1Xxs6FXpdq3gpfXka7wz/wsJ
QNNACKe0k9MOiP9s8JgVFsXc0PgtvfGMrGIg6Mh5M9S6J+xznWmZpVym+AwaNLgfXkS7pz713FES
nd8pwKjQSWJb4VjxLK9G3tT7/Cqq210AZVNTpQWAUcJPf7yAxQbMkpnlMwHQd3ZqZNiPKJUkO0/S
NXI9OQQbttPB7s4QLbGDlIi6EREssqgMB2YzI1Sj/NI1rj6SK8TpjN4q05z445KKgp5WQcN7bD+O
7acJVHShfjgkWyuxVREt7TGv6JGhixB51E644qEA160F3qFv/dDvaJT+j/CnwVjknmmoS/4467Gq
oxEADbtCq6WEFS7dbAp08C2AZC/3ZO/LqYnJ31s0Wn+iUX8aOzWOPm68K2wo9KduFsBTz6PwbCqU
tL5MwRW4T7iFd4OzQkSRG8RXURd68ttQhT6wvIWY8EKbEdJbEp6He7raT2TyMjTJSpF3J795npn+
oLINvp5dVI00Z5TUSc9T+NqlxmOLuorwp4OzQN9k1Y/0gPQv/jI8Lm1gr1zc9+IJAX2eDakYQcbI
rhgcZD0OmEhacIRydIPpKLbG+v1L8haIH2lfOi7+nt8Pom80JtqzD9J880loWKrMaMWO8xhW6VmT
tRlC5T1GHlcG4576y/O4RoBULwHCiXtSn9dKc7YvedwmL/ap64bQ5l2IhqUF7ENS4Dng8wzpbyq1
c3jnRNieU5K67z1uepWq+P1/Rqxxec1ZKo9eTeFhmCcQeOJu4szDaQNpeZ99YFBlYEOFq6u6/A45
sRKQPAWqkRDCC09pArA/3uZfIa92MUIsx10RwE5Ovuk7qwP7upLz94E4r9hyXipUaew3q3s69ELk
bdrCNqpAhBdesWzu6WS4N0zrRDEOUp0CEbc3UNTDfRV6vAV1W4FR0lXyoIHaZmD6XZXTKZR5aJWv
QMt8lIWEUTeGmSqWxrtyMREptnkS7dAvu9irmr0N+kB2mQJIwbUbFQgMRtWFsgDIyu04Bxb325fk
XgrW9VxERc1ovECEvPLbzFEjedPc0Lo7mRcevEyi/UwgVsnrnoRAD/B9ZdBo/J5UZNsyFBtFd4w7
DtkydF+sOPxFwgzhw1hNfKbJgMH4Bgyd8JX49wVtmXATXPxeD/jxXfIz0P8nDHBaoC5vW5xORbjD
auurR3waheGtfhpa6N65MESbJ1Ia0Ze620eZov1jROQjEttEYv0cPmJMDExW4TfhfOIx6A88zywG
ccChkBD9DlJHFB+yqh9c1N54CSo8myVAswZNnLDRf2k0Dmds7Yvd2PdR00E13glnwfLxgmcVewqb
ezvvdGbmsfEIbcb/17rxW3tJ0eO00YnH4PWkTTb1HV/VuAqYiPfaMfLJOTjq030M0cuPSqr+BEj9
5zY3f6+wNk66tvzZyrA7AhQ+KBDmfN5Jzxvkt8L3lkdh5lfD3Fm98DRcANLypOppZDZREwaO9PlX
QsC7JjJCX0TmFWFC/8yDp0tt+Gd6/8BFoLPiy00bTu+iJl9LGfetpcbPrn9qbt+f8zwuk6gio02T
hyzZu8LWgWVoTGMzG9roCqfBze96096c9ggxqKP+jVpevueo5MOkyZvXHq9I5ugwxznQMz3otjJq
GBc1xWHf9nP5sU34i4KmqMe+V3eEW7+017ZEXkc5AVVc6hjlXTCrmC4NxQv1OCa38Or9+ZKaZFUX
wLupSYs9AIRguEBo9yE8FTznpTLcbsKpesb8BqAaU/wfs50IM0moZtntzI4JnF4nVSvUTJhlOMmo
i3W+8RvK1Y0o0yfoqNw8kYvPoOSbLyufLWczbR6n8H11u+6v35x5PfLhFV3/DK+5N8B7RcJ5to7k
yNxzNaowKvALxl44G0P+kj+AgckRiObIUXC37toIZKTP6UYPws6uGECpoT/xwZdim4iQUF4Lpxu4
G8rrsmDLYXeFM8y8XDtRXSMUwCWvYlC7UbB0jyk7xDI2kFfis9JIysykcau+Ms5BgbRf/J1KWKrX
Z+SLjfzCCIrshTjgsmlbx85p2TCImtqBvFdzpRWhop2LAOzO6kT4ArcddzASAc6d4ISbJ/0kP9ZN
T1V0mOaT/SvoirJxNJETZJj0gEKVOymDDNQgG3G+ob7QbqJDwfxGOW8g+9yavPnEjG65JYl+KzhH
Plfq1gKIIOH8Jr1W+Kkm6jDzLcVxzVQFcJpCK/z6zqBRmmloNycduVoq3mP86EqGfcp2chA6SJpc
OfWQ0NfcvPw0Pqd5/MAlsW0mQFmii2M0K/9eeJxaTBonfOJKD03EdXFrJ7VeDt5TcdyKfOaYKySj
M5ferLgfM4aMUQewFDIBKtH9xYrFIrcBegi5aG4IDoUWBjpX28Z8e5sooFBYBIShJsK2f3J8stjQ
DWyiU+XTMwb+I8Rv0Upk6T+f8J9TpBfxPS+rV+ocPfE4FqEfMhf1adpk8A9jUQvhPDZ/0UM3FDpv
ExCmRC+qN+IW5b8ccbaztdd+dBoXRLx6v7zl1jW4UOe4OGnKFE2wcoGOJuoMIuZkaV7IjLfR3h3b
T2bCy+GEis7soy7ngQXTHns6GXR4+bZpqOrYi3OhRC3eC3mD3hEMBZwGB09gpJQY8hu/XdCLG1W+
0soMqTlDqvi0ru4Ka9jABloDUI7n2vkiN3uHBcBvx2vqYeyARhUUmAkwosvp4/cGCrjOQUrX4SBA
kczlMioCkYOMCZnR/yEwtmxwNiys7ybB/YUY0DnKCXs30FLmzd0NxLeOdWYqmenT4+NFCzh4sR2R
6w66vItU+KtGcuirtmouJztAMYXBaV6l/6shBFG8gaGZYXNaN3A63uCMzpWOwHKGHrutD4KVsM0Y
hyu0PPhv0TIrm8pf9NW/v7xlSO2iwSgm7j6tEC7vlsUzGXWvEsS43ENG2EW+bU4Dxi0CgCNCFJ9G
lJRBFMwscjyOuOlSuh5EzlF4AxJI+EYOZqI7ChEq8r4l6gLckGpoS+SovaJUXcoqkWzwfVa18ThL
XRpSJJLaoC3sEpN4BG/Rl78klCpSlVtZiz2kfzoWt2jbcEFT+Q/snN55Zp1CGAizKqGwxbQUWfLP
qfYVf/Sgr+Q4rQTYwGIqwItXfMHQb/Sp4CBUl2yJwGwK6R1qCRkW0YyRNjlljAii3/D+zQmTPFmH
+B3DlAEr/zoyFPacJd/5EpO1o6HPRuQd1UCnyayz32l4D7/o12acEDRxnG2sFmb3k5FyhbGw3RFU
QUWb+WyDxNq1mWaTfH+ORxQEqGfPiMc1WeZ06AVPGUMzXqGWqC1z8GF+es72Dk9ao0jyCjVYioBZ
3ZMXMiPgP3snQW5DYugawDlDHQMeXv0CeLddkek5TV7lLhsOKemvzJFOL1SbCicfKIPWb06ypkpn
T33mVPIUN50ufAl3gxBre/denDSzX1YEm8ir2SOox7diB1qRJQPJD1WYXVpCgsiwEOP62yDXR45o
lECEfzKvljeYeARcZCxVz5XtJviDTJ6D/jz6nu7VebQ2vLmwH92Ylym0yzBENcR9yNGchfhBN4fH
3e5W8FxuS5bLkrSS2FFYxPpQ/IiSasT9OonX5D1XciOE/9c9B74pDzXgStpb0EejMYtiVd6ve8Jx
G1rEUcrg3/ehpd18LDSl4SO03bbL0VIlQ48Lym0dO+tNtLZUvnRs7RWYJTsc+FOTe5B46heTMQZ6
F0bw/snSCSjwvdp86DS57B7/HL2sgjLg9MUxOppxgUURKYesxoFk7eXrE+skPQLiSHGSXGKdwfnw
e60xr3VavLFIhfbsZTzpQp7YSEKjD7UpeMyPkGeC+3A5snRVu1as+IPNcmlcw58U/jl0jMIBkNm9
nc7jCgVduuX8HOXoNEI7Y2uLZ1qyz0T5ainku6EuwCYUz6OPxYsBrimwSltS2MPGUxxSETKpGHkk
ZET06rKUN8qcm5kHxNrDjJazae8DUzhhNZGaLK0k8GgJ+8kIDDn80JJzYBMOzG0FZZGKJPGvTCuI
DSs5c7dq49RJXHUAgKvxKJDhEYjGS+Cc5F+2y1hUmYsIHhGzRCugxmRdl3GNDiHaLzTyQyKPEP1C
zF5+ziAhKSnKrLSS/gAhv2R3s+DuC5dELjkiSyHxPjUm54RsDU02QRRG10UtS7gkF8XTx890nave
IQiCwKAP7M2kF7MTmaN+D8Jr2Zq0SuWVisA38CbF+z18282IzmHd8MW/GfTU7dSBJXC+4JjFCpsr
asYS+NZZyyQygqsEsRtuVozBKrSVnXAaEsUXyYKcdxVNTjtxpsfQ9qZQs4cmt07n1JlDe+UjdCql
ADHOcQSQw51fBwPJLlFTlg9gVbcp6bfKfU7zCI6irmGH1X4oPT6+hgncKGeY3xaK1Ot6EQFQvs0z
wWD7m3wpCjBPHIOo16qivoiWBcKCkysiaBHxxe1NoRyy/xUddXatY2XEi6IzRgn+ZqZV/MfYyHbt
mvhBJnA0EPnsLriaKr94SolKKeV2sKV4iEBH4zsIPVjRv4urwdNxBvTJczOVufejL2qQCne8aGA2
8lDqd659SXv7TmC1aOx1ri58IAQ+5ysRVmzfHctETbMxK6SWqE4IOxOIpn8cJd9bF+5CA458LwlE
D8SW+25uPW9+Rbumie7U33PS1iqDdNjkqHjDRPsQ2oGOlHvBYsFANdb3pBSicGgoq8W+jpAaW/RM
Xo1Vhc3wCb7fD5bb0XPNngmGKtbk8pY8BZtQZponT4hFCzEnZ3X3BVXusLuQokqYxBgyrdCG9lHP
a9pi6rirrnuC+FIGPDXZVyZZBqCMZy/XF2XWzPD151y4AzWvVR0LJS4ZDD9D9Fvw5RWJHRXy2pch
opA++9pYojbX3STiRAAt+p1AkenSC7OEsAL1kscrlnEvJ6VkPh7x6/Cd/T71n6i96D0tRV3FUQ7k
aOr9ZO9N3EOV65DdungKfVH8eSX4gylQyaHXhaDespCOkh8ZrRA9a/Jmo0cyg/Hk4WGxAo65lshW
haY1tPT2fQrc6OAYrOisrqoYLtUDi1opkZ6RAoyjyuTDeZaNpI9FDiBAhWQ2SEzgRcEK+QsfPoUz
uwHnMi3W/8ktl84zIy8sWAn+d0zxuYfBW6rzYY/CJoFpRpGWRInNIl6evjzxO1wm+fQORGWJ4Cyd
2aYPE1iyhwDgJ/K8Jo2R9eQgn1utyJET8nGqHdbeFzXt+VhUYOdOOtTCmYXWYMZAGI61trsvRc8/
gbvDuQqFldNevsnNVkbyURl0SDl9MH5UvzgT537Z2gkd9NIE5FPq6if5VPCZ5jan5hJZIo9RoTXH
bDVywiiFYbcVfojJ08ifCJW2A8gH9HIKn2LeGos64zrYBm/uwZTNsNYI40E6TFIX8YtD4SgKYAs/
X5/1Z6EuLFGncz3qOXdUpuHm8gPICJdlswWELz3pC1wrrjtcoegUoQRscWKrGCzDVVxoWVqeYIW9
rSYM2sfx3s2pd+UvLMxlsP+0AAdWIKKmuta+OzNy52J460nYY+TQetWOZw/zLx+V1m9VleJSXdZp
Uk3Te57MiT3lmxjK5d8ZlvjHz2lc7k/Vld4h+k6loIc/E4JcdpeS5QyJeSD3Dwlx8p0PuCQiFzBy
+7uisupa4LgFL60X2GNAoYbqamVpbm+cl/sjytvSAdTumdtBRwFVCmCfSpwfBtghDqIfppRbmpJf
7N4pNYSv1HiOJ7kCWpIuSq6RznwDV5zhJUukMnf2Aziap3s8HpTASfLWfpj3tUWzorKQ2e5BHJ+k
H117X6pQy/N1Gqyybfh0FucDxq0/Yl9u0dYV/PKS6Jlat3/n4Eb+6vHjNKg3SPnlzItJd7dDeinI
q0LEpM1QHQeMk2zUWA/SOHWHlgyQrjweZhuRpQKmhLtTWknuOIRyvo61uxhHG5vnnkKkZvdzjuPI
dKraabCrVI5xLG+AGtJueDpyvGIIjnM/4IIKwK3tZEWQhO79fWk3tb4mkzbttLJWQp3D6L6U6+WT
2+DtKEbtZUPfr2j/BhE9eyfJIPogsS98Wn1Ix0D+0ARnmB/orkmXml9tcTbuWIQkESOpGdDBy0Rl
1Evk7sRYUYIoi7dlnyoJvAoLSr8V43tkaYPYWjszbitWD27RLQyWI90g+ycdtLApxvTaADD/HxgL
GQSjTxk3PFi6Z0y21u3GlowZSsuTNXfBCO+ypOO8pRShutdEzpNaQ347alw7gep0e7eZe5KwIswh
zPxPr0mHD7WRd+AVa1Yolb000ojI5chtUo1PXa/PAEdEdVDsJLsz/2Oz+qyuzk+dR2G8PXIelLuf
ffQbwelHs4vxkYZwRl/mQ8WE1FvOCoPnyUkrRvtrpUWtLhTi33stjooiSvHz+7FZLMfYV9YgTQvh
E8Tim1UXEy9tV2ptEHy3N1OIPinDjceom+e69DM5NhavbGZgDQHKLehaDXWI5JUETBQxVLVoo0WK
5PxvFRKxFOExqDueBgZuSkBm0/gL4sLJ91bw9yK5rvlv9wfCy06IoiZ+L4icERBOrwbZDlmUjURn
LQzXjjXHm/d7GCYqexuC4r2UaL/Jno7T4FZci8+Ferjclk1RolgC81kTXmBU7RQa//MSU/WFmSOL
INz3XBHKoKGqj7RYQyFSWnhFNt7QHePdvsGF42xwwldbwymEqpDnDnFSKQInihH1dCSWibMOqApZ
cSdGQzSwBNCvNHtDB+FQCkSEOGVjJ3P/CM7uLkd/45nofZWEAInKJ/BSjf1EBak93LisfLpp27PX
Sj0m48EHPeHNhglpREv6Glo0fEVuSzZu32Wf47nKqxpaLGifz54TmeSElot8cm06a7a512g6m+ZH
ouh0aIIeV5SzvA+9/lPJDJeTtzh1FoZ7QL/xUle/wNqA0dZG/sDH3CQ3449ncwuo0T/pyj6ibQ6m
6P8tbnzjb73fYxjFGT9xM3qg7jChwMNEe1sCOvMNQMYDE/c2UJQ0KtiiYur2OrSfA5ZAE6sNddL8
G+gZcFr3qI6DMw6EFAWQWYKbN++iEefxB9BQDQPMLDNlS7IakxUnVXdPndrrDXtBYVDCRqlxcDr9
thmZo5nLH4336aUFfuHARql92U/zPgRVPmIL4YhOg4xsO3u+GdAGRb2kyugcDEPFO7/C55CLdMly
DlEI0VxlbFPsoY56dOvxMTVoRuxxMQZWwO4v+XcXVV6jgU4NzK1NylWkfU/9sNo4NKARFtwLakEB
bt7ejXDkrGUQI25uaCzYRz5PuRcTHubY8Tn8qEYPBfQnElZs9Z0f9GLh11lLg678X6bJwJi33kjx
7aGxg8CCzuv5IG7CaDFcDYClHNShWBGsg7/33InPhvgPeq1D8zdDuGGJl+T3zwFjVTWzzxmxpNan
pEXGopsUe9ffWtkhxQPqviscBGqPxp2PYPNFQxlztXkr0dTeuwAmrN4zFKG80ISSAsrOyBDDuGRw
szI3SqHY9VphD2cIf4Pb9bcZuHDyJs/azevMvNLIEgfN4HzT1nJk0pDfcTMIIgNOYaR15c7J5aIG
0MBMwg2rbdnBnYJXoUVKelFq0Pkd8U4pD7xOEfZ9zDAjWXKwFAAAfg0uvWbDryMFvzMXRpG3RDiY
IF3/mh2meJ7wONq/jU4fqhC0RlBXbOtNByNlzjHkhCqZojJ1BQc6bAk1s9CvQ42JVTl6bXe8vtKg
HaiiY2XA9rQ4A/qcurf2MHFoGk342u13iYbBt37SQcv78LOmrD/MucJRu5hhGDaJNOFwBCWGgNdL
xj77Zxuk6ffFFlqFi5jKIYpVi7EssTOPIFlL4IrXTZT0KpNn8evp1MW/n2qCZcSYCWSsxUn60s8+
+6GX+5bWArE8fMGFYmQTlrDYySE+r+LrJgibvKOMZPIqEvWXA9Lg/Vbp5zjhxk/udUPgtR/QK8mj
GF9lV23e7xhTyPSL1k4OjYYpZEXBKCkv2JW+Z8KMdiV59+YuVSm2gZsy4P/dwx59Ehlu2SUNca9X
LfsgB6Ay8LjwalVpDe6j7YHsgNhRCjXR7iLFVQEO4TAMaizQz4JNtIzeyowu4eALUkjbjZo+bbsk
67PhYfmJvZLgdfiHoEsWph4oh2LGmV29c874qYPcyZ9VA1eEVVT41KEAvg3yb/c5iq/OEo2nQ8EG
OJGBYdssJGpjmO4EdIlABJq86h4jVTDNjwk9yxh5IhpexrDCexBIHykntHXaHrY9OBJVJPPoPwMi
cz2myHh2WRK20q3F2NW68gud0WiQAt7mdjnKGIrH4mN/eX8KenomSvPpGnp8trcSjU3nGo4/+60N
kI7VPhMLRRk2q1iWS9jenYN3niZ2Z3sjhX9zifpyUHv+xsh8LJJkTeoIjhTWzEIqX80UsjTwjWIM
bMeopkLSSHm6hsoZpoHSn8iauKe6Ez8R/vG/vZWj6r1GzZpQZmvHcSA+7wXwVgb6hQFBWlkjaTnA
Wb1ohH9uwwNoiuXwgtzCMRk9iDipJdAXTMjkXlmuGz3masMOQdgNGYd7u/634by7uXM2rq0QkTjT
u4QHHS4ytKtCIPVyLhkr53RoLLKJBhw0t/MOQt2WnEhD+FFq6ukzvtsLjgC7h16d2UZDPgxkHSPo
9JoIjgvpXFA20IiidkIcZGzvJktF6jXfbreUQAb+LXVqUQlSdz2HsatsE81rCcklvr5OA0mXgrEV
atRd+fC7y4kby4c24Q1mimjxY2idT3f80jvWq1XzMDeuVzqtREG+t61lxsJN54WjEjmweQUCzToT
Mv7aeeA+k3pRUuQ/YqMuF+23o2NvEzg7uCTilWxc48JYM1YLw8NLAUnfzyc/EgnvTOM73t5gECUO
g2mppkTBnk5eaPzzMZxzChSPT4TsUdlkk+Q8E9sKr3iPdBQEHMrmBDxXqcrIjonZKphp6ndmjFxe
6T4joJgday5LCs6UC9bseEL+xG8eif3w6oNrFoSCrvpKYij8Uxoj831m8jqLC9sFx5b2TQV1bMn8
MUd114CfovFFjIb9i65EAdhLplPxVzVLTYg+4mX3XHOgungU33kangZWNz1VAkbM1jKFcqDyuSv4
CE9f/iTQl1ln2tEkz1+ULWsbPuBqHm8D5NHhUua6YgmNbYyW8MT2x3ZVYGgGf4WGjbNA9rUT2q6/
yZIXC8DxY23BktkkKJAhsQ1kPEcpGzz6sG71TzDqLkyNtpaZi4QRV2v68EH4nb0EnaL+ixk6nct9
C1j01WjySzP5NfcakQrOV8Zp0KQsXFwk4MVZi1l47Ergjl60m2Bvi+z+CXbT/CWE70v6+Zlfa7+4
UHE/na3E9ScM0ttnsBabQ4EAEUv47r+aI8+j3LALDWcfxWV+eR8NE7MtxRFirrRffls1asVc6eHd
Ll+SdNeAqeTnpiqZTlLYo+lmpmhxu3poRcXfJawI0aJJWLa0GwehjucPUp578TBa4ORF4txvEvgy
7PFE3Nmo18yYmPeqqraIHugLY9yh1LUcVxcG200DR0FBK0O/PD4VIHv5cM5eGXhdG6e/kdQCpedQ
5cpNw4vuKQ614pLVFoQw4RHLXhlLaLe4Py/rLqj+P6JWWo1GvQtzYI1BbSgDk9NDrW+pkSSk0pGw
boNkT3GHgnbxQxn8vc1g9MbWb1e3jIdO4WIC66+nAjMNlSfW6N+PTnShE17ZzEs0rjf5+iPtWfDZ
mixUMlWSaG3LTD43dy1SkIYIm/iwyv3b4ArroovEdrtAmuZ8MUyhRioV1vsTaajC95o6Fy6ZkU11
JxJpdHsCc9N6XWZQP3xatod8t9ngapdVY30lUWgzOtJWeF9tdt9DgsJJXqb3beOLr5r+MGcT7aEr
Agj2CooDnkr+D6eucwUyy1NDjtRnjAcwdEFYorsrkEHeqKqMZIAs5l3T7qX6+edKgkjx7lK43rPW
0GIHEKfwSPX8OB9OWA91PAzXwnAqAMM2rAaUQdv+oe4E6GP1rlD0DyDXC99jJJwqRbQknFlWUEXD
XrUo8V7mqUhPPoCrn3hH+4cyITpBq77GtAw1ym7367Ktu5q+nFHLdfGMDoVcPzE2R+HZIn+CbZ9z
FsGvPHcLIoM+CJhHT2KXtL4WdBHfZhabKMyns4riYeN8rYTBQdCCiZM7w9UOv105i6dEquPcr47Z
3CKsZ/0tWeJM71mhttwhPDoa80GMX/V/QB2sqRmnduCLw3xiPOsbU4iHAzWs8nDCRA49bI7Mc2sw
GIT4eIQ5bHYveifNUfMd6LditeXoM2Scow5jGQS1qlEUvBqDN3XniP13f/fv60dWQnQwAlS74ZGA
9+WCW9MPNZ+t8S8xSuRKkyhZfYAOe5wUTU5xTgC4KRR0ACnKzY3O/bBVdTvMk/tezj/afQjgcBeC
D3fNtw02RnkXWFnnWZKvU1iJk/nkTtqpmaup4A0xBwOrjk8DAmDKGfnkNVuNzrHDJwrCC9NqgPBa
NbgO5ToTP8Jowgo40Ycg/nF5+i1Ym8R52NVsN24tIdF+SlPZbevy79/AVD9L7+eSR/wsLHxxetG7
OAEJmaupTInal3aMNdEamMuk0fbfFdv3Mq3JSVwOgJPKdPZloG2JepubvjlLc1GjswFrDQ49JCDI
M+KmpdgY4h+lInDOc2+LuUchVCK1nGodhg82SrGXzSlPOFzoUTbe9SXt/dGGz3oXlnuFb2i+Fetn
BE0RCsPmkDF9WNq3UAs8N07OCDICxAMg6w3h+2KRjrtC3PzKnHdtCXoyj0TsZW+jKEgZFo7Dvxde
FmmQLxsjEp4Hdy32287xf4yxeSGK1AO7qxVQiyZDPmzvocrwHtZP5gLS3u2ZeY7ZCVfJQ/I1Tuxi
B9YHaUInmx+qlWvrYUW3H8KVJtWzS9oNKzDyT64lnBikDp1gtQZ78gIk+CP79AWTA5ljQPB/xFAK
MLukA34TSeIliDMr/appm1yPtr7F3Ys9EBr3lAICvCkCAW+G1GWJ4+r2hM2qKOYhQcAwbTlXquWm
C25GFRlGJY1B5m7VC3RiLUBKfeY1RFcGKvpQ0SWYhSqMgZroUi049w9Pp+tU4n2Fz512NGKoXgkd
b7mtaDMvDOtRsULmtkB4kJiOfVcg4dnFSHfOdMj1yCbCQAewOraJjmFsDO016Bqb63KLBsAOUpF+
bLAMwbphnzqX7N+zzDf+1W1Px150cq97VJIx4bkxtj4igPnbbuWxyc8XHJYD0n22CdXGqXdS4bEb
xIzxyugApotfBxlG9cIQsA/C8RIy/DJkkXtN9MaHXP+r8rucN5LSMedAK2YZsSbKOqFmOxDCyUqO
bAksEK6cNJRN9dCm8Tkfxxm1MAuyJuwBiSH/5enmF8yrw5yE3BuFZbRHOgL6nI+ZqZykUvJyVQLT
6qjLEl8lui4llPX7ND/gq0m2lDPAY1mbILq17ksQQ/KM243bEAUVV8hiN60171oRouptMBYkoQ8p
P4S8UKd+sPO9KJA7fV40JJ1cINaRruYYKFBY1AMUiqejOYeJe1WMjyZn45D6Ni4EqF2oHmme1s9p
1qQ6hwoHdPsAUML7P3TNZ6bR7PyNL81I0WI3eDW7qmClHiWyLjmAjG/t2zV7O2jvMgr2DRJz8VC+
HbrtUbSJMYcNbqfrTRlRPNgER4E630fRpG38+D12J0hz5iiNjJfWmYU5d6Zvohux0DnzcpDSl0qT
1M71Fyg2SnZQHlA8eoD4vHRrVmpL2Q7di8U+skeLoXEid3o4jfr1PxVeJqabl9eNvuJgGLW6j6dC
LLmC6iJV33ILQp3DDROR5sIb/YmAmCwPnZqsY3RvsrW7qMd4hmrrc4TBYtZUHk3Y+OYD5nNAX9wF
+8k2ThtUoAsUGGlAmhp6b+ar7VMEqeMi6Hk+svhgrYFWlw6D7J4dlH2LNJ5UlH7OvOJNF694Bwqv
BywZHEIcyWJYnXTZUFSwf5cSYSQuX+4FPYkj15ENyfXqSJkZ24CnHlk3UXr3G4TpJfXXwVIO+O28
MZQuqOs4U3WU+KXbREUCLVEWSUJ/EZ/X7N5qEj2h5H21WTCs06NgCf2KJMlTwKPyiWLzme72yGpm
qzX3FPmYtK/sEbebq8jcy3lSCMrMwyRB0WwMYtJLyR7FQZWrGhkV9wIpdbx3Syr38/Kyh/u5G1//
YdQ5SqhByppydLlnR5oyhsR0+KRlP8lg5Br1BStd+OyiX1bppJQiD10UK3xEftmgcDsExOgnjr0d
Rkgx/H4FTqf3i1TSoeZoUIYyUY0qnWzFVivEFOm+/6VR/HLQwRgzznyqt3fleRCVTSIVtmCYFAWP
lnYTo584J93WJ9RFjbPcCeIBTN6wzSQKtbtHV+MmxJxzqBwECUbGo4wFR6u6ckNCXuMF8xoeR+7T
hj3JnTj+tVlMHF8WuVgmtlJPHacggQkySQD34Dyo7RzI6+HDY+D2oXU+iw2FrvKJkPewZcxYAHHv
Qz1bnvKuuWQEqWAnddxeYWIxib3UlqjXChQ25YeL4yjAsjCcktdYlzM8NK2zM+RxdAzpg98LYhUq
CiL5GEOkKmzjT0qmfrrMYxi7EWIrKnTlGsBawybUH2nBR+szwTbqGKjU3OAyq1K3JOskylChJMu9
dkRQ5evUrJ9da0mQ/MwCKs8KfnqQg/oe9KpIGNOOgIpeCqleCDvNUkgHnOzNBAeRyvmyBGSfaMPV
ix5A/ZL/oKYdBDMko2MzoORu2dhre4oltBZEaUvMJlfPxOKvYhcxre3nvIHG4qPtIcyB5AriFW0q
f4ow8HfIeRJKXRSN6d1TrYi/bWxkW5qAUE46MYwTSHRvhkNWrQ51z1vDRH1yZ4uojBhqwwjKRBeK
R72yLLz/EgudLqEzTnKoAFfSbR5USB2cRQiySgTZUUi3pgDi+kc5AlO4WcaP+XxG2K89B7KPGjYT
ywoGNkf1+riiLce8HlWtwjQWHuR3ck0OLgCsYe987JeQZb5eeG5K+kRSXHOGb71jkMzrJDabBKLo
HlVBa4MW1iJ1hEcKuCrQxkkFDOYvCVcNITsUVQAjyJmrVzPJ7yjkTWMeMXNCb4cAzaKaPqpBH2b8
oYXsxMwDnzGCvjURD0CTE6vv8D6nOmWB/8v222+2Wn6QApoideJHgbVJ7Zh10RRrkYnZo70RONOd
4LYN64UzoKIxH+Foy0PDIiog07r70Y4aJTLIBjTQghVA85g/coCjjR7mULlAHZekQs7QOv9xuygF
cfKhDhf0wVleO10iRGNQ2nC7TxZbdXaAY5yBMO2uuXIFxRezg1MOK7wcgaZ5maAL58oQYx0y/POM
EU8CjmmT2YWLtYhKJy5SyHtjrP3uBs65qBVyG+9kP0s5KGCqrgmvmnY45a1wM/pQKV3p+ItodeFG
1v1dn/WMswU1m416Vg0cniwUKsSbOLHOq04xbv56ArMGNOuhU+ZU4A4tiU5vCqoc5M94HzchyJU/
RF8qzHmj2p0ILFNZIBCtr/CVusgmovJwyGpU/NtbceYoxYu/0LpNX1BedYzLhrkz/rCW0sZVcWTd
TfR+qCdH/tXDYgmTAYxZxuSXDYM625Vg1nSU18rCNNiieXv+Hlr1toReGi88aX8sOS5nzqrmPH+e
qMVGxPSmmYD6MqcKJz8vYz4FQEjAzxbuAw1sL8sQyrsGj72PLMFIEhvu6Q/RTNgNeFIvTq0m+lKl
TO/hEDjLHREPeFDOAu/UpCUWe+vKj08w1kwsyBncjSes9PKQVemeyp+adZDxj+UbHWqZlXl3Kmec
GyuaTMe2AOIUp8QoDyFo9CD5gBVIWhv5xiJRf+nAu070P0Dqr65CnKwfy9PUpjjc6deycugctihW
sCphWNNaCzYtayK6DFjz6Lsi42qDEcViqMd8J/6d7lLFlTEUzJW1BowdhkDxLtsG1ASwsdBGPbcv
cqv24C9E5gB88hEBEioNo+91k55178vv8AbR5Dmdln3bTwMcXGUHjOIZNK2C5lCI8cBxDknKQRx3
6S20hr/KS/tlSZRT/U3xcmvNCDqkliBfUK9mZYkdQMM6P9jW7oIFfLHQquOYujYuHJPg6rhoS3dd
eXRsU2AvP+N6O2AuJK28Uan2KKLyFsnZt/M6blyWiFkJZPcdFuXsOFxCxy2lap+av1xlohQmvhau
KUGpD1M2DLe9fOlz4RNgJtohF8viZP2fjKXLYKuTFvzBMleL8vQVXI2LXG7pmntd24rywJaKjYS8
Ow9nYVZFK+hAwewq/C/2D31fOv21DAAzXogpmdIO7i3h4+GeRv3PZlqux/BAe/R3VbZJVouiyY0c
Vm5RwvQnsHuPzTGRfLLKlVncQengFh9SgSkYu9UW99K9iCBDw0LMUlyEgULVCLwEQRn7U9sdhib2
Es2Mt54A2ICIIqwMhuwjDOmAKHVmwl707+WPat2Shl1KcqxADuTYil2KdLYGj+UAKrUy1/+W2IWo
uZbvMotu6feNDj3FKKDCQKLeKyQsGb65z50zFixr4VPqP6UiTzsSk9TVRuwY73NMu6v+wKF0ravZ
ZYNg+C4KtXfCed/VZEmMqi2HdMMPo6cTDyrBSxxQsU+lQrJIRMfbrYFMx0tAlyPmyVQgLNPFacS5
VaH6AhcE+fonlTJHoKdSgwkiH+vJB9MlXF7YVsr8219Li95ad8LHLJihul22hvk/ufM9JHq77Vkq
4nCWS3tKTky22tgA/cmx1bszhZ6Cq9ebs0OZRRBFPQXaymv7Er7UyZ/6Ruf395MwLIZgUG0l1uyv
8BFr7xkpxLHkm3AZy7G5sNyAakO3Av//QNRVYcmg0gwLCzUNn+SyPYWq0cOGWXJwaS8m8NbgchKK
lFixFRJ5Mi0gwseM7CH7E/2/BUGjBusaFTlmzjYFDdgnbUUd0pb0aWASL7bfXmbQFF35gKxOLKK1
vRHD6GcjhuSVsUIlxQ6XuxenwqrozbXuCCrx+DEwBERQP4A80UFtzXxesqmVcKXQAwLbOn87prLd
sGO8Joa+867DslLKaTsgOitaP8i1X2dvajf3D061X3am2p7wbE//89jz8ds75ovjp7Y5twMa+5m5
PN8HQhiuWNVRNDv6fTkG27c+P0px1AMyTOkiIUgPil9A7sIV3zisDqlLNeJPV4oycPxC0G6Kt8mZ
COeDu1KeFAx2qNq9AzE1hAkcvyQ5pStm+gs1Zy++35OamkUk47fHLMB+Og/5zadO4UjBiOg5iPDb
4YbV8+qUQh9+sUr9S2VDqSg6hhMGpI07LwOGLOJp+T6V2/w4ZiUcC6oKNzyRwBqMv1udkK1PRZ9e
5ytr796zSnALsKpuaj9nwUo7fL5mT352B4f6MJ3i03zXNyZNtyYhkRgzZYZVTvgtXhKNe0EzJQXj
JlyLqdIPoxohIIQ/TP89Snpm/o3pzeZBx1PhOwnn52ZNHnLK7nSME06mPhSpwEAmXcijIcybGJ/g
qEiCUGJbxgrAhG5eLkIJMk4ktI1SLVE4Q1YtNqIQpu1dRk/kjLnO44KONBUR1wZAgQ==
`protect end_protected

