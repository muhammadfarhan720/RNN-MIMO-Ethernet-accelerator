

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IijDYFYeRdzkel5iYnZFe2NzgYX9UDO+g6PdWiHeOm5P1+m9Kt//ktx0y9l3PqUsSWKKIi5tWbDg
OqtBZeM3zQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TXFD8G5gE6CUfZ/9/aBQvAaQuQ9Q6vcW5KJtFkYqsiROk19a5PsS1gCxUXtSJ+Xt20njQCTMz6jx
UaSmsNRyiV6PuCAgdQYvfeJWiNmQq7kXQnkYSjycSJyNe/xoXEYIK0mHX7J2x9ouXxNx6jQFR5Lm
jxY8fR7N9m3PTkCqNTI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
0bdD7I2gr0nFDramUUXzPCEqtk/eE+vK1bghpNlKE+S5t5/NbqJI7gNd3XLwYh6qEIInU1StLpm1
ZEERnCmEf4+rQBAW7x7u7nIsJjSOmPWtDc9DLn5S3e1Tg+IzLUqT0rFFh5TiwuYq9A6oIvI4ufWQ
WwoeY/gITSdj6C0JQ3GFyIRhxG7psQKO9U4fj8El/Lb3YXG1+IGuXZsygyLPjjOU5LRXKo6kKsub
X1PFDvdm4rWaB9AqoPLCqp654KCyKSCoufeM/jiWRTNXwf6kL56WQKDXuyAhrasBOno4KOT3c5VP
WEHGNdGBSdU4oUFYiOmAKlCKGeUNCxMxx765QA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ppkak8ss4yKmNiAZjxFq8nn58TDV/6CNcvQivN+uaaTC1viFh2EDUvJp8zqZ2dJOE2mTN9WJY0VD
93fjF/bEPMptIxFj5D6ldjwJu+xdHqS9FJ9Wajnbu++DCTUtAQE+y05rqhCz8aZWKGNejsRfG8bE
xGYNUIbFoZ9PYrDIdRcDSdZRUBadrAC+WcEM6+/HxxJq4Ly/w0BVbiEq22B0+4wVDXszrocC0mKJ
RPXzPj9v5D5aBX2ijUGbICpT6JkVGAjlIEP7HZoc+Ooxppwgc01k8snVnPVI4IVVYOjjlTQgT/qU
t0doYgFMU9nD5a1hefzXRkszYn9RHVZE5bl6NA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KtmDUKyPqH21pzMoqq9CPc/SXFhh6Oz2JrLSFRZBS3mGc7ebGc8cQjlvJpJA0WNJlGqACicdvN1t
A7mG3V1xKtoRdR+2MhucMQ7loisN8yDj3+zqgbM5bAdlz+62WovuGfaM4EK24l8CXSfBLVGQ35JP
2zB0abBrel1cOw3DxvSIS/5wueR9/Ul+GoLmD6yF7cV2ne7eGwNXQ2OsCqdcb9wK8gNO1YfC3kE6
WwdUtjutDvyXnV49wmg6nCC8RAPNWbIhHiMMtpDjux6E1Rkd3xdCMDrxrupZyNQNtVmzcN8ITAn5
BYoTBON1CKVljCmLov84lxcdcXGcSaBAtLIiAg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sjMrK19OPSOpuNhtGVc8GPvvQoA4nRSUShUtMXVan8pbxWL4SmeH0c+Lr407Kf0YXDBqUDDkheov
bvkczAmQfT+dVPmRtr9F/s03c46gcXSPX3D/EHROl21MVjaptRm/lAFzU2JR3vIcBrSyn9KnB+G8
cTUA3hZ8VcZWUlsE5EU=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KDe/Bg6fHbQcPjNnYiQKwKjMy4sdSqf+Gty0JJ0Cl1tXsbqDCM+FOd30mp8wMVyuqAm1Cs7QT211
JO6FwTQoTSe1+Ag2KZe6AMFgHaNj0EL+M24h7wdNN5Wj8M9n4Zw2cVNCAcQuMAGYbxaWpNTrYMXH
BpdQ50EQ9/kLpocWC2JhjoxshWpofJ0tpp9WlfLUPTm7TftCudU0M3dMNjnbl+Mfa3yuTHWt8aDY
6w/HgH82FHAd70Mwbh6CrcIChQUulExaSON/uCwutX0SehA5/ooAAlnWv19O8kXTawUeKwYKQikK
PjngB0eHiTimSxjDCZaaor8VbS4WfO6DyMwmEg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
cT8dyz0KorR0SYhMOqj0aLFC9aXL8xkJM2yMH1HrCo3usx0cNxJoobQDZjv8vqYF+p+PqyyO+p/q
UJguYwb2Su11/9omuhwbS+PhUxPuwTIKLA+2LcHSDiHI6VpXNDvIlSG9HIu4E4JjWZb1fmLagent
yOni5fUREZ9wL3C4dRqfnEtfA+jm9dM5dWfOiDtTmFXmF6RM/LOQaw9Vk4OpEjqtKF94VMab2y4h
vZCuMtca4CpDODUlYomFAELmgMnXcFuen4w9tiG66QZ8Qpal+Suz5+uTUJbX76UH/uGsQnTWYFOn
VrKLyYRI1m155lfgXrThSPk2HF0AQZqN5OOhb0UEzdK9wrnGNnfGL4v4RNcvl7mRkYPYHdi2jphK
QAjRP4k+Lhv98u/zax7wrAk9vziBaEUJAVoyCnge9aOq55zYdl718moBJ7PbL8u8BrT5RW2nZuwj
2pbioIEkWQBrxr6l3osvfssDCthSi9C2BiaqRaPUwP9Udecas6pTkghMnQFU9LeWbrngxycGX/Y7
NeMKVVIHeJPf+tOwdL2fJJKrQgEcBu5MjCka7ZHbRQ7+XUEtWIRDop3n15SFCquBulQfBsZEB+gu
SwHTyBnBjYNfizmh6IlxcgEw08oBrovwuOCdKZ2s7dH8Pg6Zod9Sj/3l47UkU2yMGcLMJ5niPquD
s4wcIcmaXDlOXADF0FYbfjo1PZR0S+z3X27rgnxGmPuM2pllCvBtrOhpFWPFSJabg4iVgmg9/s0U
8borF05k4UE7vsIFe1OrQjLFe9muX9zmjFVA9pePnsrCwcMbJFKEI1WGNieGzh+lRZ/fwrsyKlUo
NP8EdJo4KqNg7zpH0bWNSdFUS7iJaMzoLUtzL2BKI5ym/mzl74uLlc2dxXVZVbcZJETodac++snK
FQa9B1SHAeCpVD1H8WxuFwwcHW69/PLYnO4WdF/gyuVCsTlsQuvFWaYVkd/gxd2w9Pg7kd1q7ZwG
iE9Yfu4KKZccb38QLBjNqWOsWhtM/Xpx6B7v3eWb9bPTP9DbXOFPFs9Yrt2g+4++afkMVvVXvHcA
cwlgxYjeM7neLRY32emQ9CNWDXIuu5X+OG7rpQO9osmswbvQ7bD+C3Pu4fpBI0FIz7LMVfQ3Pm1N
Co07xkTgZZr2LlydxpJChChBek/Z/ONwAV8VR6gu6GbwGZw569qFlTzUwaGaMrkIgaXm+3ffQ4mN
iwnZ05hAe5cJ9l7e9yn+OZrFQTrhaEZEu5ZC+ty7iVpHJWymBfQ2o/GwcL8AcWplO/yVzB4gbNKx
64thGbli+62VnCsYNz/soez6UgwBR4ErQ1N1FZzx3H/Q3DHiAX8RoKDfAIQofwV9j0fLadghPgGy
rek1sKaWnU+xckNG7sfrtJlPJ7yMUDuVR+FDLPlpEHSUakamWjj1BJGxj1EZWWQ0xQx5MbOa9dwL
HLKArtfgMOy0+x7mV4LQpGYXNfLgCuc2+Lzza6IKnM3ubbneNqw0m0eU2UN/yJd136gUsJBrI+eQ
ezFNVjBhYc9K+dpMiftmo2t1iMxSFYIFbRdewQOKnY2vUtyGoJNmA4nTM9lBUWw9PKCQnFBt/nfz
aRuMnKqoPtp5jQ9gH7Kp6QVr7VOq7N0ob3zYRA8oyN/I6Va5WtU371qz4jcHxbvvWGC5RVfeM+2o
1clpdr0TIXFE2wJScQt5+rF4P6swQ5E4AJtLwjFLDBjJjE3/E9CyoX9d87iEy0KqZyVcjcA6Z29p
x3o8bb9OssPNFSRMNdAJ3hcPm+eXKoVORlEilqt95LcDjB4mVq9cbaidNRsutqDJ7Tkf8ZnYaPp0
Swc80RZsny/NOzRVxyIBlZT/Fk4YLEqfrpJfw8t4xEPPZUeE2rlYTzVy0W64r0RhUTOELOdDF8DI
w5Do9GgZDrNxrbT3FKgiV6SfgMB1plvo+/dswd2ti/lHfNp/s//wOBxMl+tRy8LHlPCBEYp0hdP5
pNg5b0mjd4gMk0rFndcI+TJQl/mGR5yiGVdvAJPt6EsMmxrTwTJYEVBeUTdt8tQVqMtqFfao0zZC
81Xrx97+Y3FmIkqzF8a806bAvnEcKpAA7lo74LSOTCfFidwbjy2edHEr9Pez+JuD5+HG1Kk/xZxO
O4bS1Fpb2Ybeq/q9lhZdIk25ZvVog31PiZVIk+yh4PCgWmLQ+stV2UUCBoyKVWm4CjINaqwURPnV
9sif7ABOFy7yGPn9fo9LG81ZA0v0aMsNQq4yV6naZruu8xjzF7qWkVskvXWpwD/h2X5ow5Z9IBz+
gkACrCWAW+D4vqrxu6ML32Oqq7XnUxEYvjr9k1YixLNKB8oEZNtHTBjjM379aZi9jU8tw8zlHGzs
2SWD71Cy5yG0pbELIi9k0Q/LyTgeDpMSMPZP7XV993B1mjlD1zv4xD1KsRqCH08fmMf6bhY9HZJr
uB/jpme29AKsYJslSFvdPh3Kom32ldboGXR53LsNPdb35NSxQ65IU0naVDiNr7xVQLd01+ufKm/R
khtbtHC0QO9gFhwdImXi+2JAgLZ4qUmtNzeRuN0Y5ach5rnl1TtyinU2sVsOBRB54BGLLx6rK2lx
iA/8Sc5qOc2IWMPFBku7LEZxX4C45xmjjsNlWDUvYyGWn8JAjrLDkxUE1doHzkLvnZmoIxi5nSWs
tjyoWN2mrF/MigoBb0Kj06Bj+CXWqVe9sfIB/zGmQEl0aE+we3NeIta2OCcUYDOozPMM5D3wMYMW
qI95ED7/shP0ak2BMlz6YHe2yLhYcJb1TRrrdAeUTIevBR3Pe8Qd8CILYNV1wKQFon1T3NVhqXpp
7UlCB7zH6OfDFAmTu9SJi77qjwc0FCMsV61c+21JaloOGIMwCS1aX3GShWieQ7p1Vz5k5LO/Wfuq
4daWsCM0K23ZYihp3wWPJGOCwJOjeguYdoammKdGKvn4sgrI91GLI7ZncNEeBPK02cTLatk0ig5k
glyJVkBMvGvynA6hIJFf4NyhAqmvUo9ob/3ZlwGjXntJCsAmUB2oDwd6uYu4U2rQY8lYDPxTVxSG
35dMBcxxAgARI8nq1SU5GUztJjR7n3q+f9mqY+znI/wpU5HHZ8SbNsLsm9LT+uimVKnJKKMgs9g4
3wMu8CkqUKzhKWwl1WP2jIznD/jvlrUFtJcOQ1KII4VXblvNvCVaPrXX/W9xmRlM8UEtFtGvp5z1
/satzoob1/X2SyMd6r3ZbqA1ikanfDkGZKd86j5hz4jChW8tkTq1Pa9vpNELsU5jsws3giIrHzpE
VDOFloWELMPUvanZeBaEeum1iLCBYwuicac/y3XInSRZUM0mXm9zcsUmseelUtiNZiHOwPwrNzeU
UKCi0GLLvOdeHKgH6cV6tRCFW1mEhMvvUzizY0dAFNr2LaRz8LBZ5mZhTpeD/3wHwUxgQpFRyZ+Z
W13Ilf4dyBR8O5n4zCCVyzeAIIaVbTb0fK8bSQA/yNQG+o4rkzTvXBLtOcVShMT6DhmMWXN9yhfh
BJS+XiIk3XFf1hfnIwqyWrzDmmgESAfWJwW/q3TNEVeCmFEuxRKZXDy9LYGhDj/izwHX9fPSaH5w
xzEH8neYanzGSPWk8hHNq76IuREmIIqclTc2IOYYuAl3r6Usqp9zlhqtKYypZnzl7Tjh+5hFx5Pi
KNb+xmLW7HPPOiksOm39L8b9mUj/BGgyJUqT5PuQzoGYA8sWgVqpKndvYqNUhh94uBuwgjJzUsev
hLQhQ4MbV4GDQ3fisuLs6xSKvnbeRFUmUJ+HgQ+W+QU2d24uuHivkpHG6GU6M7mvD8NS70o8p8VK
EXPTQKPEqJqYCSLm6R80yao22HxFy5wtxNdVm6fojh+oDgDXTqzdxbxkKiVcHoQcd/hBo1p5zm9n
J2uArBEVm+Gq89NP5aOAf9TMm7FLMVrUrVjpNxz0qo1PYCOtVR+34TQXkfjg9hDHQsR09VFaIrfd
ums52IoMHQvMYWLZuGCGlVs3DmLDfaFI9bLnRXO9kORbb3zGOGlr7V0r9xNm3ul7RmcFKOsBK+mR
HQUJorNt/Jr4Sx+vNeXIrV8js7qKewofTFteAv+CSf6PiF3lcZgJrggq3jew0r8PJHEbI5Tr/Dnc
9Qulp8gjXzkwJdbZB/AelmRJwX3bQ5I8VqgbdHifNonTmEeYxNcR9T/ZtvIDOcsz+b6yna8WOKVa
f9nRLWuOKGYFyQSq4abBEFTDT8T1pM8OQ6tSak9y94L/JzjL6Q0gPs9X4itm3O27zTfqGNqa+DLC
0IR0atOgBr7bIbzvZIAIX37tMQXYqdfiGtugqv+xygv9FcWv4QttnfeL3A+5XWjMMj6YY4vGWuFD
InhfNhBta/ILI3+WhobYuZsM57HVgRlm2tnKi1wj7CkSVg7yZHasV5U5+EvR4OtHe/thYUiBFHS2
1xkVKxZJUHB4DvAsmDDv+96RhOCLj53yEJ98ANWA7PTJZD8lCKDNjjTNwYxA+0ZYU6exxGXfakS3
V6ZE9CD4Kkvli+lVcUGGBz9X+KC2kS5xYB5KSPPMiUixZFed+eWVrYNCEDr8hiB9NiSbwb/Ig8lN
mrzen/3Bv3AGXiaj5FQ+njV9JwXGq5alSuHaqEYcUOc6mThoqxHxIJ/KVwq99axeF/obmtu7ZhW+
7qmHufXslfbKQsGYD1PvgiXQiK0v4XDjl3akquFrxYjAEW+NU6Kg5iHvb70sTwn3nqrLMZZRll0I
XvvnQ2MCQKMtS7oPjeKeB8om6nWGxEdw8LfukY2/6JH88zXfq8QbLLY1dw/UReuR1RigcO/C608D
CVP02LbsDmJjPKduRtUNwwvA3DNmsgJmBmaa7KNU7FFWJe/fwlFKIWiS4bskUXVdSHBQ8n/5PZqy
zR7pAorkYHNkRdT3LWRhOQyqoiy3CvZOG+P0hnIZU5TwmM9iBBDRzQnw5ZoVVErW2IxjqzjrHYXy
taFoK4HJgFbb23lq326Rm8R9JD3UB8tuRKYjmjbzFlOuZUUl7hqeWdYlcjmfK92rcGZl9RCplzrs
j/QHMU9M3vmgUauWswU1nWUKf8EeOywm8ro9oKBwQMmWU9V5x/P7JEyHFazEn+rEH+wjgVi3lvu0
kJfaVNk2f99pKoYIAArbehpKWEQo/KG4FfsyZYcrx9AUK26craFAlui5sfyQuHuk/ztr/EWWvg8i
XJI914BXt48REB2q44jQOv3cMKQuSrZzh8qp8xQuPT63ge/wBQ7qZxC8vQUhswuqAUcepozcRi0x
jqugZwSV4QYQpDnFYJk7ZBUyU+xvu6asshO1hAPvDvMd9ow1pPvmaOh5Zn3gOpTzz0PWjjUncDcG
I8Sz9zgL1oI9Lcbr68Q1OMD0lPzh4X7EptnV8WtmraYG2CcNqWAbD5GTkkZmmmXAwi+NLY1csJpO
s1I7T31HiMY3DxEEQUmJyAJc67BHu+NVsrAacu4UDJUjYUP6Mh45n6aFVRu2UvTi+B6uWlH0gGF6
JiWyFHjqh2qHbp3N2zVy4xSRVeNo+ZPll6aDBo196oClX+aXpxTNzj5AcsSg0iQ+KcCymOb9/MK5
e8/PZEs6rp08RnZDaEPQUDAjt0oWu+6xF5VDY1V7orGMaulfD7dvMZUVwrn1iEA1qZtybc3uQOyg
LUwYk/Zlb5W3bDn/mB99olMvJe7uEC30pit6cTRBk6ugl7lMqjlu+Z4RSRKJLT/O/OIA8KGztDhB
SXWs6GzSqukd0uDuSJKNWE+BcUhmea1RZlSQBslcnyI6veiNL/7qjhMZxgHHnXgib6oofNOC+APU
taStH12Kznr4Y+h/6NpkK/4NKfhKdNAAi5czx0o4LreN1QVFaQv5xU3rXKTmA0e6zoHJrgriLQoc
e4v3MhAoXhOiwAX/3BwfX1xIoLRXyU0C5AxYuOl7C+e9S4CWFiG7ZwR+xkiqNdnLovJEahFDPiDy
PEImU0gNBmgprnnQ7QwkBcYnzrrxWMIW+Zjo3tTEfaauXwdGcaMg0UzPNa6GzvV8N5EpfPvq636J
6JHOsaypVcvaSSh4objRKe61ij1jElmHngmfWDMOy0qfPTcy4XOmUCXg8//NmyywMetRKxztEqto
HdTD5Cnej64JvVjh/PgOA+vlUvH92glyYMDYicK8Q63Q13ducezHW0O/VDxfbFSfKdannjerkVkd
j68MhYctJF8eKc45iDHnFeRrXqouwvR3Hojdrs+chrQFYEcOM4eo9GzMlK+2M7TikszmxuX070Px
vLG/cXA2rCYSmmTcsWPw69eCMsWHaGtwpTn40CX1PdanoihPQD3hHDMHQRapnW++OoGuZLJLknnE
2FgXFWfYcDL9Sm/5qBsQQQVl1N3TH6Xr3VXAMqEdtmip6qRcT7Qbcn4q96K2+DFRcPTxQt6lyKx6
aiXeQ5UMXnVUqIrMxdbxT4jgBElmUMbShvEp/CyvR6dof/SGBjDC4rq6d5bjXuY7ztQYxZtlYWV9
Nd1Nl/Ihp7p2f7W3JIYTymsMD6XDNfeLlgCNca92P2OkAbrqqM5ItJbssnS0Gvz75iNeXt1GY/yn
rCB4N6ybd+4gbDHJmXNVvt6QAjjBebmqLqAePljDmb/2vmkF0Ix5QEtv9Gt9NNP0ldJ03sXhU5KR
78O7tQ9n15Ue857iNZ2It0hzAYyd/VRlyaAKvhRurJIIwtG4q9FLv+/Fp9xd8ytLCXQnSesorkyM
q3MJ2PtWmyRuTCN/2w9JAOrQiW9VIT/voNM0iZ40hzIuTO0nZtHEgclQlz95FGF9dizYRsw5SNVB
wc4rQMkFI9w/k2KCy2DCvDD/OJ18YkDmZfWmuJa11xkhue5SV+FE1toBB2MEEV+lfctUd7fnVVKe
Hi8gaN9XcszTMmBzcZ7CR2lbHscB2Nm21kj2x6UOZXnez1mMkcZ5yjuF7NJfLOm2Whi5emPx87rk
xWqdwlE2vgTHh/3OTbviC1maBhYNzp90pvwni/zdlq6yJVrxwJbQ8E5LHjGMHNo8j8bQvwWW3Rld
sgKzDvKlOvgHWefjgFMYgVjoksg1zyW38Y5eP6ys+Eq85mFkas+O7Nu501aK6slbkWS1Xj3dAOVD
FQJnEyCz+nU4BRJqcmFZJSFMOmSIb53u6Kos2Wd7nOhGomScwsEpC85rvp1FAxSbt878Ll2/R5/Q
qkCUKIa6uV++XpU7uuwsKGCLVTilXljLDDpmtViUOMYwlzv+by8jy7W2bJQTa578qDof4VHZBj9+
uCbCjCdHZzr34BYcEHJ9x/aTpb9sAaIsWN9GPt34ulQUu8162194OpZwVP+pupjStjolmkLKTwvC
bCsPGAPbFbLH4mguA0iTYGzEv/jwuZiaXn6yOOwp+gYEiHpe+d/0ujGcEu0/tjUsR8DHBuGTfKW1
2noEOJN+9SUuafNuz7uYIdlkQ3yA0jQ/QiLDzkMovCickRB+fETaxB6Jc0N2uyjGdYkqOdc5ARvF
BrBTkg+Y/sufuddoKcIj06IfR9sHTGwVYWm0QsMBRicxthpWSj9pJeqCqOZG0IhQzFPj2XugoB2c
cuWAd4v4Fw69DRmXNmHQKcrHtdycsRatsETOMRwBwj9MKtQad4Snt19VCvJdnVe01lGL/zaPKmvl
gziPeK5hQoo+fJ/odN1bhZfG35OJGdxfBLTTl13k7kcNftf0r9AEUt3hF/vnHLhwa4jnyPxV0iJ1
5woVTdTeDP/t1/wCwTJ6Rs+22dmVsfCkTFT8ypW00EkpczyxMESlYqlukFUMtRG+xxc222Ksk+bH
nyVui9U2pAzJ1xxvtsDzEsOlMQ8imVqoggh0HTIVRTCv31LPDggrUhGGnuZl44aNeo0iKATcz9qY
nwR4NiSbbbgp1tQ4oZsMmoNlTaxiYqah1YGzfqWALLEgEpJ4YvXnUaDIrc3crAlgClo2WcLzNGZO
x7siWcqcP8Xtiz9Ophy/XDBjMSm7pCZa26XCcN03uP+7U+OcTUJdJQNHAlvOAyEy15P3KH/mAujg
Z7NCM+7vSrts7qdpPj3+fFq6Qoj5SOOX4xIA3uV9jeJpiBS3YuB/tc1+kiVCSFkY4CCSpxdH4uKX
WBb/2FF5jHJQQrqlaqieUlmkaNvr7wJqKBhqHMFXuGTmver2vI0NVOTaA0kSG+yhLJ87hmDNrzWL
NA771stuQfigbwXFkkTh7Dl/j5KVWG2cakFqg9ilxftyr/ZjYRlR+2UCDH1GU++K/88W+I6XnFhs
Gd6UcdRDmUFvIt0EGAcVg5HjINu+eu5d70UzJ64LcHkZDsWNddB3aMeCxsuDA6NXxnlubuzHVWrH
VnMSihTqcSw6qxMNxaJ0NMakNU4rqTh4wEtz2O1RjfukdJJbdtQlzmyafGCvoUV/qz/aNMjWOIaq
FV64jGmhfHLwzI2mMzEnjiUIrbZaegGbttoKK0i53TVwstJ2C+A80D2P9Jww6FSThQH2YxSgtJXO
Qs714oi64gz6PIIUx5IiiXD0MJZ3wwRwlr4vIDV6ChHqvSGX/BbXuEydsniZeKPeuGBSN0Wb5QSP
j1UUMYcVgDZPo3VfheaEqcHp+1udLM+1DlN2WnuqwWgYz8K5b9e/olDg3pQnNdjp368iaGYnYjOM
kdZY0lORs92ZgRiuGOUa1UctEfP4nTQIQy2Ikne47LmJurE0iB6nzudxLx8XUpHoDZJU06Vtq82E
zA1HmR6ap65Sot/1MWsxlLHOIGU6LgOwHU+Fr2TDcwo6BCIe2f5S1yBxLz+i2ABJpEAtl6dM5+8V
HavJym2b+2oDRkA5QOzck3t8NWtsvBbyBH7ZHebwyrENi2qEYja7HidiM6ynZurjSJLTOviThlAS
CVHNkkMDk8qd2gHJPN5k2y7MTO1KkGVZGXM3k2Z2ToqdIeVMIXhchU2hvDOLMzzNDuQM4f27JhPd
wtbnR5HBALpWRs9Z9fw1qV4BQbSIAgGSGD0mbVIEfvXw/7KldqgnUUZNdImFQgoWnEjhG/l7FL9T
ZJsAuDXjUxInLDqoLiwUSynZFKl3ztuzAhFDe7auW4ZiSn3oCNRT2l4mRy3xR9g0P/335FWiAHpA
ziQXmbFug1/ebtTkwkaIuJ2VavTyi5q0hknICcZOYh+vg/N7g8H6BVkzwDvGwD6Bw3zcaaBVsz70
jNtRfZRDx9tnSOOy9w2N2b3sWKhGB27flRnumynHVrp9oJhWNoM4Qz9HQvczrFaviWmGolxM7jUt
WTJm4GU6zTrufA5pJldogIowcA/nREBmtw3Iqi1Q3YLSVfEhwCo3/XC+xC6aVQpMF4f05CHQ+pdD
U1N46Xc1GzqrBmd7RcrFla/XTkFREBFhVnN5yOkZkoyQqSmcnLVeUjP+h6HgUNrwxA0dn1e5xzgE
bUDljW2MTqvR7pKuiRkhcPSrRUxxA20mTKXr/EoBlooUCOdUiXtu/xjgpR1X/D0eLTWO8YvIhn0v
iNSjXbndtgJd9H/WMDc1MBSs3w6wmxsVrv/gvoYomG5ILOXEtCxInrBtDPcD8egy6yHY6pREhlkc
8F+Os+ZWau9CASAWaJKQWxt5lEXhKTmUMC1jnjxR9N91baICxm1su/W9YdkHPxKuCOJPEkSNV9M1
F1m9NiF5P2XBPrekl8MBNZn4cJYGgRYdgpLhlvnByZ/4Vd7i7XID/kXWZ5lGlU3QgR1GVKlQOklt
cwm73v6wmWEVisLhkmAhNuHT+idHLj6+p35CGRExRLcSXMQWwOQKKGyiKBbDdGXgbtU1BkwqM/c1
UPfo8CV4hfgKe3F+NYgoTkTdrDlwhVuU2oZf1/rXO5Iklq54Hu2QzSHVgjINLP1n8k8MlMcup48P
QIfDuktpav38tmOWCifRSqFDp2vji+VXneAsvSdqBd5kSrY0hlVX3+msY0mWJ5lUVuCRGAC1LJ/u
kla1gcVy0J7X3Qj3sXS/dsVZqu1jeM5++zDF7MorNJ1zFGWOV0r7KHFwXNqJwGGyvuGGdY3v0vyt
EnyMdNzwhLoo4x1QpBbQop6jlIjTx5wKUVHnJ8JScpkCdfrCm+8djARwKwljoFgH8CsnmbxzxXAj
R+b+n9J7/7jKwtr311tM/r032divYgvbmMaFSSf3T1H/3MBkjomaFOkhcKglBs42InRb+P9pSE46
BMoVelUqnoFMvCxSCFuqm8cdwgY9vNaIBFfCj1+UjXNg/HV26exiM2SEDNVQo5S8iVF0FcP0Y6My
RKrYS+tDoG6ij+8itc9RyIrw6U5/82NSGi1XCxr6QVwtNJwxxJQ0qDrG7Fl1jgUFRZsOp10Ww/+3
hkac+C7JOdv3roftum0OQEkbzJkjUf6UpsZlsNH8zUiGmjzCiZmfP11f90RMaFO4NT8ZHGG81Dyr
CiOH5Oiau0hDTZKu7NglOpXLvnbgZ1Ov+aWl/0tqaFGV1K8vGSxDJLaDLtI9KV+paxM9KEP36Fdt
+np9ioOvTXo0+Tr31KU9uW83LzEXN1GCCN7NwmYvc/Qdfh57GHfuBlC/vvzc/z9RnUGgx46J33Bd
u+7DK8YmV6DCug2opVDLIfNsQfPLFX1jXwJrXgwCl4gGEgEdd56vHCeyt63X4eDrlnveP3Qi9TRC
mEFcFjxgUWJhn3ctUFkmVrrcniMRQauH5ejz/0zOugPgldVjiAW2i0IxOnQQlvVab9zhdpOUhFni
svVIhTnzbzoHbLAtJBfWSnBNUy5G1XQV+pH+dKpK3h7XKrZEQlIpKpXdOR2Dvx43e1pizvb+OUzR
db2HV/tHG6qEY5qEkCrUmbOUYJBox5G52HP7REz1c9PuHEEA09JVaLbsG55c+hcIKEv+5z7vmyZS
sjNiT8hdtp+mrTXQvqi7VToqzySYLIpTFlxSd1bcTvE02IfSVq7KP8oC+xJHNW0uyBXBWMpdtroB
w72SXY17gOEj8iRGoHPDrx5wOoXweRp/37xWUMenixn/4nz2Eh9UO33jEAuhmDMcv9ZB81Kf3T+D
8JZts4ePJC5N6tzqKD22/laxdmU9DNGb6GWm7NaUt04LhDp9uP2Y1Vu0L0yVh4LGqGgcpo6pbbsm
V6W+WVQ4yEJV6apgpHXQzmDEUbgfFlAzTwVtHc0vPBaDd8kOIC1eIyd3GSfN0alhA6fsQGMJpV1y
l/U3x1Llw8976SrZ6tKYKUxwiECvHo2scgr3OwpCrbN6OY6jpTJtHalsIW0FsCKl+NT2M5WItTP9
Of371xIGpQouKBAgnRf/FnZBzola1wzKx6JbkT+2vc2meE0VSu5WWhXjKOCpJIaIV27q2t0jt4qr
XPvBeGx24GXJWPa1NvDySrkvCcCJnrU8YGlBEkf3FSodQtVM9Q+PwnBKoANosWnmXfdduxF+zQFt
itjTeVldcx+conFS+OeORQiSRqeuBPETUPospgylLFi8M35CBNnruq9pejmP3f5CQ2c+W46dHBCP
o2yByIPwQFkUXHakSHSM0tHCh8dG9yn8ilyshn4crrMcw6Be97PUmzAwwHYFlKyTICptfVTfImnF
XUwH9uh4yZJvLNuYNdYEVnU1KiLIjwIQ9nKSv4ELThVKZjHACKuobxxd9D3M11pqTSnMRvI1+uFn
laEXO4/+6mxr2CaYP5gFX3MDqF/CLXdSIBNTuS/VQqLxQti4n4bj1CKp0YRLbuhpGLqEDwIb+B1a
/Xajx99YcrDiPY/qHv8Ua9JdOpHEg9IJafbk3Si3CsVk3IcSjwMkeFtAqBLVY/Z666nYGwSyWd+e
k3UY2k7DT+pw5gPdnFeRN55OFbBHVyE+z1PGi0/z+vzuqOO/Si6iOGJ/rA6tloH0fqU2+V2lVREp
BbNEU9gbTDZw535jkNNlwJKFSC1vFaStZjpyS+t5bsmZhHodKL8pdfqOwFG5J+NthRDx6+980oBF
L+GSLa4ZJ8EYlTzvEdFrUBax6aOBclt5NnBFmXrUaQ3mWTB8SwoE3lRY+v181pGOUpRA25DYcDAv
xYoTmBRJgJmeX3v6PkkPAvAcrENxpvr3wp2JhxwLTTzBmrq5FNRPofUEmD22GYau+/ktOR5xY1+c
wxzohqucUwzcv9kLww6b/LHgsTNnpYj/jbf6MtITpLGHPpdNAulSmBHK9U5t6zdzX2bSUoNSbaZJ
Xr8Qy21AoEHgRLzotxo5TJpMeOImmSYGg62mD5r1lkus+OYTM2L1v+Q7FqGJOoLyIupuyxqlGsuO
5B1xdlLil2ww1sXcuDaJCEdWswwVwT3P5cb4PxATjCCMPkCG3zD8dd/YHHpleojQIkOXDi/PgVeu
aQ8gmbkBc0h3N5gVmb3ksf4i1V/cUBTycvekGFKB/d05JdDmYEXuZNHoLMfRVLBBDycywAOyPiT2
FyxwyDepRIHliYqvtkad041uv3dGMDHOtUnwNAhsMuTLv/kf2LSXLxcjyLTZgXLmA7AXdJUZqsxA
mBcPO6qyp83oR+7FNskHk+0q6MJgPqyum+8eLksullvtTnox5qB5XiIEZpAINasePbi4ybiElQ+W
ioSNXVBjTQnKv+YCjJFVCMaTxzVdzJcaNH/gX6+Ft7jTJpG95yTbmUIIX60XFYl4b9RfnoaEAYss
qQ0tX2MVCLAJHDhuzu7MGv6UJsP3yrq/Ehbww4Fq2lM80EGWmpQBvwSjsLh6yz2AL/3Ya1YZenys
PmvKMUjuK0DGwFeVLGBfn9y5EwMfF8d3piEEJj/HeSBuFzKZSZ52NaOsHQc1Td9MkfY0Fbwp6ld6
gzmjXrB/XAULQxg9XgkFl+qdpx1mS5GTZ/v00umsRugZRYFAOi1Bp28tCg/erlZKRm5rlFfoFYEh
Je2ypyPl4dhZySRoAXpYjZ457cv/vfOBBjbN4NT+eYBdG7bDnZFOYyGtXhORYpeDWW/DPzmu1jlq
TpGElV7PUVUKk8Yg3UqLBss7z6EFE6U6PzBM+3iiB53Ef0mAe1QKaLSecU4tjspSVAi57VUZW/dN
b0+mKfzmcxAB0/ieNzKqQZ0gEGi7Jlr1X4lNm3GlcYPUPNzK9m6k4ENvKrE/BnYK/wUp6dne0Ruu
wnG82Toeng2KGQtGHMiaPh+PhcREnN2PwbFpHbqE6Dwygph+Cov+8hlXqwP2b9bPGQ0zq1o1LHiu
oTdUhNtwGfFZ+89O+s6SEvoTsYtUSNnYwiUQaD/0ddovlJcH3vFMA+OfnGcg2cLCHRBVW53ZHQVL
l8014UkJIk3Ku6KsYpTsiKNgpDMGOlr3dI1fwQznfe4BMPsAr1jThLKzIxbIvgbtGClh4hcb3SRc
eYKAZerWu5CqwVA0XzFcQrSlGxGCUxPBGUFjBCnNmzv11d9EW3Z0AWCaQ3RqJDKUooA6Rhypuo63
c2s4rfEv+0WGY68vnKk1nUOTZd61xViBDWvsaB1hlrg3jgsUj1W0Oc77OGwuDCzQ0XliF9Kl1PIw
SSO6YICn2oj5tsj1Cmp/O9RnypN4Rjxphj0eRIOzRvcC0lYbbjsb8ZK2vQoog/N8H8jfYcWYqk+f
npf1yzozWepnh2RmnDWpUXvjI0Qdv4f+VTBspyfMiXeC3TbXzRvbsl6Hdi/zY6KS6L/wJr2LSVXO
kQ+yisvPTk2Ar9UCPtV9uqKjtJzXmMVrzPYvRd0nDGYC+EpTGJb/LlNiYeqOAltGcUYrIyVsVuGE
LrPAFVdaUEj/2zAvUEVMwgrpTKSNLqFStmmmUSPT9iQVQ5pBSq5gPcBR3fkyjkl0Yt+0jTmdbecp
5bdkljSaoCUNxhaRuQvQ24nIZXOi6gke5HQvFK+qRtY3A6Hyaer7/r85Fzzy1JArxSKBkXCcn0v/
KJBAwSRmVBkY54orV+8YHXqcj1Mu7Bx8qQ45PcXknCLahCBIymg2EzYV+yQ5/Xa77CLs7QBjaqoP
X6mQ39Dzku7Dul0Dj3R7TvW0dpDRtLMpvE8I9KTrsBY9p//yRrAsYhIO4YLJp/R4Q9QQtzz6fIzz
E3eEEiX8BaC6iGCYSTZCqcJvllCWSyWaofWULddaEL6UEsqw+rmoUPuM6rQ15bomT4IEtSNCJFaw
dhSEOjJNxozhh7DLq639AYW6Oih1DeSINAIIgpj2LPqGBYGeqr/5BlYdzsNqHPbW9w6ABh0siylT
KF5BmmgZUsiimRRtFrO5qp7P812iG0jqr/USoAmsalb5DNgnZeiB1m1okd0POy2BS3IUEr4BpMzj
lmIQq+zydSGNGEG7rvvBsdmlBj1mbbV8Y6T8fMBxnT1gE+ouwrXOuQgabyCl4cXAWjiQxnx074aL
hO4lzzbqOBK4v5ltSGpcDAM/xzBjJ3FOVQzsqjSeBZgo/UHt8dKhKyLSEQ/uRkqY3QMn9c/w7obB
5wDi0OUglOBHojpK/nj//wpKFwczDcBFrtMmn+7+3Vt+HGNBpi3nz9JsNq9Rhu+N+7jd4HSVPuxP
uwku0FbExkyknOc05fT2+yigKNLFZjeImuUudeuZe/942L8OSDof5LH6i4l/Jr8byvetCVFmckM3
7nqd5uLxh+crC9dst4WIvhtFyzJq6N1mbzEoYmLtYLNhMqhpIrHz35g3rTOM1/8HeYB1DQtxoms2
O6WhrbNPJwE2DNDTjN2ka0pz9WUh1ssvgP5SPvofsuFti0+SAusA57bW/anjiUgClaKRyEvT9+sB
k5V3vjyN1s3B9MFsX1TsNxD+Zwfaltm8xjXEaegmiKVN61oK/YPf68CoCImQ2BO5UlYK8AoZZu0o
y/2h6k2li0NqvlDi3fp+Y7bP4ORSa9cbCANRaGSb2cRl5XHblFdSin++LHX+XUNi3OgQVYkXGiyY
gOpAkKz7aZunPjv51iyrxOeNvAy9N/x1PLUzTTsjsizY0HJOK1Ne7JBPXt9OR6DoEsLD2bXzjqrj
Mtt8y4I5UGQEpzwN61iG1cwmGOAddsgoa0xl8QvkpqA0Si4IDnrJ2sH+6QQ8lmCu+0pp6WcQaJo1
KVqCrLXij3BMyDRFqul4t6Tr+7+onynpHgTc5Vj2TaQz4yp6B4DWU0D5ASqi3eW3hcYQIt+UPxFJ
dmfWcQm3Idue+7rddDXu6ILb4Tfvim9iTwRxmpUSWxAnAz+tWjbbZz3NhihGw4+wQocT57kQjNDl
mDzOEhCIRzGA6W6x/Qe4XQLE0r/SICDMS8J5EF8z1n4xxkk2RnIQ3NnsjdL9KYygn9x+rx2c8FgR
eIrN5p/dha99SK4sHGqdI6i+Ax9F0nByJaTcMJ81D2CYu1KFqnScnvFKoAdjlIQ860rx5p3tQoJy
vlj2hu0IN7c2VRgFymLGv7PaRMZjL9LhFeRkCOWt+j5SxfsXnSh8tsWE9Z3AkmLD3eSewBeTb98A
yAR5v4W1JYrXTvF7Dpq7Oe4Jx8wCErFPyg7gwWesAANPUagUm9RXKVB3ofw7/inkmBTDYGVNKopp
sizdn2RF7N3bWAemhUWNIH0ec9nk0LCJoYjNdiQYSdp8xCnO48PeGyIXPycgQcOKDxJ1E7VTvuuM
B9Kum8FfRQ9+JCU02UYn49smingw3ypeusbgJdW1GizAzZ3ZwMapAw4ZEk/8s/vJNELKQES5A4IQ
J1DTP3JFMJp5wT5RPXHP/M4j5B3hxQKAQRYvR/y+J5dKhUmipEYbFblHh6sFIYHlXzWmedrz5NlH
Af9CwX2s9X7+eHCX6JrqPz5iEpy1IqPmu0xpworO5wt/T4FAtTyzMd9DQO5QlHjmDGypvhtGdG8d
U46kHEg+aMvAXg3qOMil7RKs4rQyYqwpH13sDcB/WV/SfwhnxojLMGYxocFmta4IUkbYjKeU+apN
WgMf3PAuQxyWx24CFi8QWp4C1kSGLXI9P+T3XkOcvS5yyhqXzBQOW201BOgFpUIinZD/usWoOyyl
2IIZ1ApVkqPRJeoWdo5bfi+aNJSGXJ5mE4Um2SgQciSch8PTq9egFLzYg5eqET6GdmjeLCwz5dzs
/s/8Pi+VSb1sHBOaxWzSrRUNsmJQ4OWzrwQidZL4CjdWQ5lSDueOiFbN40pqwSRl+M5aCaw2q6ZH
ZsffwJJBcc5zuNNPTn8BrSsPybASx9U3obMMZ380/w40qU4DJY6s7OpK8NCcCdeRX1Y+lhuFi8Au
inBvOYuODQDHaRq7CiEUFaBiLWTsyKuN1eyMJJQDrggEyB5dta2zCFYEAJxmeiQd4jCECvXXIrla
j/BSz1Lo/6Rg2RdKppqwARQBZREeI17nC5wVCwIsSxem8eNV9HOgRUSza9XHJ86R+ESrjV//nma4
tN4lIKweRRHZxSTq3d3nj0jZy13ZTVODtEivfXmLPvpkGsP2n72+xrG11nx8v1AzwJ1zgw1+aTwq
pD2dgdaPD4L1nc7UYJcIx4zzpIEizAmkdwKfeAqCX7PPkkeW6xWqbISIDhvD1j2wHdokQ/H66HM+
fbP2ZhpH+wfWk/YVNt37yjBx0SKOEN/DzEenwEY211gWg18U4rIxfc03eui8y+Y85UYv6xpxRzl9
4ARvGi7yF00hwFRT7VAB9R7XEYGVPZht2iZlOqAFbhTb59PZ6rVxDWFXSthJMIsLELqEqWfk6yBw
uEdfaoBEQV7iMCVi4ZTFE2v4WWqgbOOqgeaxg1bEvEIWbTb8dWsuidk+aRJv34W4XikfUGheVmQi
+CmE737G4xdPzNkeEkSlfurerlDR3SzHF1gPGfQOvL/cfD4IwdD+cDnCbSJoPQn3pfsOP1eAgRay
cfW/Sov2fQ35MO08xH3c8j+QZhn1iQ66Xnc8WjTkhSjru2RPKsnLW2itzWG3F38p2rLryE9a5umn
58EcvjISEIOqjjgY7E/crvhVQjp6DoVu+HF6x7Wx22WqSnaw9K/k/2jMzxynCI6zCmXoCEop4XFI
1B2xQOTrRFEg5TgwcMNvwxHiQdceGYW57oRxxHhw+a1T4+PZfpQ4LclPpxu4RVbIwdExRW8QzoeV
XQGgXBY3S9LoWb7Q4pngdNQ+hnzAUm7sZm9+jVjUEl9ebTbkji4VQDSgpz3DuqPxdBPj30XbXveP
V+gPyk2dwr81QkGhId7IIkyQez7Ghg+pbIVKQKwT4au5X0W8ZAWSg2gFnZj6kkuhyvDA2IOyb9ID
K1lHa3fj2Ep32xHKjHBUNyji6WhDYlUMikjuGeUTYvz65xUzPh/1ZXLVvUMfKfeVy/lj1tylJoA0
v1gEp5PsRavSDYjlKRapUkSbfzdPqftNsgzGO4SJn0wIJiJN2ejrPJ/39K1dsblD1ilAz1+ut6R9
k8cytmcnnI9vsegDaLwNV5yFMQ/Ihq6LelgWyrZ2QWkMMo5iX5O+09ZkzN7Gb8XbJwpd93GAuLAK
kvkQw1mzMB7P853W9VQQDbajpkkSPXrUUB7XI0wobNF3CGpdyDtAC9yxz4ZZdRmGn4eJLzDLHx/U
LEfU6a+VURuJ3Ff0C2mSQf8ZoKnNAlEUKiZCm4pel5pHuH40HzGQ4NXSjGZlRs18w2uKzEec+l3d
t9LWIYubKBpfEU7pnNydJZf1n2JbsyczyuSxNA/+/l0kIqukI4DMTZkoBbyl7FfQL2+vEzr41gi8
7EjI+sJlZD1SIx2rtJq5ghZoMD/bYtWPYgjZMhcsGFlPZKL/mIBgccz8fZPuNMWdCTXwZFy8LaVM
HEJZRnj6RdbKK7Zi6ytc2g0QzSr8RETETlB+NnYwmr1xVPGjoHK+gYceFKONdQmgJOiOYiquHFgD
PLOGPI/gzxIdryBBp6pFRTzxPIdqaeSXCQjDJZOcgf0F8KTXiAdaiscpfPay8Ka4E3vScP89pgwI
XT6CYf/SMgY9wAs+8QYG96bpingFCMPdDrSxuPQqfNOS7NgEEELjxuH4ecS1JeI1pJF0TwLuMnfQ
3IIeVCpw9R1UXqdlFjuJD7hCs5zbAda3PmTY8Pe+fHEuJnohDMCOt4yu6RvMMa5GodS5WN7HNkq5
mD0hWf/kL2FS2OEBAxLziHHs6389cshXIZoUs5AV1g+ZGG3tFBZNEp0fBPHEq5801Z1kMgzjgjkR
z/9QmmGV8ejKZCd2Vtzdive3T9Namiz9JoR/EkYQ4eAWN+l9mKgbB6mOqg8yQ/jIm5GqnkpCSr5E
5ARuTbfGbg7SrPreVaBWfGPz0oV5vkXlbh2A9WxDS/xMl451YZZQLlkb3J0zaevHRmhK56938ZQx
ZNpfeGN/xzpUyN5ZgGbUdQBv815l8e2hd7Oq9TORlBPdAycv3pxnVhTXzzYD9Vv/z4I+kI6JeWt4
xt4jAbfJSFYt2UfKwRSdl/FpI+8Feh7CaR+w3Kvffg3aRkQcszeg9IIRSlxl9vzX8TXkODMclNmA
MYdp/PJlXaCIdrEX0o94SdEQmsx5d+PsIaUobLjO42U4T0lsigVt37yzFzDMuVsXx/JcXy7+Jk8E
ueu4Rqus6N538jb/IqfBLYDln7GzsEzvL3yBjFkcRsndnzzpvCaFwqntAiS94TvcFrMjc5c9PpDK
7nOtWopuiCwqdV++YZyP8AGoSBwCREsM05jB/6ZFjiRjNh1Ww5tyxQEasrVFStPMqZB+d1cbqR4x
TOsc1aC1WANLWnGzPUwnQwCGuQ5szrDK3KJXosiQ6vWR2poKiLmjsxG4LuVYMuRzXYkD3FI4Cn9e
131LlR0uAFYqhwxeMMN5pKZuLsMQpyUYhSFX89Tw9KubuoGHwi1amTvxLQx5wB0slYdId0RmJyfm
zYTyG7UlmDBBMpP3Vr/VLrf5CARmFaI/oPky4rXXYajRG1d/wf2xGaGICaB+fH2MkmsItxjEpRiN
xO/hgtJsJcjpqW1p35jY9w5k0XOaU5Uo1Dl/xLMvkHde7g5dDTZJsSbfwDUmU1wsYYDZbqS026b3
o0ERVUGYTvV6VYXvJAyO+od7tLbqU/CmzT+gHhT28r7J0+LrorgpCcCytryPe8ZjgknwJ24MgmY0
JcpluIPC3+bLwhtXMZFUEZB9SKlHzwff1xr/PPeIgliZNNxZut/LHPd3/7sG5N0M9vg7fScCWWnT
GEx77HdH3D01EXFH+j0dxyafDzStrnp7u7Fchwd2AVWY7Ufzuh+hSCMOVcEJCqXaQx7peFC2Qlgd
6U++TkJrkDQ8Tz5Pk8UIgrNFVOejYcleZ72G9PcLOWDt0wm6DC7lyMrYJ2zo/pA++Lo3E/GVwGoa
NK8esYQf5rVjixw8D0XO5y1NDPyVeLaQpQZXibtPxC5lvCVD7O+0GTdXIqfbKQh+3wOLlBuUpgcT
IpLRWPcw9se3JBe9dFN8m0KoecWFJhUyDaTgy6HtjpVLQ9t+ky/v6CXYXSGWAlS+AXesvu8IyTDp
Oyj997dQCgvDnwNR1tGd/ZUJv1B6feQ3sQCZBeyWDNDlrNLPiqaZaOZ4ihIJM11QmfyW9SqlsajH
2GYoIkpxo0U1Aid6igegL5o3+sRtZL6oDLZnxNaKhAzol+8rfmYUhO6fGxWfKMBrNoNFu50amYEK
DXOpsZMLBrQVu6Ioz/dci6+cPMV6bZQeEE129pPCkw3TX5yAy9q9lGqvCDV+E40rTM0PsP69H7lh
jpOZiV74xGLK9a0vk/5dTUXy6Gj582ac1zV0l5jzn3g6rLo3Acj1dqg3EFgcCzGld4ua0Apnt0gb
J2RrpTm2NhgpzfY1x+Kg4u9digmXIprgR/VDEjLNucPmj98/uTbLNhe2S8b3rbBhyILPE7CXk1eO
cGU4hp4Dem14f/a5nk5xDQ8kuw0/Wn6yO0uUHdOFsGTwzYH4CqDZi854QKvlvFvZs4fSHV5GTp62
A+DTWCMq27EeCDYQip4yEpOftpH9liJKcemn2SZeuKXHt3syKnB7NDgdWA5W77LIUkXpB0ufXDHj
JMDIpUwkxRDgLB2lbDGl1qDsv/KtkesJDtMPXWscOqXlxyDdKvaKzm00wvsC6CmUVMS5wDLdFX9n
mjCtM1tX1ugjTQFwHAcaK2VzOV7jG6gqsoANq1VVyAlV9C9CyiN48FbS6nNE9VG9pjpofNDig7wo
JQehoBpPLVWvhZ/VD+GAxB817bB3Iy/Z8Nt3fohHpgVL4kL7iI0lUQnxeuHX+CMMahwbD6ASTbuz
GdZ2KdrzBM13W6B9s0ti+OTbrS/SAti7vVg5YTJ3V0Fa6QjK+0JNW46iC/eqZ7L2XYVcDKWO+kd3
ETq5Piw3d4Euz/L7MdGWBrqLYV2zWhH+TJ8OFnnAtbwX/FMW70A3okryGpkKYeaHX0NbJCp5HHf5
hmpVk1WlsP1MXmAMkMZcoT9JVm1EGtCMWrHsyj1Pm/xN9JMxUQ6q71ac74g+dk7OlH+hm1xr6m/p
WrOaRwyCL65bLvYAfC39hT5ap7y1hQchaH9S7SN4RMXfutKp2PwGT9hAAfLb40tGscavNP3LKwoH
XA2zX+L7yyUqL7/s5v8s2oLe0LO5XkYHErNLIFZ2cZtMMsQjCY+3jbrQFocPA47KYEcgJ4fdyT8a
Xr6DIaCBGLtUTJhLLgPD72T/dAgMPvAo0x2uePcMEyJlt78Afc4HvAZzV6JEQTTo3Fxn5P4YzPcY
Y9t814uWyjd/y4ZYvvnSgo7B3Y/ymspvOtbfZkgCQ1F5pFVBlHYiKdnlYJUgGyYiR4wBUNBc1C6R
v1rskUFPhAuSXI78ArUIlwuXqJXKpLXE9BFdeTJ/AkMcR3IxBmaWXFti5EJlbic9Sg/ABOH/oDYU
tMYyDIxmZdlGzGdTMvi0UzCeOiG+KiWLw4aBO9TTUA2Dzt9F4RjZe+ZA6kCMmkp2/7qSEexaEYEM
Q+rrGRPYAMXK83joFJw/D22o6+9SpQeQRAiVELW9wxwf31fNSeDJkwf4n6YzK8aBj9uXMUbtVyIL
NqKuw+FnNTldSTQqBq3j3H09GGgpaFyWAH953hCMR+yM7YF2u4mI2A4b/Ti7WDLKatpf9Xbx0cKe
hdGqKDytAYbt8vBlgCOyOkM6jhTd+hwysg1eHvbG75lXcHHdfzy4t2PGK7iLoEtU75m8QxMRO2vP
VOGdurN7bnNg7VPOdG1vcCU+KUH5DtGk9I0O6yLJ5RrGmKq3OY7szyiNmzpPI1EmM1tjZd4GcPWi
KPn1sixk3v/EhXmTOfc234U4po2hMMpx3m0iWgoYIHuB7QeK21prkclnsVd5tNBRqzIabupdx695
1eCfqtjWAF0USu4lmDcAq7YSVCjwAIN/EOt60QrElbZHNnhPLJHH68H7tOtiEqC81CLLwmvl5Bx3
jDjYR0nDsC9ypJCh7qeVTAax1ONFf7u4jrM5WdECA/DxV3ZiGW6dyc8x2R5ADZSKXhDOiOgnSmwF
1690EWW+Vf8LKdfcAau0qGW3sFBrr9mDV+Fwdqmf+uzSU1VuzlxwPOdv9kdWx0DBEJmybSyeG3su
lCY+YR/VqSdEcl28oISoUApbv5EtcvQNL0QB53WH5261WxxRyd2c6YM2ze554X9KPLeYYtCQU27i
O4Q5GnidYS67MiATV70dbhRVs2dGiewMk4Ru378/xAOF4jZ2UF2GPE+Nc2V4Ncot9qU9qJgw/DLs
4Y+3kj/+WhGoPeWrB+BU44nhJ/YUUDYwFk+Rx0baMMQVO+Cm5rFz5ZJrcHLFHWazZZ+vbnztSSHl
+j4feSb3pYQZ/l/yrBq6WNzWWrHM2fcI+1EdJ1EexY8/QG0rE62XhoYYD3w457ce8otUX8XJccNP
taUbKBaQFidBGGB3k4bhLk+W6Dk37qMNVJJcwC1B0qY+TnaCigVpXc+gYoOeIXnuNEPeF5VWbBZ0
yysoz03iWUL6k07YexLeUR0yNjfF2ad8QnjQ4/XmpaNuxiP94CbkGT86WqhBTOAcRG5bWXTHVUXn
5O3TMlzL2lAPOcF83YxGQ1IE/3E76zlCphVd3bteE+gIWVMGar3EwH6HmabAi1tKh3v8qeP1dhla
i/1HHPjDCb1QmwigJFYdGbvBeLB9OtSQC+ldIchI3X2XoVseB55PMnA1l519Qq6pPb/LDB4WN8fi
9H3gvDa5GM8PI6+0w46ZXThBECNaZb6UvQDxeWNNkBW798QxnB+ep6z/QEud0RY1npy/y+j7+duB
8dKaW3L3ca9KJayrT5c8M6mcDtYbEeTWORXuONQWbQJykU3WHny/wAuD3jR0wQoDEzuxgU1iH2tC
8CgoDd6hHG1xscbHtqv90UUApbdKJYkBXT3KmL7G/9r42pwjvMhWVlGUYwlectw+hstJOigj2VCq
QYE49Qpl+2r0Pzkyrg62xUbhnx3kfrtMrdKbxp0t1xaKDFk+HjgF66iO1yKk16+iHxXTuGELUDYq
uzMzVIsKsVlxpUDM6Y+GRuUPhEUp97h2+6DEhnfhP967wp7FqMTkUxxVpI+iAB7FNk69jjzjg9ZJ
WO90ZqHauMo85txe87CWZtLJW/di5zTYWkBfpAKf60Rf9fpyvuXphNr8jVvMnCBnnqLg3S4kQl/3
ReOHgvuHJapMXXKJoZCmWK+ZJSdaESOJozJDlg1thZGvSQ6UbiDHHMpYL/PutvIC9f5D1pNWurEp
HO6Jy4J9m8iQD+k/ZFqsW5HG+1lTQdShSMQ0u7YUUrEKLmFMw7iC7uFBxgSuFR0xK809TCmu0zOm
zCvD05nBwqCZTNq+33Q06QLEo7xzaN2Rso31HznjyA+GrPirJa7bkloOEPdXDzvtNqQkOU8p+Qfx
rrzd0snn84ncS+zMluJRQDnqMTCGJG5bAvcF9U6uy+0JbEXSUVUA7tLw1oE/zVKl8sJ3lxx+jMNM
pWQGA5xaeKPtvJQFWiEkUvnNzdSuY+jh051eZktRGoCnPBPvF6KyrOiYH2g06sePDfoQO8wUbgta
eMKQaIQCg2mjR068gO9iQbxBmJ3IOSaJBh8yEbaL9sETE3J9Rh9rv5I6T8ir9GZdZTnnrrE5+1ro
CexI7x8uH9NamHNUAHTr8uwFGc8L9FT961V+qlsYyk4x66XaqZjQNwqgc27Hnj+qwIuEuVwCJiLS
JLVjT3eyr6r7LIjLMI8XETU/dbAcocZ+W6S17nPUQP1R6XPjnxE7dlC9gNjnCnDdxNrCiiBvBIu0
eR6hD6gGTsGhk+ZF5B2uUZ7x4wfjhapXa2VvUkaU/YNs+DzYjQcWBw7HbTKM07qBw5jrr68YVjZC
/GdJdmf1EvZkXZpVehjUH74rc6JQDZ0ThaIXzmuv/lL074tQyM+72Og9S8wfKvRQakWiE8vJZHHO
GgXGxPsibM/os7/Rxvh2iPKCCct+9YoVm6yvQNLjX+0Q9PSfzC30XufeRf6wkh1p87DEha9u6xwG
moi7PXZlHZg5vXxR5BpNMgvslgEbfVFOuFVA4kTdlRKQNcx/ftDH/sKspTfTDMTu4nbIVHd1Ldhs
s9vDVuPa0+K2KkedmO3u5xdGyEmktgNLePCqtzMuEIf+nX8wvhtovJdy7Cry3cRAHIy6o1kI7TY2
jrUrqvmfzBUuHV/m1bEzqhzM28+Kbe859mClovqZrpLlVKKKn26dxL2zTliXK6PiWcNMtyGx/Mf6
oTzV4/yCINzxiselijDp3CiWBoQiPaazPWyqrH0oYk6wKE3V79U6PAvrYEVRhb4V86Abk6dAUupE
/UhsL6FgsMyX6n6tpPsQA97U0rllDVKhxSXd5zZWfR/FFYbwcyU6peOwxx52SZ5cVuARg3SIBTZ5
TFKaqqVi9XrAbOewqeECw+JF+2K3BnMduEZdA7L6TUTfDwuZHFgV7ZRTI7KdLC8XFiEcyamUrSU6
dnFbc69lywQ+giIWElExH+cmHY2PhWVnjP5sOyHuWamrRulbGcK9ugEZLrgJZm50poAqhIjrwIIU
XsL74UHYQiEVXKPpfuo5AtbmmKb1SN52DXzrYgp+sr/Kc2zySsAmT7+yxnrS3OFggVI64VpV13O0
NELGuCiP/PsVOsmw3NiZ9vZtWIfeR/RTWe1u4chNR4sBywk9kCqA1ujSvaXp9avtrV6tWINFz4do
U1Kw2P8Zoz8B8nohe9vGaeYvDaC95/Kro/iKRMQBU1sg+DGBGUOYoqGUHCDXj+6aH9Ub9HmQX2ri
uFT+XddXfHxuHfFJlnd3F4yU8SzFrOJWu1in4NU76etiwowKHhOeq5Iy9iHzybSEuVCMjZMSlmXV
EQfBsWwWmY7AN+OPqragannSEqKL2lqJz9v1aGZBGCdl5FEVKHa9wDwcNrYzYlfKmr0EUObYLtfN
6ALdnhhrlW8q+KNCKRrYnUNhWfe+mNHRvc/Z44NTKk0evJnn3LDIa1JVj4gE5k1Vkz+fgVj/EIHX
njgTRLGQ+JeyAyAd9cxUq1r8g4Ivuwkqk0hIECI6G6GlBBo1b02h0idTo7jwgXqduVOYNzzgUsmj
99kwQ4be9eE0eZERIbrcP1GQBiJuOwlNFnel2Vlw7RQv7QxMY/BBSLodG6/N49BL9g2fm06UY+A3
kJMy7V/B1LNkXdBXzp50514Bx4g+1ZWKlwCcs4Fh7ejdV8QNlIiWlNqmE/59NV8/2uxRHEfwWy5+
YU1zWNLW2p+fdxsIEO2GGX19pEDkMrsEd/KjaX8gC+DcMlF+OpYdr5fTd9c/S3KgQyCRAjGBSXPt
AsQ31WhXA2snuiRjCJKS0tzbG92hxl63wmdBSeXfaL7+5vfwA5vBdbml+DScvlpwH+iQiYiyeEjQ
K22QctIr0cO2dROboE55f3LKFyNJxdQznLh8TZsqhiLETF5G+ZOIjJ2xZEsKOTKJ2Qo6gyDMJNdU
DDpvWn1slhdfWmUZRiMJNs0cmGJX/npzwZmLFgEAzK+fJ3BLcPVhx1cy3ri82FGBIJvjE0nPPCik
7U08ynpl10MPycPcGsnBwpykUovbl/EP/hzNwI2+xbT8sT5g+tGFUBhyCATns2Apvz34QT+ntKSm
OvjtndW9lD0n8BuuiAbRduKJkB4NcQCrDVnlUNiht0/wEajWatjkuG/g69OLtIAirZwZnLxEssc/
6EEMi4jQwQz+qN/M5/b6h4zaTffikLEFgmJ/tkTGogKrzkR74EmK9P42O8HuW0bCf9NMiPqQipcl
QXFxLORgjWQpviUGrGOCHC0kjVh0NgmCi8Pr04Jc3sQcClORPcceA8vLpu6ixlHUAAd9K4qal4i/
bIniHnaVtVlYv3JopB+BMSBoPDE75Nr5noWIoIhUSOSr2I6BXs1dr0BMFD3SR9b1lf+Fs28Gkgzu
z7HsSi2xKmm53hDRhqF/oky3ImbtSzlZENAWmjJ1As5YH/LPn4B/PRr/7fiZbGopLtZ4IG2LvwN4
O7FXDvgvNwlwU30gJsvBLd37E37xOq8ho0VYQKYGXJ/Q82Varo0KTZrlilNegTTRCwV9sNvtzdq5
BlteCByG6R+1P+2CgZtveT+9u4k6fHghw3GHtel7G6OF4+LY0qzft2Y+jhN89r4TXbT4zEiNMecA
TeOL8ijO3mc9gzSr0BZVBeC+bDHKsXfcuValzgkOMtX7b5kuKajFJPUYGO96kkZR/oDLqNXM4C2U
UuYlKKJlmL9A+D+40+TKMHX/Nb3MSD0rwYnO1a91ZBA628Fe9nOe2+5ss9xI9RNNuFZ+vhugnqwe
R/yLCimhWVLtsisreDm2cVRSU/E1IvSpGpSNOfTUTOzLB8m9c6QBMEMlWY1/P/Ta7vwJ+78ydZGQ
hokVO1mnxbi6TiafxfBhtBG30ctkguY1z5nvPIItqkiXnK6M03lqn6jFK4lwVycqdJ7uS+5Xlf0U
AXj1rgYYkwb2ZMnjDWLfiABY7wl2/LG7VBOS4OHrF7fdxZVuB2NzqOBwGj52vroxqPmRCHifc34/
gg1rPP4XNAGG0op3HsE0yX4juPohMQC/4KUmP0KmYRcgWDwefdCQQxqbNBqFnOsgt1rzYgSMC3A7
GaMg1fv4VPnzeNQqDg5WzUCIq/HztQznUUKTqP5igDKkz66dhXFM0E3HRvWQ1HPR2UnD4T6mAnSH
qyZgUHu6/oJucdHipe+kLhiHaI1DkLQ6wU6wdSZQr9jwMrd4jA5X79dffQEBU6QKMN2iE2HNrK/i
Ts99e4m3XjKOKvXmDw1+m8JDofBlbO75iL3hwc52wx7yNCph6DFLcB3EtTgWl0T3lkrsqvjcgSkY
6txhVDRl95wIDu2UYmc4hyQHNlbHdRaGMRct8qOdXhtWmEzu+wEKyaSLl8N3C9Dv+lpj1dZwMTzl
ygUqUYzldzhk4R+wXWTGOwQfHzO8FNEWSZfeNWpgW5vYwz5ePPn9BJ5ZihVXUxKyz0F+Yw9yUrT1
ChnDI+6unAoEtRwRDke5uj18OdvYnARG4jg8hM7xjFMJYNX5S1Xrybm6AoSCUsjlTmJUtY9SuKzQ
yDsMU2ANnjpCKnOgmJRhfH/oiABrwQCIiasWBS+izrD72KikvpCEX2r7UXi8buDpxfFheW6qGOqH
YtwO+QTRncTTLGUh+kaV+rZmzGhBy1I6Q6H/3r/3jH0XNcJ5+NIGSQOISRBP39sY5MPhImzCmfiF
TQ2AZf5slWmAmiPIZx3L4Pv641GfdC0VE3ipW35XUB+P/djRa8O9flPg3SSClFhMC10RTD+Pozhp
8aTTht8t6vRBqa5NqVKH2rhz9tel8bn0uYwM3pC2JbN8BNgJHtXmUyyLxrhkaYECxNmM64A+STLA
olKyv9aSsvq4+Fm0wF/37T/q/fq2G4ahPaSlPtlaxqw8MQ7m7kA1+FyMsv8NsQL+NiS1i1b1ZJXJ
1hSWuOxJfNdgNaezWpfRNiJlAOD8PnxGppR8v/r5KoM0KyALQgcTl7NXIqFJkITMPZyhiuY6aUj7
8SGkEKo6SWTJVPqaE7pI0lve7nEArB1c+FzUvz7TRQgWng0PS95LEd0T4TXfpaDWf4XmrwreKdeU
pOe1qvELGDaadrtq0Jgp97emWUtnwevAYyqt46Fu51uXxT0tXtdu44cC4sjCZk2udPsT7sG0fmSQ
nrSDxkkPHg==
`protect end_protected

