

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KXJ+KQFrskV+mMOtKobUOdwBU1Q96L1VjuICu4OyHPs6SXeHG6wnV80Fbxov/EzzO8x0Z3emKj2l
1HeobMZFAQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X4MwXfUrUSWPkQbt5itoHIH8a6wAv/G8Rj+yp8qV7SeDqQStFUllazNjiSTqZslwsd31+6cYFL96
6zDC/D+OYJSVLVhGm8PIy5CAObI6vrQTlPLpCyfSAtnhsAtbpB+/xlglwIui9BMVFAHugGmjRC+C
iEY17T6TvdLguPq7/2w=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AY6GI+RVO46tZSokl+Im9Qjzoj9Y0Yy5iXxh6iX/9ufj7UK+y/Fu/+jqZGCXnL/D3x5Vw9DvYinN
OZISR+sb1tSrIdKCMSqiOBiGlkfXJX4yx+M3XhT1daec0H95htsSln8Yy5K1heMbTBqwINepRZ7U
JrYhJ3Q2JY1ank6jhbTfC/3R00Z4shzx6DiyAkPWDlGj2jAP7UB2UON4rM5Epg2pIBwbbWQAAHTT
liAIssHV0g/Th4AG8Bf4fCEvKsyZbGuanw6XpNnQFIByrnhyynf/4UpMhc/cwEDSo/e/VIetTjiO
8GPRl0paJ2NqqL3iKfepGqCngXHn6d7TC8EvTg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eQCEBXw9ntq2jHoQJtOMWv98AZN5oshrWog2KHmvb0lnK4113pxvwRuEJXr3iDkegHdv+cJXTbmV
8KSCmD8ChKWkFXee/YjyBeJMc10QmohX4Df+J9wImo1z5bbKXBwKiQUjlqkYleMDscVyreupEO0R
OTEbw2wpFMA98KnrxKGJw/X3jY2Nad/7JCJB0vTE/g97Kv5eJ7mB6QLrkoTW8eE1mxiIT95uwU9/
Y+V0S+/QTWiV/Wy+tbO/lKYDetTh+81EC5aPb1AS8kQr5jmAhi++8HBlocjmTsLpnBT3l8E5jdrY
fTh3V2oMq60AdOU1465MpStQpJeOcnyhacy5fQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iq8QZZRvFbiL1D4/Ut/JYE+zjq0864+0wF2SilIWU8VHt5TtRRWIagETipUl8rN2FoyGyUg5scS6
d8nSqHAHLTg38L4QzRQEvkmHZ402zq1AywpH+KMXRCEpOzPVOSxNEW1EfktEXBy7EkC7JSpUZ+Db
s6JHsLkDPJ23VSMVSBo1gc4uOdYpop1ncZh6UN3ojGOenKLJibChBpSW9wy0ARqgedKvd5kHn9qK
QXAuDWmqT6HAXiRLvFbXFOQ+xZuyNr+SpToYRvXR1xGUXnXGMCWcv3DlIhK+tL3TnGKh9xBMt+SQ
XbY8H5PqD6F036BBQ+C3yL16yhDmA2o9cdOYLw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OEkw400+LKMrls4nTgbVTZ3P1EKeX5UpOnw+zEzf/LSzF3fV/voU/boIwWGplHAsHALpt4XBOVfd
t+PwzEfEgmsMqapviTLAi1nHqL0rSZoU/TtoxUvPAdVscAAzxs+QHMxHRAQXklxyhzBIyB6exb7q
otSeZ8tJ3vVmgyJfRFg=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hjbrFSOsnBewHCQJmsQwWPLXEBgWWlMnbjbcjBor8jiUxGJ5aN5yhGN+Z91PBg3J9NjiPcN/OqZv
1nBcMWRDZRUaV7niwSRKBFH5EU4hSshIo8qhSEXZ8Enh2wk8ZwP7nkVBjpQqshjBMRp47ZvVeqSS
/Qpv+YGPB90Y45prWsH2cdu0en3QY1q75Hfy3/hSS1ueBggYNIzz5qVQ9qc/N503Sl0qpujT+f30
nPcb9BV9jXIJ1ly6R4vCvu8D0cRs+hv3UTN+gGWv8t+bTGV0ztqMojNvBqHUTIm3rXfaBrqTfVAf
A+9yth4NgrpbJBjDH9nw6zqU9a35TRnhmJTLKQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74240)
`protect data_block
cvFCmWxWK98V0pkmjx8eZ3wnPYlJK9/ZdGeX+K2C/3gv7itF01w1D78A1LXf1Fmno7puAqHYbWCd
RAEdRhQgNScMbuNxWDfOHL8ATp2NOZ4GwmvEescK6sMaxKfHt8yjjCmb1pBDBvyM/YsZqANNlahy
d7Mq31ujkm8JqEsYKJ34rjhTkIUC9ZfWzNdy4YX6vJdXJp0IJMEdgJRYdhHKhHqzW8gWuky+uveP
acXD1iCxBrUUkye1a+wHos7f7FBqq4QeCJs+64eNsG2SG48iX+aRuhzB/EL6ZYdFvqxDT+ceOc+9
A2yPoBhxzfauwhqsUUS3VAr2yMA9ecitR6v9zyMPXGJBomZwYqkr4awMPss4vWDu/rMw4JXvWpS3
9hDRI4INzcQZlT2l2hF24Gy4C1I7Im10tDZ2t2tmyl54cEF3p5SwApfmKFgKS/6tRFMt6T9lsczV
j6DMhQVB0WLUvOizrVJDaFgd4Q9pwZoRHcE5XHh8b5xpo3BgllyPWED9sYaypsOH2FDlWE3NOOFU
N6KWJQAPzEodC6QP8YfplLOY/uOT5UIZ39IXyhYnnqDte8fCkdLK3U8S7YxJ5PiVFNjudF7Zvtyo
VyfQ12BZb8PE+Ojefh3FRw1AtO0Sec3exO8/wPqNwrOWzLFaJvB1607kO3yMYTXeP4JdGyK9ax//
xcMlYMFycTpnlBxxidBSd8OR94Hm4aDxzInCbpdUZRzbrWqVek7AAbgcGxUH67ImaOhJrDiKpDI/
BhAuxogR5JwUxgCPCAODg1ToI4QqMPTYy3rti5FoWd1yZEq7FelutWV1cg7qoMCVhfIQjyXSR0Sb
VpzuEsKyrWXZfaedNwrSiu8W8f5+9kRCYiwlMwPZCNARsBWVevnqYbpnDoSR0+b5Y+hY6DolIEO3
1IjcBrZRB4HMYi+Z9ExK2tjnv7Cfr+1l2+kvjLQgNwi9TTNDKTjWreyc9a9Wm/vRWwCsRiWcJ337
ftJVwNpf9Qw4reUSunEv0vE6j1yKNp6wpgPINT12nE8lYzwNkNHr5+9NGsnGKmc8Fcvjs3E4rDny
JB0rzWJFN1R8+AYjR2m3wosZIdRzqvYVeABw90uNoeqpEQXcX6hnAGo/jC2REPsnwuRcV+vAl90j
DU7rgcFJ0x+O7ja3Aw2pbmzh7WR/e1KAviZBayex33PVsIE0IqkysRT77bv+ViBmkFYoV3INDWa1
OrwBNNazqvSumwiRei0FQJRS+CWOljwk2hmWIYYz3kkBsE0xhjGjxvPbzSEYVwbq/A5u8k9rTcJa
JBdtCO8yhUe9s68bgJq76nGv+LSoCmfrEgymHOsVSJpiJdFbbFWOnrTVvniIO48BN/Z+PTwoXJOu
tMSSbBGykNhh8ZpuMbzyocIsqt2jw96JJmXIu/xf7Ch8jhHzRujPQMKzEnfvOSHV1ggKZzvLKQzO
pT7/Y/adZr8ewuAwi22diUD62PEH8ZdgRr9K3NjhMKc6BZ7hh7hurbJYuD6v31dOYVK6Fyp5rZDC
krhIDk2veqMGmFqCeak3+H7/8y1MoWM8NuEdUO6lXbxF3N2KcPIQvV3/NZZNUVp4kx4TTBnyGlVv
GU8J1v/ab4kdN52f4qYkX0VazlQoL03E/IeHNU8tpcedzlYQCPmD0cTQBZ2NlTNqWXXNmnXOnIlW
o9gbw57iXJdz+EQn1C9vuttVnnVjjS8mRssNfAxjBWQ+g8sYijmAwNTlk/kKYZbi4EZWwN2Gcb5d
JbpNkYD5VkGETaBFsyWVTFchL/NhcaXubL8WIqekSGlSC7gZx8SZ4KXvRMkdoqJ3IvEreRbk7Xfc
JgE+bsMJXnIUQeoxcz8XfI8N0IC0akB0VEw7pdI51VwUHQ51xjyrmf0EEvgKyX3HJq5CuXLPCyo0
y/u2NHv98KFIGFiGTjTx/va+PPCCPDZ5baVRBnMkjNq3/lE/4SpoxKl1SkAQiQjD3vBonuZdIt2G
19IOH5GLPRTNOfQfCsR+EhfIpBiZwBXOwXFWLdkZ2NUxTgyKl0FCZnuBccOSa9CtOrmEVkbWBHvf
OoRH0vxOyyswdl+4sstA9Mf9eQqiVCQsitDxYK32GhojyKqh9EjSCKNaHbd54pLnnyb51+QPDsPr
gArL+HlK3mYEQCaJ5eLVfsqCzrwVJLs3aJO0fPvyaTC3xZMOpqwhr1HvhAoh5+KS5byiML3GYpRw
EpjrieZWbrka+c8u+omMYyZ852LGzl69VC2yK3NPPyKwYeYNbClgI3P6Yssz2k7pL25hzneOSeCM
6clMvGWncFfIAn3AecmVD8tx13LQ0GdoNPzEwkqvNkx4kzaYI7aTkKFmEB/CS8h/1T3SVbQZOf9d
956vcOhKHZbXi9hEyHzlYvIJlH7Pm2kHoLEnR+PwRAmi4XBWPU1dfCV2ja2ZMtq+5uLjzsWaTE3d
ojcHaGoqH2AFpHARb3ZAmI/84mI11Lu1o7POSX8tVJYT50EApLTBzo9l8h9DknXBjELsRvHkVORO
JipiS4oamsTVqlc06nmijCNsa3cXAkVgPiUUZzwRQISo+ADnTYERczs609SdVW/uyhsIh8jd1RiT
paVjNo4pkBczScbx70EYyHFh6m+SCzj+26LWUOaU2+F9eSNW9OKI9MMVfo9lgkiHg3X4q50lig7G
bzpMwNdgiB+BYdmV5jSdNjSyPu7UE0QBX9gq4rvmZklXGcoIDAcCLPSbAO1pbNAtDUZFKT7gC+1q
Q13QEOkpAJDG7YrCWPnkBNflS5M8aga5Lh/kbAS3xuYSA+whSCvbGkwNTr9YV0OosWzcahTOTX/a
vO5FYWFGDvnpbimCQUxq6AHaVacSaY65PLoHYwlT1aRe0eiX0P0WQhI5Hq+iZL4nxn807/2kAWnn
qrCEb7l10GWTvajeIZ0GXHUNOVbPaXO43uaZI2rXUvvT6d0WjJpyo3B3akFdWWWZ7GfQqTavByuj
cEfA/G+ufiiM1cndvqkfQyA9O9RBMgh873gqCgxokcG69RHnIsc8B5+INGakqkqISxh2SlNX/7GL
Y8u2Cp/WDg86nVnQPTKoKj8BvaPcb8J1iDtyLvmqkTGPBe79DqaP9L7MDdbQr22ZSNriDEXRaqS5
DeQkg0RTg4tIZK5tzpui9snWUOMV0jLXJck7VPJp8CO0RjC2ZiIbMKpZWvqr0XyzvC9r3ZRTXvwd
p7CquKnN78UawUWxhjq5VBO84cPhijZP9fzk8nDZios6Poa6toWPe2UmSBXFuzRt78t+IMBTR5i1
36hE3RBHzxxJ4kM69KV9RLuHW3ssp9zVWk/R6xeVAeKtKBPYChXUUH4An9e5DjmACNe44PZ0np6a
OMLRGBlWVMeUE4/Va0B4vISUE8LgjEj2enTNrzX2g4oklV81SdObCVBCCzDYlz5b10K4e4hOv+eX
HTQBES9ZtWlK+paf2kZ6WVvtn2YTqg2/rxXO/+/hqNyfeOmdLyPgYFNC0KZJfflGFk9y5EdG46e9
HL5qQlGFV2pAp3M7aFei5/xHUYL5695ARsb0qqEqgn3qPBuIZyb71pWjtBDKrODBpUsbu1C7ztcy
B6dxkg2wsUkVBZ85A1hCihKO7gKYoZQqpIHajVTAc4CRhtuCcD63Qv+FqP1tVrZa/SyrQwT9F4wu
TnfJoxmY3g+ccWKc2R/v0SfEXOF3pL2iRbUoIeRxLzyK06AtDsH8MT3cYYqpCU5JWRkWkMItY7jp
QufnTRyb8pDqSnBvt0Co7qnzrSPFcrtKM/URYYAr/xwrs1PRlqKUkBu789NfwdhhGVbEeNTC9a+Y
f5sCPqioyZHOOpKnVn6dNIVdGd3Qei69xd2yOa9os8wznJMk3bYbp99pI8x6QABYT85stYM1wDsZ
tXhQwz22DcNZLBKl4jqS3sWsN6JtjhXIczUYgpYj219dECiX/gHuTmWKf8T97wfsT1pUxSkwEAoK
hO1RfC8KW0uC7HRvm/TzvBREgKIaKEvyKa5K55o8ExNs68WbNMctdNa3FFd8kxI3w4VRcRWrVhXW
DCR50QsuFtM+8bl97Ix0M8jSq2OgDGlxDBjzm7vJoqtzOipNsqMGZhexOiypIdQZwK7Pfw7bPf+M
6NDtqwRargl5Epf6U2Vd4TrTL5TlXMN843DSorXS+0POAJ+pxAxYj9VzP6yy79+FH777W8jVzFFx
/84STxkQ66dSvvbbGyiLmHb9RbC4/icK37nlmVVICTT03D5Ved0moAWx12StFtcLD+705QBv7PbW
8LqbG3RRjnXgZKOr80BHleNIq8gPivJDeegse4jIA3pEfXbdiwfeWer40okWb3CzjS9VZnc7Th8I
ens7oEjJGBH4JwUswBtToKg/+rjVCOMkthLACD1nmVAGrfaA+cCH93BhA+DVf5oZ6T0dj7aVWSR2
/7kQlg+VKyzi+zELeS+cNDZ2lKyar7wtz/gpOgiU/hLWO7OYsxDBah9CiLr4pTH3d7vbI5rgzyu6
2EZaT7oHQ0xJFrJmoq3RJFNa5dEORKht3pJ/WrzIl7gFRBtvldScEj00zhjtnvW8Hc5eb8nIih0e
GdFWbTYQqTBDVcBLs9nyGDcXY7IMXBxHB9F4MZpWhi5xW2v84OWBFjTnipHYKoWz2pyTH+0aTqw8
Gok60ElhKuwtxqxSChsjQIdJIzXfrljeGePIE8NvVPxUjsw1dFuAQi615m1wRPcKksk+Bmma4qaa
DOdC9VZLKgOfS3WJHSDDvWm3sFHoedW4brE8FLbUWX3Hgi9XGHU0mzK2gFk0fBxYcy6+zALuDi6B
88fsdlvQ7Nil5T5gl/0H9IuVuQGsUfQ8OGNXxSjqlvK34MNfPQC5YIDLjdiYjpDUwU1XPAJjIh/R
YajugvVSe5+PDkRKoIUO6u5SoOezs/iZ11nV2AtG+wOFYK6RPBbStUIQ0fsOwcOalf8eMOLCZAou
4GEgphjz9jXOJsrfWNXLn9ZVLQ2PqaeFvQyouHaVFlHE5tasNUlccQYUiRZYc6Jjy8mD28znqyx/
bXt2gJXiDoSldaF+VSZPOA+KMTQc7rZU7/X14tz7PpdadQq6o8UAtGh15Keeu967hcWM/k8cpp/t
VpTXKvene+S0IwwTjn7Q72DsdjMNM2fuQlw16KpA1tuTGop6EhH13ws9BWj1VpGqLNHNQmmZCWzN
dsrY3ETvWHQRuzdB8ptoMerucGrG59U52gmqiTAEvW4TBL42bBqOmSpsHbu+J3GG6JakeS/gNBdf
+AZtb7AAeXSNYqe8afjQQvqnr2ez+7yQU+BfAdrDuWgScGQ5oR5brx2LLWhNOVL80fFjSozzEj8W
G6DP3lvgkGvHqAHIAmfMebGD92vN61AKnHYh3EHCCdrzxhpB2obf0BD5ECB/UQACPuZ5f7xbWHMe
KbjEhmGKz7JbRJgiGIeTqrAgZu8hBZkaanaQemGgZOcQfDW52+X6eD+wcUag7+9U0Z5MOqyJrEYl
4+9uJADSm86AhH+vbKFIPpykVSzO8dEYkCDFH8kAe2YEdne94hNfaNzge9oHPyG0VIug81vO9v8n
xQwBXef8XqVN9I40K/7BgK9Kb6EkZniEoMMoMw+4LYZHMu8G7trN5LMt9KY05PYLIDUPremsDIN9
JtyYtL0hb3aSlYlpoonVOg76lVTLGktHy/WEQSavoqcOcjx91vAWILJy5kMo50pFUiVu5jmBGiVL
mUtH/6Me+h7IpQ6T72UVB+nRI/0hw7e8XW7kpVKdJOPWUGt5SlYxrf5DqKwgHj9EbihERAu0+CPp
nZRBHXuoJ3lrc+mzaB1yZzf3+nF3R7tmqlCwa0+Cq5N0LctB6zG91wpnULOrP5C4DxRpUD16+J+M
W7CGDocnrWN7MbDcayNeds189skljxtrRWlIUAl/krhAytI7FrzBP6j4l20Ln+MvP8RjWuKgWOaP
4x0jFzHEl11KNmE/WDbo3bjykq1L/vrNoyf1+SFds4k+UYoLQ9Xcgmr7x52XmRDfSaJsYn9lq/Jj
q65AdiG/YgPi+wMtnUB5dCVhEOdUtjGleU75wjYMiFux92vTkfOJpcfO/PedTpQnLS+7+uDJuwFm
7T4qcsRA/VDMFBm/S1jRzV6GKqK0lSdUnvt6IFuVqLVr1iVRjrHoI4huwxqclzv5JwcQabXlX5or
lkb4vF6xY9CnzKf/7LtsDPKd/Xw4PZ9ySRInyZ0MdyYHgTUzTtU4xSvSnNcQIvxgRsFaWUu2KVpe
EmYKfM4ZQoGONZnau4SI28bU2tspwh1wl8EIQT/jwKEMcRNxM3w3cFM8B7U5TlNZefUdbKN/tpiU
0GxD8Dk4UNgBjH0tgKz7j/ZTe2mvTQ+vBwLEexZkVa+x8c3BDl1EiZMYXsssgBZ7zQpTqfG1QqkF
OFmYSC2Cv40NLICSB4kCwXigRUuqdjs65uuEhGq9b3NjNrr7PM0eNCkc5TwdWM344E9nfm0gB67W
d5EhVEZ7RJAImEwFjXs+b0wE66aTJBgJrRCNGl/BLTeWwp//so6aj0LMf6OiGpuLW6Gst/fcFXJE
n9tCCzmDddzRvLt40P1v0m+eEGO3zhKq/ULWqQ8og0Pbpt0TonDDBjQrTaKELScNAkOZJ9At1K7Q
WOIfSU51k5SDtBsMd/2/+Ih9M9zncd6ucahYPtLOyjahqV0wJffq3n7tbhNkqw0snFhYp/QrCptg
DmJWfZ3eN8Z6V8oTsqNneh4RqEgaakWJpjDVwXqcl/B8t6R5cH+nQ9O1SLnnSrg40aZ6hy0oVBiy
dKAIfPdB3PZfS/++PaKzTkOiN0tB+zh8B6JAv2unajfn1HTheRSvTqUwfKbUhoJpfNWZZqVJLdUC
4ngBVg1zKoVdq+n/w88EWSWDJ12tuRyq1nPaqp1xQpfwTxpyPokU2A24pkFKLKCLzFdR9sPuPrNx
qIV019dV+jzmk8A+L+3ARcpODXfP+35DhG4zI9psc6nPBgqqgsK0HXfR6q+Cmf+cp2raHtNfgU9g
E2sXr59fR52l5qtO2ang1bkQVmPEqHeyjiRgh7p+1NnY5RD82ZpXoxLj1gfDwyVy2Yj91dvvwfgA
86NYN4zJsJJBZGWoOSBez44Oe2t10OzAlEkfbAKIU+M8NAkIK++M8rWXtJyxNSM288QpIOEJP9v6
0ZpEYpJgtbxmdOpyoXTVKfj4oGztliQPFjOUTaiFKCICggGowK6zMEKZC0/tf3m5szpsxt/GnlKO
tDX/0WkPYa7rf/Ayde+D3D7NDY4Q+BGDgFyCptU7ciWNQMvh5TbIhieNxSfqfYGpCjVULjzJrctQ
jRGVkmZ/yGGkoCciZXz5hYMJtHAVD/KAm4yI2Ul1PyGiIwmshD46VUl9zGOLnNtLrzOqUgYCSTDA
ige5v491kp7SzKWQdED0GtaN5NhUGQni1RbV7/r1qUjww7z71mUYetQkjy42q8BnBdFk32q4bSEr
A4D6XtB/KDJJ5IMFvM4FNamTN0TFLP487eWJFobxmpizxTUD1XqJZspN5I9ffRdAEW/g/C6Y2OFO
W5luVOx3SV6OpHX1FlSWByC1sJ1i3gg9pbYiiZLUmGXTc3UgSu2wAqaG4795olnX8J9eFdLTWG1q
6VOxA55cola1HZ/8gm4cILVCgLy9MaotzjqjSf3Yvojs940v1SdHkujzTZ1kTgLCrctbFXbUvDou
EWjClMuX3CUsuBXxUVnQPAEDmBArnSMSz5vqPlB/buR7Z/QBgOLdJ2sDvld+fJlEj/k4n0W4NGgf
BsDDnnC0PAQkPaAL6npAsr63dBzyTV+W5+S/KCq3rcJtSp4zwrenu7/mLs0RzYJptAw/bVe/5eUu
/co017fZa+4ZUJ0EKDHQBDPhxHd5DPBgZ0C1/a0U6cIeke2ieUGa+rDewyl0AqWT1osPo3++uK0J
BOINf4Gj+f/SRTm7GQLESQP0b+QlihZx5HW8n4+D26AOjHilfDWhSWsiXV57F6h0bxMYytIlMDYM
hYGyEaNhfA0zklHjukgmR39m0UysOWHKZnNcP7NBUDeh17mXLw0Wz9aHKPYdJhvmc9FyesucvnT4
O0RA9PNHR29bNSAXx1IuyAIYgVAxfroMGA/PWsewJ8qzx6r4p7coJQHAV+JmhBDRy7G8kke5Pt8s
W+mM8aFGPZ4BlQ8t8MmvmYO8Pv/oNd9XcLMRMzXy/kVQ6O/KLvw6HJcx+d+ID079297qw4F9fHJt
Y0iO/aa9fwpVVVtE3yFzrDoEMusXSEdEI6WZx5MEU21lbI6jeTW4Ae4eBQuRt1jNxl88K7sJ0Ai9
yZIVkUltya2dU+B3KdCsJfQA6CbpRZywa5x1+GqZ/03dapLy/ZZ9ncOZpbgnyo6RSwmEz0CSk/IS
X/LllvNFW3VwVZoIO7PwLNlZYfHTMXk1c7uxIGPna9YhtpcWvQlDAYMqxCdvjqHgGrJoKccmiHoq
55Ojn4bQnad90KlytKbnEP7+Kx9hWzjosDibn4KqSIFG638UuPXu7k3jfDlWI383kChjuz4oV2+r
uAg10xhJI7VkFpfqsK4x8RHCqvyHABVqvQDLrTTemvrSVZH3wksBh1pWdI1HDaFrqIeUXSBbx5QV
QM8+qWgjunTGjZ/o7zaT8e1d4mvbS/ymwGGj1rfrQ5FZCeCpjNO8xiAIhWF2yYP12ulY/0V3OfCR
HdHB64INVz94DLsfpHZVsov81y3oj0ap5rFEZYqXkyOm6qB5JBx/3QN6tKIe41Y5ahU7sqpxc3uH
faJiXyY0HYG5rJqnP4O5ZZtcXXGfuqSxRbm+lbjytpKpKD2ic6UpCHp7xFLqKiz9suvyGPcBD+/6
2wjyjGSgC7+XsdWOnaaX8BjmH8tDV2LJF/8+Nqd4P4hedTqDoh9T+82fjnhhSaozIjfOA63cGf9Z
zA8PQuqF4ttlxFLRDG9lm4V0/TDXfkvziMDh3711NNGsRU95c1vfrIPyDqoo7s+vkJmp8b9qF1d3
DDmvyS/2P9dEM1PeiC3DPIyAR83TJ5EJwV5o5kxpxY2fQcHlKz64/IbwNWjAKkbFkAvZDAZaFC2h
auogKLZSids5R38+ZrY/5YQ/iNWDe2hBhqdPzbucjVGYdkoVJjOyr6BujF6ldMbYQSDNdAU4awCd
jOF7t1BV+8Za7hypPlUwN/MNTBaJDE0Yme/WtMtm6tjRZ0DllUD2Rb/vhB10fGQyoO7AdpipwDeJ
7rRt3FBVs9A708dMHtY6sMbzGO70A0iJTxT0/Mqlee88Cs4gcmNE2o8a9yDhT0eEBu9tb/0PcVcJ
PXwYRL+7wAetWwNIm6LfT9BJoDzDZ50zrdErdja9rpNTfu6lmL4JZSzJ9SQURzbFbbgWNP4k39Tu
mfSAoAASxbrTFq/cas0OVUKUufdLB4qI+4P1hnVTYRJR7P3dZKxoJpKbSJC3uW55cGvJ7h2+PLW3
KcoVVeng1QWjeWyowzfkb2TSFEG1lW2NT0VIvsqvlK6hBPnVu77zEvjHXkctyablPs0c9vWpkaap
V6Rg0ds6NB+joQkez2sC5SvbKrEFtVvp4MY0xmLTT71SNsuaKXapzA1mTcwCDmYMxUG4Qh2Max3D
BrGwNgbDZxAa/pK2E++SfjJVw1VcorcnmqGcTWZ7OkLhnDPm+NYdd//xEkig8AaA/VoqluKgUVty
8p2COkgWbwNNKf/F9sv0A8lOTTLaFOBx07PyrV41/OT/7JAi8FHbocWT58koYDQTv6CANmQqH95s
qjqPXSGmWbxxzhmxJUBlB2U/CPZMPkwPlkCnnocxoaBhTV5pJCuVhaL5RLf6DEZu6c/ioPmFv06R
SrYgTQsURabsjtCxxbfhaTzwfHdGHjCMAL0Ta2y6oAuimJnSCAoDHJggXEe9taJsMqsVh+7Bk375
5QDPUxO7ept6decrhBxuHmXeD8V/fk5ofWFai9HaMkogihfbuFXPy2+LCFZ1M/kORfyRwhadgOk7
1qetXfsHM4nkTzRg7a6Ee+8P21CvPtud7adjbjZt/coxQmDAIYxIXdJOY35b09QaDd0RVgJZ+Ll/
mpdKZUadOZxU8dLFCrRYsHwe+nskZ4/be5dhBcZzF5Dwyrylprd2CZl/HrAMLclNJ9YtUz42R8bc
q5F80AiFNVESXrL+fX0CA7YSutAr8ZtW79bwnYDNadyJHj8eXkIgs7tqqBBU6Lnr3to9OJ01ci0U
PAXiIRvuC09exahtdo7iG88MMigUQxcQGrSWUGwEYiQf8JX8vAL3+OLNKGUfw1kTsNeeHLSki2P+
2gVY62BrmaVf1RIAcCa61n2BwkDzk1ZgBqEBkOMV5pCYYUoLAYlj+1EZn/QaJDenQP65agSknM9k
fNH0BwZK0/Q/WvF8By99FZmx2eMdeUD0P5Ml4VWfiuI/VnczJoRjq1f6Cjzht5XsqOPI3Bn3LsRH
ahN3CX5+6iA/nft5ulxzdH8/nHGRnG9/evvomPU9Irxcq7uII3xTQkp/uSHMWgKCRCTeAitmQ6GX
p2LNU5CBOnrwgHma6uLJfOBqfgb7drLlVK1VKng5eF+G1QcSPgV0QT+oa6Nrt7zWZtBuckSz7ZxP
zjvK2cB+X4OI2ZgJCsgtlucHmpLuAffRbLHY3oCx1MVPYc61rt7nZD+5sg7cbngR1zPjoXITwOSa
aIcmVDbZcoDhV4p3K/+WPqe4te198bcO+NgVJFtjdRViHGvALDjbf7bibozoF+spLD9l+ebQRfaP
4SgzdYYQBdnjdm+folTe9dpGnSJWSMlGVgBndsnqQbjMIppNVryzfXtR1LFynJAUyJ2EKnOZTjc8
qse9jEhDwSgzeH3Ih3u9l+rvvLnixyOGuigA5gIaURfKd+UNzxSGx+7bj/EAALMAGkuIz0/ofA8E
ZJQh7zMBvtdHEuIvNh86v/X01xW2AhG42U0CyY4qE/H4dhsO2f9nxz3yGcie0HlqAmJzlWSfrdJI
n9VoYBM7F85vlJ6cicQ/kAVLmeTGPu2PRf5gcx2ujqmmvcHr3YD1v76hqSfw096VMYue/XIaARcl
f4DxhaTD4BxsQeTEmp430WKJUhj1Th6j4/y8Vs/UHhNYfZ79XzKnUbU9m3Mo9TIJrkstxfyVsLGB
JglWWEQjijiCAj4YmLrLdptQ45fNZlXJVZyISOglfg3z58eALecI4p+EtiN06Qjy1k2O3yDunU+s
V9aoazhNAMrsiP2UaNiVXZ8iUfP9LuIwDOY8jEr5/Z0zauuuQkncgJGYywZ4ga+gQ68yW8mX0OW9
1CDh5jQqhoUTQoqUt57yddT2THfYnLSHovDxjhzQS6tf0FzjYOT8WaqaJ21oEW560l9K72EB19M8
BxTkIoVz2fd4AaFNTXMEl1cqBYWIRwufc3G5ka79HEkRSibaMJB7O26Jl+DkwIemvW3ZFPHZEPHl
9Tbk7uK4kCBhFYsi3WEynfOomxQKcgQF1JZAwLNNly1gZJIFKSM1mrjJX8gijgm0YiW+zuUTQdP8
uyocR6oLVt5OLQeGrCbZ0JT+v18DdnuE0LJkBZj+w8iII7a2FgSpD4iiPb0fZWhNreamwABwg4lD
g3NFn0O16h1Tmvaw5DebAYKowM0oCTvV1bq5GBD/75c4umYNh+wVC9GzWWOQMVWWcPZmlnmEE+zx
6F9CB+XPMmK3V1BoFg89L/JR7xcSNyUu7Ywa/1OQ7QeE+1dYQEvfHsZtUXM1ECdtIGLOk4m2EJKd
wDy+q2YHesJTIVuuwv9rquViNLdfBTremKjq/PMFVNAq69NVFe57F9PN/1zbduKT8FpVSUdZXH25
28+TK8nWKtT55Knbme/Ua+Jtdk5bvymRfUaP5mnfP6dfD31l6WiFnPYQH7kt2K6tsj+fuy7ipQ2g
SdS5qcCiPL76itajoG5O0ym89zWZMa2Iisb9dUcyHGDb1sS6XGEbqmQWZ3ZgYYH7iugXD5+vodAH
tKZWUGwybgMS3DEIyuBg2fkjTcZDjYYI4ewHz7S4+OlISdmm8qBLxwBJgZ5SFb29lyQV0esNabo7
rYDrdcnUSUmMt80yP1DZCx4PGkWFzV+2Oi8noJpmMXuntesWXv1S5OUBWem+q0yVumuephgRJHkk
6ywYhDe9jklILyHYsgQTeZjcWjOFp3CJeKXTdjQF6fS9rMiPEJ3JZOCyat4ussVKKaaSi9l4xkru
GXhOZFKAMm5ot6nqhsWNwhORSsy3EVgShj3YdgCdkKsMKSeujQ/NAhrjMekcKGsizILrVZdcunEq
g6Q2H6ZFPwAebSskjw/qa3fsqXz9YzAJAW296P1uInpyGBF09kJfYbDP6CWQ54uj7Xo60EdfuWsK
BvHkX1/n3JXmgjkTJ1JipjPAAV0//1JNTjNSO3zyqsp3NfV5znIHngRAxtCHo8KhW0vYqDCwMIHr
tZbIzNTT0pKPyOKEAb3NwcLT6AaKRVB+hdzS9VFVDxxkTyH41HDESE8DPHeqNzbNgin6BpU0sMhT
kubEfsDznoSd1WVtzyueJt9xlaIJf1kB82Be5RyPbTvYWDBEgcOy/IXg8F0g/X+D/bfNxu+wVH9L
SHiw81l+iU6THfH1jamkl47wni7M2hmKNV2Ral3/IQ7uoRQeeTgmGIIAYXj8+/JV7ViIATO3YgEo
NgDY3qWZ2ZEsCFDF4NrTbKi3ahPo/7VgvG6sDPW264F0NPdsTZGeHC2xmmtcE/gM7bHsGwUxPmbc
ZR456+Kmf1qOgdXFPB6RBROucMeSAbUDqZIi9Hu1Je69cg7JvPG+Ytc0SxVpGNfH78mM9l+b5Ai+
oxAj95HqBrL8+wd86TtyM4N/HmYb/LKI/BnU/6dtcvVdg1aTs77ykYk6gRltkgAnOnAy30jLSXgS
5ZwAw5XMnO0rBXfW3gIx0kyEGbXhfSecN3eDCeB2+JSOGulhO/6Oz0ouhqeKBE7U3iZL5mjhGNTS
qXz7HttJqJz0n1TSJ8EJD15aZ2wEmnRiL2/Uq7kXHfCdy0l38ik6VFlkDwzUXs0yFNMfVnJ8gbe2
TUKe7kf8Gqxdd+O9MatMkjOqNkBy48zFuM2ofz/7iIwOEL4GfNVdksla3MJtXj0ME5wmeulIF+g0
wkjNLpoAoWwfk9mJzU/gv8FzkXj9Tg/39Y8vwAMbWm84AhDtcfe2tKm5XCrtz9VhaeAPVUHiigF6
XfX4DQIVu4aIr4Br4Z/Q77r7VPLPxNUoTCW0dwRLfV4yu7nXI2LxX8blRavDePeISBKzLABmzUK5
hlhyt3b/N1q1wVlFNfWvtk2GoTHI9KhRQbk5Rkv6HJyNibd+QUkcX2Uctf5hfrN+/AH0F5VhzLpE
2eAt5mU/0iGyCK/SvCOaFjIO8OzrdZ/um99AOaQUO57hb5eJqQN6g+Uv1vIQxbNA6JT8VyXWnwVH
6qa51wn9Z71OD+H/LBv9Vv8OfzCWuEWL8aANm4vB3LlMolay0pzTcZN7QltWYPdhxQULZQJqQsy+
0ZyW5ejZrrNxcdKhvjHDZ9DcI3hiPvZXFrHf9JhL+imevSBhxnqN2aoC9+S3C5jLACpNh4ze2Bux
+NAIEW68xw57YCLxFH+8g+XrOyAHJx6/O16A62QelyCG33Nlw8D1sKCeUxZOguZusMZrPgE/ugbi
bC/Y/4HFltzTPN1uB3PdT7iT0DAjVcRujdEZP0q39BgtZ02W67FWL/RpjJsiLlUxMbUISMY/Txb4
BwBhoiVViH0AShspPetvr3UpXJiIOjXxet31bsJDknHLRU0z5NEebzsoi4uRcLztxOqpRCCbiql2
cpFDp2k+H6SAPipd6FKYnozUFSm3/uaQ92qbv0qq28dRR5TSWBGpB5c39+AI3gblr0oO0RKkNt5L
ijNIeU359nyanx2HPvBkuZW5k6htaUSxUNxc7+XjNBOJmySghaO+lKjSbdkA5KyzOSdsqKt/wEpi
ugN7CFWJpglmmB8456AqGdlqJY1lYCOxeubazeF/XqpBmOTKfQ6bTlbqQm0Q07WcCHd54/cMwbxL
UJtw5ciR4kdDLF0cZiBvo9AJblQVwR49kWWv/y14t5AJJWBhmbxDRHS5X/gd9c2gyuQjYTnVZ7kJ
Hu5T6npQRDL7Uclbku87AaR43+VDP1WMrDyE7FHfldEL1rxlf1oobywNYj1UoiA+f/buQ9Z3MGYs
0bSyNkbPCWyJaK6S9IsTrbde2bF1pECs8ScFL0PDu/FxoEsSTIh0nHpKlFcpU2oncoWcvOej/gV4
u0tjCGLJlZV1V3NEiFdAqXj4QfnJXV9Q1XyNMEmI+icxof4dtBt1dVKXua5hcsMOmm1uH9ks8s4q
CwknKKMdBIZTxZy2Q9gHKHLAdQoePXztWYKqC38qbeWSB4tOfJ7nKtoaS9ktNRBuYV2ddN0CWT9r
KTlL2J3gUqiKyH+jTR3C+u4Wn5I/axD3b82Q7tTeDLfNtNRmddWgInzT8DEleTm0yqCdcYxprtzs
U67hs38Mq1nXZBNwx0/vDb2yzn/bVlHOqzjNkKeHIIg2XLo2shaLE+A33avMeimC3nHN+23Yznsr
ma+2dV032/zM4uT1G7RJUOQlxJTdiz2SQ9F25TCHjo2n5TDQPMVTU0jJTjtz2+GjEEoMRajpSgYG
Skz9Vr8cHRkAP+OwAgJWjfjBpffLvpIxSw26+NIjPBZUeZrgiwQCVCfpfvGaQi9VQH0ir2kRp0Wt
2RgdfYDywwSqfUJXf2BRwTCM8Wyi2Snl9vLYcg27cpwut1eeSZbQ9+BZa29K1Kbd/pEF3boTew2x
XtEjK5Af3ICLXi3ljyxzUCq7WADEKGOG/hCUG+OF4sp8U8FVw8q7Aqp1zYrHKdevwlFs4dLb6eLy
cE9FHGzzhu80ZGfYEo1Kl8Nh8okCVOLDy5cd9sM3/9GW7Niba4GILToxPtz3Wo6Zv/UkhlfUxVOA
30+HLiWqISbo+rxwQ67VpcNxWIeDXYVGwf7u3ZLZkvoF6KtwD0MiKyc/JvRxXgW6vvMOFL7ZqOsE
xFPEsLjeQZf5ZgkRVFU4U2yAX1OLAwIBIqCPoyA8tVcJvfFjpQA2k95x1ovHNrucXM+cATvzWMBV
wn1myWeD6Bg1c/MuN/nokWeN3RGirxd+7MW+JujqYPL16CQ3QZwgGvc9SwcsxWSIZYq3V6IbswuH
EUTkc3iH5uWwzQfoiTaodSDCMT7NG5v++Zso2GKmwvHbnHV/6JztmzYEn10/KrcmmWnIV2SxZBcC
y7G9naPfEi01UvHQRcLKWvn4TCEcMUY1OX6OUzTwCGM+17+88EPy1e4cfoY/L/mOVq+JB4ruaEU7
UDv1xiytiezsq07nY3TMFsVqAdyxPqNJ0c5t5nAU8E1g8TQYUCaAqOLPp610TxE6nVGaggrCLyUh
8FLnUO10rzJhWrGnmPDz8MBPl4UDqujOFU6GnZCH7fiAS1m3f3kSpOPe8Whgv0eVMZ8LfpT8psfD
idkrTVgGX0Adv64GmOUMAY1UNdFCWF4iJMng13NvNoBe7rIki571XQr/xdIcSQznyAMJ9H+h+UZE
iy3vGPu0bfjQzKRWbVEzARnLkgR4Oi0B/vEMNvsaDehExnBltwboHml+nP+xtEm+uu2092lalZ9q
+RRLqTIg9m1Y7ut6c9UpqYmj079zF0mtrAEDAmwogf7OwWMkEfg3m09VW9LlaEcGZC6UZgtofPiP
Lyvzr4+8DmCdGzA7ilyWn2fS/4FOBsfOtXkwTNWpCOCHE+Z7YE6hknQDAS3vxX9cfJebg+6iFTYc
6PxXvdKSCFdf9A50o6EYKqS+q842rBqy3PwHpXMCeVxNxsq5v4m8TZ0fhi5Lbs1MBwL2p5sENRyv
lCmXOzaWgtNgXsF968tQQdeZUpWTwJVcEVQAnIeZHgSN5Bsy96q6Fr58FgWwAUcg7/6n4lpaPy+o
XqyuD9mErykPG63TB6RjfZ7hN7N4pNj2KxDG1GM6WET1Plzo2x6exSggX5b0VZJPGPJo6WPmQqxf
K4XCrWp2+6k6v3oHd1kRNg6xh2DAZp2lvQKRMrViaKF24oI3mrS5jobyWOWYxIgFSHinxo1RXPTA
EZurTBHLR9X5GegnDi07NBnfVobG0wcRnbX8WmQ/4Bu1/ID5hQHmjo6OiQet2WTZYz0adjCIo2KV
V8yIPVUZCv2SGj44C6a+dPULvrO6GWicK13N8qHUTNouV16z1T1UuMoJYy9ogkVTK+ZTt1iBfbUM
wTfK1wh7YZJ9L1vpXCH7w4liXOtbwWJ3J/aiexwvutzOnajRY4w/M2uRKBE5tJREMwN8M/B5vyBu
T72wqWvIrCA0E1JyBbL6tJMlvFw1q6hWka2+dvgv9mmbNfRXRv/p34IMAZLFtvogS4KCbzJ37BJ3
NyoK732sUl2OYOTfAn/5brc/lVnzYkNXJXQE2ng+Tr6BoZPJdkEvK0G/Nj5wzUwHjtMCrc7Wnb3a
6e/7uiro3nGQUrRWOYZiA0GPwd2Yd51y8KKzQW1HEVux8lKufAbmSs4Q+C5/oF80/AC/n3n8lkuW
abJwHd1TqyxDeasP6NXKKfhg5Mm3z/da+GXgwjbA93EX9o2uAFe2amP/N0TSSErDVkufSfMllP1F
/0LEN0uaRsnkGTgDS519FU/ru4Hq9BX/dkCLe3joeH83uuBRPLkJcU7o+ASu8I9ek2qfJGJdsO/W
7dCXtC8hubg2K+5qBb2dmptv+dQS6fc9Lc1h6yrRfg9A/ZnHqlvpB7VGMcuzCCk0Cyg6LThhengC
D12eH6ZakU3BjFziyQpdSQ2iAEt4b+WnChy/ppKv2is7gVQTIAtnK0pzFykWio4PPp7tZUh8diOz
wShiWLIaz/qTCjd852fJt07NkacMTAG/N8EiYgvwbBV92StiuBGItqTUcsMsDxpoqK5jT1AtfMjR
tpCtyr5smwxsRSBUKLN9yDcGhtK0mjtlPgmUzgxX4MpBCp8E/GBO+Iw1e3g6aL2GZNiM8kg8aDb0
7uidQrQhPEBAWG/H3yGJ7cVhrTBAf7vllLBeGVo3k3x32PSM2y8FUU2xiT/CjmWL09RBNZk90pDH
kdMstxbxkKret/SiPjYOGNcw3SZQcX96Qi4CVgUSHWNouVt+BuSIiG13YQryQbHFAJcJO/wferIu
W9RYxxmLSmdWcUiOhzXse5YbVFI34xm2N6mUVlBnzO/C4SIBb2w4VmT86aKJif5WztPep8CDcoyq
6fIAQCHKVKgbJ5jlqlzQedr6X9a2s1Ald3JcPYzYQS3/tF2HlhiOGEE07fWevqFQJTvB/DXgDUPT
BWjcq07fxmalOU9vOhIxiF+xfXvHO+cmB7jPYTYkQTiVJ4EQ4zxH1hDExIgwPd8NdHf1LB5GvpBH
kMN7XZn4YAjt7+1qVS9CkLXJ8JoS4JEhj9jP4WpI3tkC+Pwtq1qAdnpIVAvljB//A9AHd1zjq/CR
rMgZUCzI2+nIIIqffYDpwubx0lfEgsmTIkZbMmLsBwjQBA4l+MtJdxrVgjNZkYrq1xXcUoLNW6JQ
KSzEer4cDMdw+9UhlpKZMJF2BE1t1q25uIhfDGGDMAqOADIhIn3NTAyfxsMHPAVwLCSn9pxIsJNI
lZKtfPYhdh72MHtHit1QAifEo8lMG50NEiqiiNAO5I8zOnnmtFI6savWGtOZHJS9W5iIYvW9U1rD
SDsgGJIferg1fBNv/DH7H6hejhqPUQDVQ4ySZVtLD7Qzo031MjOjvyjEaNrH7jomzekXNNmaV0X0
X0iBTZH0OAmeVJ5/4wV3h03OixztQcd/PGl4+F1hE0iduNCTtGr+T+bw116e32VDifujeXO3c2gY
ut/JnbdfbJDbKr10lS2icdXxrekL+N1u1ms4BB+VGyzK0gBCViXZbG1Sr7bkm+lo1DkqB+4CHfLN
5oIiYX94AKzHiU+lLgTonkDrcBNF+ZuHHyigM/LlZsKSRbOnOJSIeCaOcXgB02quT2Nkc9ywj1Dl
5DX3n52X4rli6b1NZ2StpF5OwudySZjVzk0upyRIrzmQTWoxVaGQ+6OdqmIo1HgCp7S0W0NGyM5p
LJH6C+Kq4bZHt7Z86K4zwAh0iu6u22Ty2BwjBT1bNICFs73L06Do5BlZwwOqY3Pl45x7yVHvOknM
3W63aoYEEsJpq7mgqBBL/3sJxKx2UM3SVV6j1Ac1mhKmk9glKIF5Ny2YF5kBHv+5g+V6rM16UnVB
nIWtu3wiNtACmf9YGzzus6adnc1One93OBp0Er51zGlJ73qOayUlq00H6TZoygMnbh6aTSO1XWvh
n+9nYDGSgcTPJVAXzdf7Sbtu5oWOdldnk0dcbuvdMSfErPu9DGNo568oayA8jTDazaGEEgv8d3r2
lM72eQ1UyFJU7PR1bX3dY094ZBsCuiL7HA//gZe4pf/qJs3TBKa5AOAjfTNKmCS6UypMIN/c4Sib
CMr/6MBUa7BCACZ41PADjACygpGggy/QaUc5qP2sDaSajCg/cJVWkL/kj4bkx4gQPrw6v1ltw+nD
KX1j4EWR3GCVmvZtmaPhP5eHAcIhkvqqQLsfh9wsF8rGEuOtdA3bhwq5t1SaCVzsvrJexBTg5Y3V
uSB3qWBLGOhb8I+o/DrlNZx6PE1SS6qbI3WrVpzQ0HGUkFlFY+DTthjnWKHmFLcPi4U2t3ftLLET
tbBhnAN/JqoNZjNYRtQquE4piYARefglnfXRjQom+DdnHMvblNvHuLxYEgapEF6MV5qD50SBl35t
3H9zhz/9Me0nE6DNg2RcD4aaTWYNlnvjXlWYK9urvx9kyq13lDQQv/zQQB2cZzsz5WA6yD44tTLl
056d6QoH7haxJSMDwBRrVp4f9xpWzvYy4oDpppXx3kQFQfdFTVIVscjMCqSpcHcNv3ahLpflqFTm
KoxiMbfpohwIHBWHwttkqS97kY0KDJ7U3rj2DzaPTDAiiIDjyb6n99wgrQXKT6uwSP2xXznXtM/h
Mv/JYDme3+3PkiQViYX7zJh2J6wimQ85ZGts5XsdJM7do4p1upDg/r680LNkpZYYpCzycE2omxyi
ToTh+ANhzto0KWsrwMFk9ee8yMWOuFWoS8rtjjaRKa/M0/u6nY/iJQqAiJ01bc46xMYCPaghPEbP
URvoLc2xuJlSE01cOXQ0CKOfcZS4S//+M/DEyVannpyTpMwpAodEa8OH/k9lhI0z9n8WsxRiBY8K
tl3CtNenNnvUwxCEZdx7arYMgEJ3lHlg0pPussKj7fh3ijZWnCuZ4VE9ZssP5Lu4hLAhacF8su64
yTfrX2CGUXmYp9Yyvs3uQwfbyg/mqUMBHQZyRFvWUHRACOVtIQyfgsSp2vr1xobXFSPABgaenFuy
/SwfNjrNVVQ6SsUwc4+Lr4MT/gOsAMbsjzQyvtvhTAW19Rjd5ig3+6Gn5sTbmnes5ouDe+fLB+gc
81/MaiRLIYihPSBIKQUyxrdXZPRuzDa5GMJwp2sy5F7cPG/mWYT+3v9zN6zDL1BcSQ5QQbJEouEI
8Nic91HnqT5HQFUDoGvGWqaYTm3ydDD+lg6cNHiIAt1ltmoLG+R6xZ2rdtQp0z6H92AFZBfuzU/5
gYsTK8jF+AP1w7dnHT7Zsg6sh0BJBMch0mT+YEldzpdk2PxgP9pX9DOffUtlXCNX6tyfreIjJTIa
zR62cJogKH5gDGTW6KoQYZ2LADZ9MStyFjLxotpyb4heaCjez6pJTKEuIHlRqh+ZbFWDJTbcdfDM
oB7cBgyDdtbhnn5PqMznrTc1N758GqPMRv54LmUcTwBoqwza8YB4Iz/TCMiVnJZJZG7pfFsMeh/s
LBVbKQ1QKKl5SYJTXSwjGTkuvOh0RbDdACN1YoysDBtUnW9E+ZmD2rRGtsgj9IGEaiTTVbZPm/B2
qqFCj8k1qXwhpAN9HsaxoYevFroiDkU6iFAHeWFjgbfn7Bjp/t5mCW7T192hqk2jnyL6WOia6LFq
SJ4yVEJvXnVKqYI+iUghNjfu4QI2tm9RuqyAp0XgyGV2lElI/ubBocAw/KGm/1h0HKBVpTl8gGK6
ci2LakOMwCoAQlC2APZloQlerfq+FYbCqYzYBnAJaJl++dnUsYVOWj8LVdPE4zSEsLSM+kUr06jv
R1zJCpuDXSaOA+egfGRO/L6FR05cmy6aDjA4dG44Nha+c7KsLDc2LiaMxn9aTpO1c2cRFMtUoha0
zB0fsURSKCIjDNHw2EZW3xviPkvM0Fa4xXQjpB6X8goqfY44TR7x4OXX7qSk2W4aeZb8zt0jegg4
pkLr1LwbeDuhHDbljcYZNSovHciHuU1+PavX2ovcHuq0H1NDWmgCDGsFSuuWmdT8qhqiLExszf2d
IjDSTfyVZWbsZgJ+WcR9+Iv5PEXzn9+XLRI2ITdTtlDKWJq3H1ozQpYSXrmsD0XHw/ZDnFLDyr3V
DqaffabvJUJd/Ku8qhY2PiAMTa1ae2cMcbfaNJlv3L8xQ9P+mH1ix0zQC2QSsXk/FujNOQz3+pZC
701FYSDpV5ppbxu410tT3nJGqt119SHhGeYh8y2KxOnaNX3hsZIZ4PtEmM7r35zKKilmFc54IBCO
fDg2PxEs5aXuBuc8ZhIi7/wsbpFI5b/vdpxq+KJnw0gF39omB38kSMmgNzReO7mMo8q/XZXHVaVA
GE/sSLw1yc6nXkw/f/W7QPUHFoSP8/Q72jzTwndhLOpX6y7SBvUaMAq0zO3U41sYCEuMNU4/YbVa
NWHhKGnfid2w9g3a+Ab8yrKdIcPPiKZKuwPFwzNQWFALIGSCXIHi7BbyICVYhuvWwptAbTQJs0fC
uIKy/Fih8rPuyrnWKWGBlMnnwZ8xZl0cpQZ4r/ZNfgTtV5xwIOT8sGqfFjiEUKNvOSII7PzA8IQd
NFmGZzRVkjJSpQ5qCPGB/MrhaWHVBOtTgOnlKo66lNhjW/NZWDQB1Ndu2FjlKH6+Oc/DPJF5lcBl
MzWsOJg4e4BTvGR3oiXmcbpoejJ7xRVFVVU7rTPScF/672wde2GkvpaN/omH6iPuWSe8G3KpzWlz
Q0n1PHg4IcT+fmcf89T1sNLn1vL0s/FUV6AgE6ZelAjml86pQnaCl9SzGPUVsZAqfRjjwzsiU6Yt
cr2f9bWEW16X8Axppdye1/xm9p9zliWpR5wmCQ4AMLFmdgtYxWCW3RNHy2z9qy/oQdmI7zDu4JPg
W+vavZAsho9OPBCfk4mZksNp0JiJco1BG0mOK/Gh5hJVly3LRt5WclTJM97HVA8dJETY6Xb07NZ+
Y7sfYlrMatfusBGlp06q2YtHXNqCpB8xq83EkYxLeACbZkd87n709OBCegE42uY3lF4u9ncn+rKq
OnbnUAVQZsplD2bz7h1qy9xtnmW8LbrbOTNDDkSXTNwFRjY3r9+HOggw+YHXHRHQgxcmIie+p9d8
PdcT+gLUptYU08H2yW334rWobRV1tXExffwrLCekswQGSPiZLKGsze0/ULVAT0OSPzxDuskvJqYV
5d/Ta+EbxXZ9Sx0bjD5K/+RETbY68M5rW7LLIaExcRT97PocWsm5ifJHy3Lypb3R/xYrZSpWXx3r
bUF4mQCqd4LX5jOrWx6g9PP4ob3vDFoKV1P20pT8LM3OZVMIzwmqyqZP8RzNAPljimDPmpLWGZT1
BnIM7oYER/FM+o33uMnryg4AfA2OZaNSWRma2ckB5xzSxfzDE/eRa4ewkzFOpocMCONzPAbLoPzw
S1kScBk2VdwqllGEFp7KK1+OJ4b/4EvURXskNrNgnHW2mZ9RbDUg+keLMlQsUbBIfR0LysBEl6qu
34Ivr5mkKHm3SkRW6zsEYkPJYLTGQllxoOCUFEhl8EEPUbvnpPbiKAC46o2cxkXYrRz2/sO0xyxk
fkcB3m6jd62YzGd0OukdDfLuXPlChaYQuHMeGK5AJdhqgcv+5Eauqg8Crxo46qp8ta3vgY7hqvIS
LQuUSumCND7ELNxYjNUnjH5fcmc6uhupDOb8Va9qst3KXYsOYzXKRqSVsLQS6n6pjdWFeEdWwE1V
gc1/uwKc3uMSQl+Ur4pKQemdXA33MBT+pFSkRY9+JQ9D4NTFBSlUWbEgYBbU3pjv1ncobP00+vTD
sP1/u+d7Z8Hz/3qwppMfa2V7Roq92j6bDPAMJ6cQY+AF2AEEHSgibdCWMMXQq6qe6N/HrLIyM0VA
JRKZIJDzwV7jgB1lF+zL3r1PoyzogpXK33kvm4U8FO+DCQ4DyeqCTvIy7Pq3PUrTd9Yk3lgzkjhJ
eyDZwJ5EViqvtEOLLXaG3z4rixiUKieIOU3Hu5MuB3a03mWXBcl/t5Hthjqr9FP16XQ284wMsFzc
pTEqfkNZuNNmT+Fqv5gD9FKuCBADjLHZaEJvdtCle+D/oLeKXy3MDcdD/Mjkc/Z1ZrEsAPIs2zVx
HxYMpeWfYHrkg9I//qKotYN3xB0BoJuQvSp5kB+xiwY4xUd7Hy31kOLG0f8XsH+gCfYsJOJV6nLt
T6+hioQ3+fpQaZHInd/rwidvlfNj4I474g0f/vthdtpS8fqeFX5AAGTNeTMKO65TOIOkEwkZ5QJh
Lar4M/EIW0JU8kLkafkxfbkHFwkv++4acA5SU0Ez87cL00iCXt3AAICNcBdZoLUFrO3NxYtOKp8U
78fg9G+g6iVsMGVnWEXrZTd/UA1O15k5j4VbmRm1o70BT9DsrPkotTfk+/k+6Opg7Df0bp47qHbf
iOTJLfEmVhs/auQ+2N9oD2J8ONnWZ/p7sn1/YGmINOd3pVFE1VMBgVxUyMA+Oz7nmTZRibF0229o
FaTVPLRtVN3sd2oDfUy/3GSgTpel2McyZ4HjuLP74jpzm0bUepltiRUs/5p9gxaNN21zDuolAa7d
mOKMOCJJMWKxDyl5ni22cl8s3iig7xAgnb6RUcGoBIpcQCc1LYpdeXPXZIafZ8fyCTrdq0WY5uxm
rh84fCAPjEkYpiI29kRngQRI+7g74D8HET34L1aeSM8nrgKjnOVkc9Y7FBKxQWcA4XlHuQ0TKq1q
RG7USTf0thR1S5BLUfQF1Yb1O6AA5KRLCH7ZiXi0qBLU+Sd6Vl+pvr9P1M5byXjIr052FKU8vCsW
OWRhbkv4zfEbrhF9Vunjm857Bf0+Euhu8rlxLUg9e/hPqUHkatFaX0Q8esypm5w5XzPUcTB1zgVt
jAC3JZr9tUitx7VwuZ6bjDhJndi3XLvX9Zg4ygHRdAVjiqQaLsE+JRG7bS+957y2JAyzVTo77WFD
LT314u9yBvyiMukkL9WZ6C2Br9RzlgyRLitYQu3ZQkIisfMbq8UscFdem/pzzEz/iePXrX6Cvxfr
scoVLhc/q4ZqgLIiWHgbPElSL1kGwRrNf/NYkLa4zsv8G3c4vIsWWVcj9o7ypQQMwAm2itUD4prC
B4jAuMqxT8WrqPZpw7rbLyNh/e5lyh2c/kgaeVLGKvG/qRi8xmUYHVvyGp1+JDLcR4XpMSpLqLAo
M3usmn49lcja/odK6nazN62OihnAWbRg9qFDE2LXiCsYRizXFwKfKGrLIenol1Z5cwMcjcqvtNvE
gQTCxktfue83vvm5ABWTJ0VfEW11yC5BOyjCdZHCIgXFrKX6rRFBnAZ7KEgEuZTE/U7ODKFLY7aR
EAAo5ejE7EUhyg+ji7Dn05FqRexdMho8rS5BD/4PFdDvz3zVfnkIRcqW7h6huOTD9rMQMZMIPPZB
aJljwbeU1dm9TCHzfk5KrX6YJykW4g1zVMsELBHMKTrIKEQ90uyV3UPkPCZeZN0FcFvh+Au8coAr
Fpn3oRswZn9WSHApivZt2mBLgEWKd8Sphvg2FVzOnGdBmbgqz/+R7gjsnnyA3cz6corupV5lj5kM
vin1p+4XlKJRHCRO3b+op4Kcha+BFtASzJqE676R5xEgwJA5m6xNWqze/mmqqHiHd+bYzukkqwLu
lwz1jexXO+hDyVcxq8IXHGlImjB4I/iIHX+/tR3o4XqO9l7luR+lTmne/5m/lY1c9OQHqq90TOeQ
ipCXDM80FY1ucPyUDr1i68TRiz7CM15LfO+jkFPxF3mmgeU9L1kVTCQqMxcQQhUlmyS43FD1RmoW
Y7S3jwH4kOcmz6gKD+NzOgFsvRDK9fYeE2JHFl1ii8N/LxJMARD8j5e7NnZal2hbjJvXMUaqNu7W
IJWwyqqP78kT5Bcnf0jWMYHsXPYGWZ6qUIFUxtI5mRHKRUX4kujufB/S2BylfRsXVJFrssk2he49
8gI9Xb2XmTVZoaEGLZRrLTPAjtUVHfVPj3DL4R3Q+SlWRq0SnL1LGKsI9EijGukCCP+2TjbvQxtv
eo7LNSKdoPZqgt/duCU0PX5AWG9/ynnZNYYC8sFM2IjzTSPuTaeSMYgQ0KOyibBDcl2N2J937YoR
DkTrU+7tTEO2rIIjm89yEkLHrMgcEQ3hxnN/Qtrn3LvyPYmSChwfxFo7ZL/maT4cOWTw7wOm4Ll5
DXyhnzpt7cwsk0cC+JY6ytTEEu0InOhx92hMWAG7DxtDWaWdDPUHPZB5cutUOnc4e8gR358YE77T
cFLTm0ENgVxhq+jq3bmKbMex9Fk2k2mJoMRfnKuLatHoP7EWs8jU7y121gniF+D19TtH9qWOnUpe
GE+tvl+NihpuvlPubNPoJ7iMozp0Obm/x+X24FeFjH4QNXvL7MdTRbAyNxw1wdn2gKpBEQM+Gjgt
s9eBokJnyOIpac5HouqUvNbs5zDCoySp5pmPAVgC1S9vlg/O+AIUoIjT1emhJ2ndcMceY8E0NnZT
kNr50KghdWmnK47eEDaBoPZRICSAMK5zW0MplBIF8JWLzFyb1LjmIYLDm4wYKiVptHa4ElbWSTk/
GG+B/eyPP3r/+Qn3sGhKpKjZ9eSwqvHO4MLx6wUdAHyhUZDNElgluhc4VFGiEqOaWLPeczK4Bffb
Agb3dueah78anReRsrvzvjgeeFcKRb45fZqxfpcrx+tbknZb7dEFmptfaPNY5yjpMAYWww2oiOLj
qtaEfEbkiyHCigtt4EZ6n9khU3aMW98emSH6J8oG3KelF67AvImROFvtRTA/NFYvdLl8mBi/6aIl
BGYc2neCCZdjZKfkgfsf9d8qLYvaN1LiUy1mczdCPXxRcH1M6nVA/MdTi+C0rHqONfMw+dVJ0bPH
aMQJYEEa9q8/KuvyTcKNN9yJMH0p1YKm5KX6SaQ6V947OWn3x9b+IKbm0io2egYidzqymdY085+Y
0+nlVOZ6PaAYR/rH3ofj8sm9RSgbPL7v7xax5tmYR0uc2hCPdMp95f4yuVGJ4l/TNr+y6x6Zkb6O
00IGb2roidfQVzoufuGhaavmBhdUqPGVAv/7AOBq1c9bLzaHEzuIDzuouAwe+hmL6QhGXgTjJOCt
0z1c/wRA6nUd487xSBN5Ho8xBd/E+/4kvO+kYFmBuiz8kT7TgreNl7p3ZKLppD/VK+sNF3hWIZoG
IZhoZHTWig+g8krFgZDjFBN/6hmAdOd3N6JbszgBBS6/uyYiOqn50e6sqxlWBjEmg9Rk04uW8fde
GKLonb3PNMewYZ4bwra0KES4a6hd4NKbx5ceNtFNB360mbCWZsheoDH8YolpF03QVv995wh7tsJS
Wx1iXTBb7a3b3AhkfkcaLIulK5thkGl/ugPI2I/eHNEd358/TI4RYfQBW7UFpW+112FYyRNz9d2c
xu8Sd73RzasvX+Gxr1+4qcH9vEoAnm+V6eML89UPVl1EFdp4s+EM7K8sj8Ga1fvo916YifG9Nidi
HL5tlqu7bYAe2mu4j6AY7KhP/+Qtek2evKQh9UW8gITXf5f+tHefIjRsVCPi90bQuw3sthoaoCd/
6r4TRak2yw2aqnKjmSFXQ1SBg+MWbRu9/1jOcBvNT3emYhVdS0jZfzQA1E5Evcsv+LzYgnSlRkvc
yUluNwx1qnQIXRtXkxzdJE1k1GPE6UFK13izX/6mM0tIYb5jfQ+SpmU4XHdv1GmAqchqn7X5+bSZ
9sVgnf9+H2wKwVA7PocYYigdCMFzdtLYHtqm5nlI66FrsuJFQvrGex1mkqzwz2zLGa69DnuxOFZO
FNq/BhYn1/riONkOccRZIbgMSTyTmXKETp0B3Lh71IKmpKN7lDBrV/PTUAPP17tcwtXj59HuPtbl
K6ShsUgSzWiSo3DEQ2H+qmovnh7roFJrIGH5cdiVk2oX8iPSNSF3KZx8LcZSSz48WjSo5+1woE7u
KEUEh7SGN2Gp/ujBGeLzOB5yTqG3NYe1ZblFLZgGK07hxHciCprQJToM0tdQAOez2kCrfmnGoTCb
6EhObt02N8i70iThRU5Q3nFSDxU3suRPKH16KTv79ZHPVeikdvF4zgxhFw/wUtb+9U8AhcrLB/lQ
NAFSJzs5d0EjxrCPF1dtkpS0N8MbSZV/U4m/2fbs6HlQW9874sEayh8TaJxxwc3Rr+fF/9PNQ+bS
BijbHxSie11MzHHmsgTgkXfYfT0XRHs83FrnPr2HJYLzfLvQ7xbUH1Jw0izzYvanA+svrzT+LDub
nrdB3myVmaKo1Zd9tsRv7M8C0+aW3YJdxpv7G3EPxnecaAhd8p7UMbOgOb25cPwg1fO3sP2P8Psm
+JWTpno+CGVBwgAyehjcZoOTv7inFeYf2e9TZeFLY2AdYLeakAbLfS7rmCzZEL4KH2XJ55CYaWWd
iOlVntrEtxqtuz0L3pMQfeTOpsEV1pbR4bHZV5ETbv9HZudSokHsOnXAUNA70kIrrNiwaUHsDJtn
Io/eFaY0XC6arZrDeNN+SLzryQeGv2MeWl5vUC5307VyOCArbBK7GaBdtCQfSje3NRCBkXD04e3S
ye+MGYMLczBp43o+cGw9V/7CwW3ssRstSn1gI4rT6OiJThjhpxCB7r3ILcd3P02yFLoeoMV2N3Lh
vCryA4Oqf4aFTjTF9HfStk2OqeokCRDtp3Hj71+1yrEdKYgzdc5cc9nWnUqU8zdJa5vmVdfazqvL
uEZJtwwRelbtOKPuLLdzD6PcjxO+DgWm8X3XJoO7wJsusR9XlShmUk3cbaEe/t3RjD6uO2Mul+Tm
19TbtbKiiHMJUux9Ojoh7TxVwOA6pWAGbr9rlIz1M4lbgG7FFRZ2B9CSiFf9eVjcakC52leU3Fxi
Q0hRLqNGayy+TCmz93pY1mwSS/ItyYbUXcD+lKLsCt+nek17yYGTwz/czSOX+ivppXEqAYJjzwKx
m65QbspNqQjORDBsbZeHA7YG12G+ahU92TkmxSlOaPUnKr18qZgjL6TLVbHsXZQsoiWR7I0ROl4n
+Z9TSuiidRx5SEdqS65REZ2EuvtCunksQilRCk/RYHP6PFbcy+YkoSv+ov1uGLlUGa3BVGdbzfWv
z5Pjlut0RcVDYBLDw5XGNNUN+EYtGcSp8Eg2CPgqEdZpShfFjRnEBVsuADU9171eh9n3c9+joiXC
QB7Jq3Hf4YwZOiWpdln4mMkgyzGGAKIOUIq+RmNij4RNf3PjhEAktsE44mPN5krf+nkK2AZtWdRc
R5KemyBgdnhOFdkIryn2iNe0iewN1NZaRwmMxvMZuZJnDFToikvBWUmqIyybn6geKRUXcFQAONz4
ByQq1kvmP/moux8RvSZkJdCiwp7V+mfCBehypbzDZRog+hFx9JrdJak6gFOgpeGNJVJrQYCOLwfg
op/Hf4ayv/fjfnCUtWw2ls+Q0SkdeXXBINkwQ6pbbJeGOT+Hl6zBKAS/P51cz2RTSno2yGrlFmsd
UHp9UXrVdD/srZ43drAW4B+NeyQEqFNlFKvqaydSLrwdTLmyXLaZ/cJZ4y5xD/cfGGEeAr638c1X
coMW+SCaE5JLvTEkzko9U7PJkXfrUCWxnWuOofKvtzBXrTA69XTbHT0LA4B89xKs8n7e9he+kHgc
xkGh/F3+fq+eudJYKbGxMWtYnSz1y6qdFc4n8bG40HuCQPv99Vx2RukbQC+ifijh8lNuZKMZ0qNC
AnRnVe3nl1bkUtvIgKbTkCgynJxUlcfSr8z6BZKcpJDP2mXyzowdbcoPSJkMpKQ2VYWzcXC0mnAF
BoWvD7NAl6QVXs4NR1K+b9TTUvrJ2YlGDAmTm/bgopulnKj12WzpReiHRY8r1jMJj8PTfG3NrHZc
aNNQAjkdG5pXcffgpj+MClnk/vA+iHwmvg0wqFzNwc70TjX7/5/SLOgYRIVQynS/fJEXXxOLmgU5
6gH7spHBrcURYX0F1NWxYNDCMFCSg6hxBTHEIB8mFY3tNM6bEzMwJpIOuV4LIHBXxnLfdaYvUIIC
WTeWao5VYU+KKlnP/fKF6GrFqxWToJP/JmiVkCCJbATnDQGxiFOsXFnD0u3oGksoi2yh0Kcii05N
cs9s854SjkVmiiBkVLitxNM15eGFokjDRj0VQHzsDIARJ+d1IsgPC8WT9EuIA7ksOTUx2Nlkm8LB
NHP0TG3nuNegh71ZAp3rJySK41Vz62MtXOz2Uvgec+UFtY6cac1x4DbH65r+dOoP+ACxkKWRtDMT
hrS1+PaohWsMdMEF4Uup5nXy8djypefuhYr8NwhOndtSkjwWWXczikVl3Gwn7akWhMtT4ct2asRe
TTwjHz9K4XC5iG8HnBcZLLvb96NeV9orW7k5QAmyaGv8q/KfoNRxNqmIYB+DQJj8zmOsDN/ClYuW
1DIRg8J1qo5Gcaw7UQ+4WgObA7loaj9QJWLSIWYoZl2fAJbzuFu/qeVSBOHZEVx3OCj+q9dEEILO
J+10qOPeln2GYlQLR9Kgncqzj+1Gwe4IT4HX1Z2SQ8UFtM2vmIG9ryB1CUzoTokqMYOcBK4XJVV4
SXByFMVXIjLKrG7/uGVaahyL4dWCNtShQOKgBrEfT8hQUNj2+4H3uMoUtXXXsABiG1qRYcE5g61x
UNZURLDmNtiwpUZ34rFOD3DZsPm7KA9pVglBNBX/YkUJFDJIhRBIO6VB6wMiEE0p7uHHqnZXiUYv
vDxgvalO2a1WFNpS4kMIb6gXRZr5PfXRl/wO8ovVcjV++bDsZ9WfwTEWy0kREASFDJ74VpW1eKQO
TjU+ZyenLpwf6rSOkKkqXEyyToJ7YovmHlgOyPYfVAUq8JfO5w2tNMVYtYyjf0yZSbDvFvTk5u68
xfMj3cYfR+pbhlL8JXQg7v8OuyUioEJcQfmuY3UL7QT9ou+xzaXm+GQgckF9FT54HLhSfx4rmcRU
X33DQYG7e3GBt2/JGc658UWTNQpXeQ/GheH6Syf2DauxZBO/WEB1MFTdzzddoEUIdtF6Z2GYeOgr
T09zi1qdqecMwGAj05GDdWepCG5ao4ogLY3HQXQw6pRpbFmVK0BcwLD28wd28d3CYLyUn83C0LU8
lWQt3VDtczbqlnyTi0IeWa5DSuQ8ynT9Btfh+uTArVgkpusKHj+CTa9mfzFVL+sHN+drPwG1fdDC
MJdzUcvj705fMmhKlch91ouL2MViHNiLzz0modsQWtNaWN4/RY51VzeAoyn9uCH83YYjZ7TIJygK
kCMW5ezAa75dtBLyfWU0P21FaL8lf6Yj743fu7xuVDT4y8VxhiJmY2EaZL4SkLXgyKE0JGEyiRXQ
5rC1reVMSKWRcu4SWAKaQlxQfT2DRb+0IEQ/IpQfBthUDjJaGiXeeZDDG9Hny07Q2brZrO19aY5H
W8YTpSD7LNmj6ILkutQPy/kuHIq/lsS3LJDjBZpecu8R3U19PyMQw+gF9QkhSpmh4U4zIsPfxnzL
Zs4Bjv2FYz0giUoPyU4vQbL/gD7IjSMe+1Reh8HzEImLhDv4EUzZCgfU+hjECFotaLNXmgKAzz4v
Q1Fg/5FyGjfQ57lX6Lk6VwJEjXX9XNFMhjmumuUjLd4cqU3pbltoLhmWSG5Onp5leHGmvjChjtA8
YIy9X2cqljXq9dPUleFN3VFPpNkLqRnznmx65WrUK8J/LkVJaxVm/mjTsUxciJ9zWl1fECp+Vb+p
x0ui4kaYbZPl2Tez669B2l+h60qhOOlHVZuOGWT7FFo5eqA24tcl9R5KQNIsjCaa3UzxnxonsMw5
ZpLwIN+lHBwDEIYOBZepO1wiIizj7f92dbV8WnitFdCr4xt3BH3uKnaDIUsyQAqfm1sdrsl3t2el
XuWDkRLg3/VM7AloqfNa0wi55OgyLKK5CYqvdRJAPn060w9uFn0LwjxNU+9jchSYlZPMTdrvto7t
F1vdzyMLYgOM8dplJFe/Tk7FmhKdYbHDvYxRph6ofJrtAqhz/vma90NA9Ria62gXw1GHHP4W/LFq
zMMTb6MdABfQGjgDx5a1NxrwarUAAaPQLHp8ptLO9ADSPIZJemYkBQm0DOQsAs1UyAaXtVLdNOuB
IhhaynVKgWF1fBrDcFMJ67FuMSHqps8nWe9XzRQAOf1zJ7VEJcN3Ngb+gr+k3M0nnJ8jamKBnoBC
MNkcvhHMCPZtc0MeFhLQ9Vu8FuVV4iuGaGMxwxfLKSwoW03jN8oJoXD0TqaZ4oSXVNcEcDhbi4W3
N8wtOOHG58O1u+MRLYUn0Yop1lkWSjupRHz5x5jWar6aPUQagAnXQhFAN+ksXoXdKhkht2EqdV2F
uQlVDg9libwH4jjIb1ppID93/bjMEMsuKIsVPVVb/4oYrAXgQXAJ45OqFGmkPLEbt/ZGhQttdTen
AzG+mfpuJSoox6mPYfH7/V0CF2Sn/ExSYjJMQewL7BlWpC+CRGvULEtLoVvGKz5hvJNXQwUvOStQ
AR26AwtgpBTm4N8qXCG6hI4SBIIOQ7JBlFH0tFPBF9Q5o63k6Ue35vyYfgMRU0LjIcH6D2X8vnor
UcZoiDkIwTMgspVE9PnKStgKNQ2S3lmLVEpNDNlV+Kk8r58xYCxHjtDxO3SyswgFVVC0yUFEVQ91
KK2s/8U7UuIo9dHeWZyn6VrOEMNgQ1RHOe1oWft/TRWu0pIbV9zyWymUUqxSBDn3yYq5grlLzFnL
Fa0tnDCoVMJdv1Wod5mJTmwrNHDXqCRagYNjXqNcNSj9dC186rHgMSeS9/OKvFHD6JWqQrJwG8to
DO7l6n4W8nNMZpa0RieRWski4+LqDduMsg0ysv3kQDHLNY+x4/D4S5mqcC5XEzzFbE9uhGMANOH9
0bCJzeONvSQ5VDDJ1UWmDyhTmIUtPU7N6/FmJcdiihxqKvrmf1+hku8/5UFJyz9oEUcEx/bo0VkY
qoNcypGrW4KO0ptGzFAlTagM4tAn7k0TQSxqeKojxlDEc4F1E4/WDEVPcXoTkrdCFaPMcAO3bqxm
c9LOuxQmzO/RYmGnB2xmuoC43oEhXyyOQbgO0tBouJic92oHuYyD4bf8sa5NYP7nAQRgbd/3Eo/J
SJsDrzBwM5i/M5XXVzluCV9in9Fk0fS1s76CNwVBkqQ06irBoGvVV3cbhL1lN00GeNCCT28arsbb
cAbVd0l5U22/Ja8pnWDOw8wyL7hHgcYMXuP8viKUa17S1b4EzNbUPzK5+T3AKVNyOyTf1/Crvewc
J+kGsIKGIZMxpJ59YM//Y56MafhxJmD0XbbIXtzKY3dP+HjL13+BFeuiqGuL5x9tsSm/a0zlMiK7
axd0WYIkxyMfBOu4Vd28RoQX1OgPlweefPMXdG2F5c6RVxVK7J7a6Xf/AnoTpvFTtW1YAXb1DSSA
5aA7WxvOjHuhuVXgBcqiagYx6DAkoEBasUnyTcb/SEnZHkq+MOhaRwu6FqlrsySoRMrvPd5UydIo
U7j3Y/ilfjN2s9mXaFOIL+AsLgirYTpVi0fFAkZlTJA+oHQ/Z3V3S0O4XOuciztaua02iAoszI5e
HkqOkMPifpLFCJ2CQWANRp9KAO8oi/olA2q3KYlJD56ITCm2JaHyWvXJ5ERwOnleWBogAuVkYery
gvDAcNeUHi28xmmSuB+sNi8f2fGQw6gJvDA13BWoaf14I5us9lA+khnSM4C8EOanBx3IyDMHbWxk
eUnBfOKbz3/fI5GM2/1tUG4WiA84FlBkOgxMVlC5K7QYmLX3oZ+UQ+GK2lgZlwLgrnIr0pTAe1ov
PBT1BwUa52x/yEoNciuKbDGsM9Abj5rD+KJa1bo6U4iR0ieKHeUnNQAVwxt7TIuAZ7lh6JY3uBmN
4Qbo91dUkSSh4UfegnOVdvJBFeEvbhGQnsuA3qI3RWCJj42m2s742AjV91sn4bQepY/eUpftppKE
bNczjmWz6eftbtyPyhxe4Es+yWecKhAerX4yA/0hq9//2mazAtsDTPgFHScfArHxHEiNi/NFfe+W
Sb5TK930XvRMsPz2IEkxlwWaakjsSgY4CFxqKL8t8xysZnGZ9ijW10QLz/y4SGhQ+CGJa1JPvhQe
rzZDSiweOu7arPDB4gxH2E0c+/an5dCRQmncbeCoiZktLAylZlej0LvIpADH9EIJe7PdQim6pbEo
yORhBA4oVymAipWLNAWB9maqETqs8hg9adiFKZ7NuMr0AWPHL3L21UhHySxkEQ2c2KWwdFUits03
NmNf4n4JIf/Bk2+Fu5DSLZx3GGHe2WP8s0taeIc0c159peEdy/SuqBfyXtyJGnNSSCFDDB/7L7Y5
9BPE3auHPTXyzhzKeTQvSV/pPV1giao3Mu1MUWBI7GP152pTUtVxaX5CKhBwUqASgCFTTBdgzat0
lheYiCrwRzYVtUuw2miFaLBVW3rThGnTGiXLHCz2EAevXxcSTipxd7N8i/bjZo2AlTrpDqqb14e9
Mf7bPgkv46LQ+XAEn7S62+s1HEG0LOLC834y2KnRxtr91a0j6yIvuUCJE10kkIJIhPuYZzjlBD+W
tLQlJ+NVvKwOj/I3/eK/3PODzThT5ZYfXAMI83n6v8TyYwFEQXvbjzKZHeXeUUDYhrfBQORs90BD
GBMZlytZZT8YGwr/pUJIXT5foTH7U0/PjGl+S5K43PTR6tTSn6+UUXbs+S4rI4Nx0zTezwKRLJmn
Bm4w+2KyDS4F7FVr0V4PNj5wGo1mVC8dpokcgCudXwCZfyj+KxuzD91+P8pdfDkNYPLc2dtF/U0M
p7V/4Xsm2S9FciTAP8TcFuPnyhgzpTiBmlc0E3prujhog9LtEKyr5Egrv21JQgQYelXFx+/ppYKt
AYI/bC6h+dsK5JnfUjSG+TBLPtiqqCHByu/zJwlg52qijytt2L8XiAHK8XfXJUCd6ImYJI05Bz1L
bRJJ/U2qsljLNq/fA4y8ZfTNHnKr+3C4Hh7bBArUh62QuLd0aHeUvMqX3ymWWTkr2ecQpGZ9yugj
nZ1N9LqyPkcSxMDbuWcViN5c5lTADLelYPcyb+wKfUQ9qsh6w/LzQliutzh5zS4Miym0hUjO8YLt
GZrrx+FTbcdTqToDDNiEMYNT1s6OJDTL4gcL2meW0dBkGTi4DdwYaS0tE3aZrEt4ib8YddrTuuSl
0FqAIMvsaWRmhL1/aay/hdDTRDdPwteE7fswKv7o8YDVWxTMrsUlQOtYE5Z0whVBmnAtpjquuqlA
ZipIlak7Pt+yGNltHtwtI6InYU8NzwZTt/0yh4by+QGBa3fyEYe6lsCPSx9LUwmjAu/T5CZBPpZL
JvP9C24ePfY0/LLQDUHb1xfRAMC6KNPnBkqA2kKdKBsPRtPzxJGG7+SSyiWMHdpTiDSstPVmkAbP
62RLZSVdtfrx/DSijQU1LgHcdohUJcPeihZCBZLDpsRAjP9AfCUxObE67THBozxd3aT/DeJRW1lN
x4Ko2977EtuRdnw/g1YB+CK7xMuFxw+tbg8248I2hyX5t09qeP3JpUWaWK7FRhY7RlOlDQ8qZzce
3lppVAloqipZd1D94EHluBZwRRIY3uzOBmUHdIbjqDzx1GyvoyeKUPZFVOFJ57KF7ZvZ4Jl9qvg2
/3uW9BmHvb/Ko2SVOEY9/FgY2E/N9jhkihm5zj4281R5wAOH+B288L4pgZmvP38mvy9fEI2ytucs
/A7EnBf+8Z8abz1EG8LB+UYUVq8D/ApnLJoYp6F0ycHqJIzQhAEitc3/2N0dFPrQdflqojXaFrnU
VwYhYfbnTrXCP2M0GywvPXDpwzI8mE78W7Y6VMea7fkVvV6Ub5FOx7XgsKPrKoNerbDS5ZzLFyZ3
0Fisbd4oGf+Lqf6B0IDA5IoR/Q5niBNsjLaqwLIOYHCV0iIKUVsQcjahsPBTIsC2QQ335OFGolee
TAwFPccHxyBD5/k5Rxi2f+cf8/kCWfGawHESttXb1b9vwX2sYOWCAqnqHYu6iZiVr9t3Tvu/5Rw3
esrlmRvW7ioeAQ73EKSVmIJKCSSaS2+h/q5Vybs6WiXMiBlHnqTLbecgtpYZWk3WFVPIeGJd6NxI
/KSVtTS6zC1zJjFWejiRwVkl08h3tAxcxD1gn2fAT1Ca+We3bkEYGI6XZystrWwNoamCYAtbzFiG
rwdFcobcUzT28edOQPFA5nkeQwsaE4NglSB7crwe3wqkzSlac0ckvuWp6D3OjXWCyuywj+/jJaSk
l+dym3cMefEVd8giTR0w6iDC/5ofSK4YLYx3vqmd+qftISWEF1nNh+QrH8Llm5bOJjJbJCzgl8ES
+jaVSg9y2GXvOr9Yd2nn8Y/wbnNm40CeQ1RpBiBHHbKzRU3HPiIe7AI4pBFG9/uEuU3su8zmdpf8
s+66ztKlburnZtG1gaFRwur3cGuEy5LdlWZFgaAfmicq28Fm+L8oxKLN+8ZnXrSQm04Od7zjjM/1
gnz3jWDMhuan8mfXBHg4ZWkVJTv5VocyQeDFWMnEPyEOgevCeeUBkMZ/yKwO+TMM0u6OeQ74qd8C
hQq2BAAfyUe7th/IcdSXF7/2jex1r2p3iaWdMMJ3pUwF8s1tAAtclPn/7hYQgQjNfcqhrOpTZCqG
fTYC6do2+r4DjfoTGR7OA9CQpv75dgGDbnaIWZ9nF8elhzP29R2Zszt7ejpXShAh7yvZe6ohkNop
BCEIApWtKHPSQs5xwaRjs3cIAstrGn2DJhYHdhMQFlwquQ25qrDShkE5U/AklY6kgZuq10t3Ua6X
D2es9iIUYXzDIs+CV1Fg7PN0y5pTi9JQmSwZAfACb41F6QdPgOlpTyDYwj1wi5mGfXpkPGSkTfnp
ISkQoLU+jNzKMwhmMqI72NOW4DBtslEK3lOEzZYvHP5tWZsNuLo2no4Gt48gTuNBGaWAUfpbEoV9
LtCZitI3nr+V1HpWkgsuD9g90N7cmMpaLc0hvT25ikhJ92BDWrB771bUod2TyRCmmwqG9p6wtkTq
tiLpblYunyUoUKeBO+RpLjc7ez6CHnBxpTYalFgiY2KItbzyM23I3DxrEkwjG4uCIgJPyztmJniM
olSpZLkyTgvInoBGdMo/VbSit9JFkGaCvvVwuIEKQkwC+Z/XyoeP9Hin/oxakaQteGeNf8t1H37z
T/r74SqBuBEJyhizW1Cp2XkRnGoaDoBtY65JJx+SxAeGENKWoVywfd4VgXYtB2/rYo4NwZ76r6sU
NEid8NIrMMxdt4V5xuDdq/gJsSxS3MudAvXJ3h04rgKMlcx2Iokhg48C32CBXCn+B1GySBFocj3Q
VQ1wn8RlFd+8pafcQaNjylV5BOblekl7bBKvmE75wStbgRiGCcjLbCA48cwzsbIr+GAOqJIOCdJn
clnL0cQGyydiR3MJ/BPtIGlSwR8Ec8F7l9xckE9TiDc8foAflIJ7aFS2IyXetAGes7JiJbbm/NYd
yIO1dTucLfD1/s9xV2HaYKjrrdG+j4YtV/nVpwR30BQOd1fzgkg5dkqrXCjgaRwgwAfvS/OjgZwC
cW/wkuwcpgZmqahEu2kz/fzkQoPoYB+RugSX85yolTheLbanmJ2D+ifqQmsIIw8LHaQZP7QTOeTj
dwYZDNDoMzDT3iuWdcPHg/eEenp+t/G5QA2bBc3FnDxHxhpAfShizarm6aFxLKA770Wz78OXon8W
b/tle1uy46X7AQ1ZhwnwDkkmu6lbokoTi5Y01g8lLAeVpN9faRhLU1dS8ogPS8+faB8PO1uzhTng
SYvsmQZK66xkA0CHHkNuFyX/J0+wv4U5kfFs2rQCEqYoEEdDkBGtkQ+/PhW0R6vCpBwentt+mluw
PXi27qWYU5+nOgPD2QR+YxG0pqWxJ5JMsik+HjKLET0rk6TaNOFkXS0GC577MTJH9WmjnvNLWw6w
DdRuIYk7vr0QSKTAuHu7mHraWTLOsjWYQ1S02ydSsdxvYX0DwBqo0+rof42+sfG03XPrTgwrV6UA
u8eDjcrqCVxX4YmpFxasReAohZwkbith3kBC8G1u3Htr1AbVrLGlu4VM4n67igS1BxZ0hXG/efkf
Qb3laME8wydivRu94jJr/lBXWvlDQSUvGOp+8e591gubIZxz6NuDDlOAlVkAgxTsvbgBkPSh2Gsp
cIPsO8vqkunPE52PyrkQDHoJ/O6rUTqqFaXzf/zm4hUCRhVwXGWj+ubWceJJcoT+3o1HgOhRig4j
M7Je21JWnbq4ERa8FqfvVh5ozgAg/3GH/0WY4wyr72PWIyw6G3XtrwkLC0hrPwnlULSlEFWgWdL7
qBGm6VI8IKViFCeZdPqwwrd78l91tKs9JefzMDFiJxrXdRynCvtLOUeTST6DBtk/4yQqwdy4OTF3
wAq765XuGELOC7NtpamDBkpYsBWXnGWBSGbBbGgZoQTk3sCH6j7gzkh0oacOYAoSAqRw6t8vhtFO
QP5A2J6Zyc87mqeUJ43PUVQ0574/MPvErPHAgBRhSokIAonMAkfGxDPR2sKzmwXp6qI8BYHY9DF6
dzgxrVZf76dkcwD/DFHP5a9A36dyMhE1t7+PN4y6OpH8HubrpivfFKNuqMNhafWP+JDKPcHVkF/f
2+kXLOgiOwWdOJgi4fMrLb+EVbaklSWmyQfIJ3F5e+5XHTPvtu8U4Z5CrHkqE7nJ5Sg+yibKX0Zb
Im5ktk2kdsDyildZNxD4ZyLGAFaIqqNqvCDa5p3TfTnr0U3s82vcJgd+gpXBu8Fj/yopS5WfZ5Dp
C1Kg5sOU7XCuUJcs8LiZgrLKIgYDYJwPcQ1BwO4bVqvPpJDsnvEOlwxm2CzXaBU8Ii7qmHqTJSQ7
wWJ+34Wbeix6anOYIegdprqpi71TDMGfBLaJG1tf4JWBNYD+iIeWYhE89YB/cRkhrT4t9t/azIKt
OwzZORUpqwse2iTnqlkAPInvGHvyBokjt1R6sQExE+7HHdvKY/mneLBu/pObAXEYZ6RbZo87LLoM
/TvQGvu5BhZmdh8iVpAC0rZh8M/6/5nCfH9ptaQn3QcN56c40v0zvgVrk2378es3DkeEnjqQGk5F
pOgeV6DhVhaqcRcqqhLN2wrWXLbVDlbRoAA5/8PCza5bMDL89U8AoL7qxiClby9i66fxFPACSs+P
2uckrXRnNifJT0bBzmjjovnlrtGCw0qamM4ifQV+MIniQdLg6baaogXY7k+BW209XDol8ABhHnGc
2vb9Krz4pvHSVBOj+Z+XjJ+Cjt20eH8xx+7aFJp92kV6a2/TgdEh+mHyPRIA3fEm4A17TobGljQG
kXDqNL1+ZYHGlX0Tf/TyblsqIchs0+LgyQNzIYl6RK8D8VHWZ1aLFj+QBLs4y8u45/d3oAWVCQ8k
TCFF8xoIGBRibx338rUemKdEtUPEg6+1ea03KvYshzUVIjsdCG5QVif3iY9felJ8pkCAN0TcutcX
TxaO9goH4fiLTr6VXLHzOkvdBIpJC5mJ2Q+5OeETimBBy8lUV78Z07hDBNUAmShnP9uNjGGm7h4t
OGbDp7qpDc+Xc1P3hrOUE/TW25KfmI6MCCP+n++TE+8eccQErECtleWfhQ2tAq2Wrr87V5s7/+OI
mPCcngUHhxEinEjbjz3YJ2L1/DYZelSwqb2hqaKICsDGbZcr/8YtDBIXjQyg5t99QXZl48nlzimK
dpdJW17CjvfChUhFPm7/ehTiA5CFugQjTGA/5ZqDexy4/xFHOFHlmrgLkLeQpmEUGYAiG5mWWrgM
V3bZ+wfaAbpchjlX28YTKCC9EuWr/KQ8evqmBn4NUK+ZKJIajfQBP97aIXcn+YruhyvgFPYprE0L
f1GgUFv05WWfk/Zt5SkZo6i18P2i+J1Mat5vVO3tDDF0Xi9t+iEFo7JHyt59Gob1Q0O3D0kJ8eVM
u+LSOorLhxiE/y7bzRFlGci3gM7TVzn2oh2+6dkWvz22f01k9TC7uLeDbrKNH8DQsqPQhs0TZVj0
ywd35txTu5v6DqR/TlzuJBiMti9ZYuZY9GQT14weDkEwL7i2UPo1+mgbDTvRyKlVVFYqfnzRDxma
rD3JkpsPkJwkuBil+q+w8C8o/mZXDlp9HbK4hemJ0uuYDpl0Bqol+j+SsmYS/s16M66X0yHIymsi
urfcC3+QvPfUyNqnKiJhUWbzQKCkT0mqqwPRwCoseINjYZN+Ax3kzqwH8A2hpth+Nqyx4xvrwZbY
OkoBiFoTTs2GgYrA0E4/dQF4CnnrEOKh4ZvJpu03bHZ+DEYDl0KDqfAQucUPWtGvyW6ZV1RMBhBJ
NXAP4rfqmm17o08Q79LwP95mOa4zK+MzhAar85oFHJMAIuTRQigAkthqXhxQzdgBH1sKhh1pV8u8
so453UbYPrb6/cMEOQOndJJ+tptY/AYaP+IB3GxM9h4OLggWz2vdFKRub3VfC/mhlJvTCT1eFMpk
9UO/OG08HjXpQ2n4TddncmBtkgGrP6zZeAfaVgPbZiWz6mW54gmjyv1nNi4ZuJWUgNopZizAYtMp
2TUE6JM0tSFQ9Ez6UdGw1S6jKhFDiDEMZTGPHB9+edDUq0jvgNefPgPOuQpG7dCETPPXbqIerohX
LyO/6Z+CqUfGtRkvDHbizs1J4cQKyJhuHygG4xfS6EeUE+enJp6h9MNqijzU1H1fT1cnSu+xFEQ6
VzJDXgVtIgEDX/qv6bTsqyHQuJi10C/YXDni4X8GsIx0KZE/QKNjeriE89X9gzHvf+wH+AQYEtk/
ZRDPGqOkPjSyR6gswtxZVBb0p6RrSET/dwU/BjaBsLRP9IwoCj18UosaRSyknzfd0cdBdot7yL79
ryM7BgPaPIuWf/eUVHzFMa9GFEdnHrGnVYNAyUAhOVCiTuxYSYPpLdp4Dsf0boQmfomrDgUw9TK9
RNjZF9gY0OZduTSFQDIXWM5qG6F9+4ZCf4v+PbcNBWGN7GksPzBjk1tNVrXoZFC2snvlKZ/k1KHx
GIN0DuLMQf3OibrSGA9/+TewH8B7iJkkQ9AQ7WFb23g+THOlhQg7velF7kq2u3DwAD86W+kZR4KW
/wnsetXg6ljIMpKfsvaIwp0SzgwQMRddy8PMqEmAOx4JnBenfVYeoXWvVlF7sPe7Vys0O/iwBq9F
rC/LKhGpIkykJuCHF7rKMS0PgcAxy5S7TPE4lz1UsBUrw4bXA1ugRjycMZYPCCJgdvZi5S2bpxeM
SI8vWd/PooSP8ypsu7xpBzj5huRFZRoD99GpoloH7G+AL5iuxadxAwQ+ZtHR+yfD6/G7Dspr2Tyv
YZkBD0bA1bOgn3c+DPB8q3A7RF6YJAU4jt/zDycnYJ/sF97m6SOab1a8I9mhDs1TXvNQP0sexyax
ZtPdt5sWtOSi41xFjLxzmiJH9mr6EvucQZapSB6rrUv9X1Blo+1PXkFDn6s6OUeFg1Xo5eO18KCr
nLZ97MOyyf+ygsKfP/H7FQD4PLnbZLMrwTbO2cX674qUJkCEkUz1ZU7qv+u/4z4Z6L3p3NQYNQne
PPqZgHhkMeCNOX4elTjMozeoxUJxq3HEORYsvjoypU3PVpT/vgPcM13+eUplBBhuhzwzTmAs9e88
C1ZBMzuQIzfKg+tNiIEQoU5ZKDT3RscQx3I3UGQ496yxi+WdEhN7AJ8zSMmWwlvHdTIxmG7OtFfM
QeMeGXFRstqNHYl42zYGgkIIzfU/oq6wc7YhLkiSn/oDk3aSI5Hy1uKhjZFQCu/FXvCXm+y3zZ9F
xYzKKEHiZ6sqlB0pixITFK1qJmqRHgYEmkcMcJlNbCgp+m6hBWaTU/EfPuL7DKdyEb+cYIRb0mO6
KChSsQMCz383QlKuJocQ+szGu1dRhPpRRmG2bteEnybdTv1t5KRLrVFR8jZwmVRPDhFIOoOV6DqF
iktBzx8OJQtx0E6pLXDtxf/Y3No/TwYWRSB54NmzEBsEjBcelna1UfhATnFNh3dK7Hs25r5KVuM6
wLj/RVj1haOJnZWtDk1jSM1OfqqLHa0O/AIa50hNze6BiRBMlbJr+9QHnKPX4weJb7dmQca3Z38F
dTD+whhB1z5a+Yi3B7oSdJF+0iDwJzEgVqVuzfo5wn0iTixevR7VXffpQ0M1gSwVlkVEZZ/jUlOx
hmGgLN28uRVCVsyx0zhhEPqxffgN1dlvLHk1gmXQyhp4u8KKyFtSsx271OPvxfxnlTcGt/8hp8Ud
ScYEOfSIXU0Ig9cQ8PcWTtS0cHwT8r3cwDFvAjb0qCKQnlVQT+l+q/7jNRGkOece98Tf/ZoSJnfq
ZtoOKqdnQCQX9e/nrdom6rz3RnRsuFp0ZcfROHtStgVtkgoFzCeb4G9O0W5ZIQetzIhqIK7NPuFb
64M26N8RofN51+TgjxJnhndn8WVaKK3EnzPA2/rse0pIPTrNsSSwTtPail7tOwDpXOEMF2drHela
/tfhgnRsUCpnr2i8Kqm3IVtlB1swpUTgDVFNNbIpQnVdpZpsEjOTTTDBCFnR9oJ28W1JIZg6QXVh
hVBi2nEELIkXVykylmaRm6RTUxgSby3UpDHF/SZUmdaxdt/W0pL+ZiqVrgLGQisUNtn+NjIbLg7O
63mKF7eNdAOfgsDS7ka/B2uxg89eB9og6gotC3OfCrncL04rBEfcviV3xBvJNPy5Ywb+3FjNxkQP
ohQ7b1HO5xwDja1s1eTLLyXNodmQEG/c+0koE9nbOSeJHxh42chO9M6n2PGy6HGsEJP5OMvaz7h7
RJPOQteKYH07Ff2aTMMQrPPV9HNxe66gADbMG/BXfjzrZKutXRaElF8Lxf3lJMLt+FEuRGHBNovj
MD8ODyuglK8uT+ZGFaec3Vd3vIce4fWXlT4C31foeI5qM0aTO7rIgN5Wc7cskE6o2rNqoHLsKEnA
72tj2GyqTDBR9dx8uUcPWwNBqqncpA51R3XwB6ZCv8bJkzFGAVClpkU31TU0kaS/xA1KezfppCIQ
TpgeFfuCAIY+v5eERDH7VBnK0ArX0EFU/1fqicJIx2P6uTx29wTuc89N/L4Dj3QkLN75b5u/fO+7
Us444gPK8TIWeRfu67pcq4/JUzwlxMOKgGzddcYUU/XULo2Z+opM2ADnEbbgsqFNUwNRxthwIXaK
yjQdtNL2edlg/jWeRvjmtZ7m60Jo9a2cnlR/8CKzImM9+LFpyFg3NIol/MG9/PQF8ERcPtxA71b0
T5n1kgybu/TKmXNP6WBRcLrXHE7j4oLUIeG1LDTlawouRwgbJYxhe+3AROck3aWk6xwuCoauNonA
5LkljeGhOAQlpjdn3u7IpoUNpUf04QLCWC5dHoFO6Hnx4kLcpJsujY+BpSHHHssjBw88a31+jQBk
XLWb2a/+MyVVRFrhTENQDu1dyBYmLNxzKJ/OXc3honLXNS+EfOOKxbpXexHfDngcuod3aLwVbvoA
B4f7h4NFEm5jE7DEhI8DxtobOuDCDSgxRNNod4XO/SPY3ExQalU4/isHUCNDS/cbGVSiIkaWedXI
eQCFl1npMpl+8NlyrATuWMuSdiRY1wlLjeHn2fZj4ExJxJfVJAW1Dst28BoCv0/mOIDgcnJ7SeZC
uFMi2KxuGsOWVjenxj79AftSs/z3TrqR253Qdxuuk6e7/ne4q/oWne3oB1ymz9KrMu5CmzUY2tlq
62CnoTSXgc/0T9uNrNb9yMIIF/soQHSW9px09Fx0CbnVSqrTu7gtG8UxMsAMMVxzNjj+8ZqWj9Jw
tRMjX0p0dC3jIRFBsy4uJjLQgPW1jYtaAt3Hac43MKUt6dHDaebP9BMHSmyMJ2y6S3YX4VKs7Icd
fsitKf2qPcIUt016PyNP1cdzolkChm6bxapmFDV9/q1/V2C0ZaXyssB5LlSromGes/slRk1cvPk5
VQpS0EUByxVoBjIMcNPe7vGKw6FtA7G8yrWZwBGebRGVRgD+c2Z49G+mc97PkUJ229x3HtEBy7ft
jI+XVaC2/saTspBkVAo7SM8xTvp9OOoNyhdes8HFTv439FVOGzpOJ42igu121sPUSVjj1QT7rokW
4iw21M1LH2MxPoj72f+tDIgP8NfmcLpulhw4nPtBmfXTWRAegp7YLwuL5zi8RWa1Q5U8zh2QOBxd
d1FFsWTX5H5sh5pZ1YoCoJnxsnVCD9Lpgg2o3d7vsu+qI+Ep2foktaov5b0C8un+useuBFeBSPd+
252IIWV0EFxSSmH1WrrcFhURO3UI7+ebLwfpAyvKYHVN4jypgxiYHQ7mz1JBAyh0QG29sfc3GX7x
lsgUU9fmtFxWi74GuN64hxRD/EsBb41Z157Aa/wJBizbafbZtvNuSH/6fjwlZr2tAUaEnSlP6GAM
QuojS/m4h1s1HVgC0wAM/ETnp4Av50ZuL8f80rmJfxxPYnQnJkJu3vYj/jn8yoBpI1FhMkXUJSHg
SbcejnOuPXF7SSpcfQJXbiilPFZftP6Jjx6bxMOYkzME/vmhWdUnhjJTPgTedN6U8jsp4D3uhM8N
OFwdJTFcJ6g72ond938v5/wLfkmuePE2cHHDF/oOLize9vvFRIrrewajlB6RE3CcxsPFCVcjC2/y
0J1s7iTKFpRL9Tz3N08b0Mhx83ysqqjXugY9xIWtVr2BMhKMaoMBdOVZ624hr/8Ec/P5AM353ecB
78a3p1XlBUQ9SzIU2k+kzIH8Rz00FhqyVmpuTmnNF6gujXIEjcba3UvKJGXZhzWySbNMVSu+q32l
NcJAoV164ie8CtN4Qb+9iZl/zJw+bB7bYd7RVss+wRwhWHugTrRWuhDQOBPgwg4yY2jaYpZRrWgw
PXlRqr9YexLgNQSH+KAIYWuY8LmPNNdhA+2yaanaOs9pCF/iwZ3SM41GmC9hjBJQp0My0VC9Rjc3
j6v01PDJBzJF5rwVlsEWqPwSxYqemrXlGaPoxWOmFHNky1GvBZiCNJE8/oqYlGsXvbAnED768Dtd
Z2TPti5DPQNWzGxaGsmM+Cg6wrdpS8N3DOsLgG8uuq/NEt3dqGRth83U5HcEW9fcpSBGMiLXVC+Y
HKrYVa0GZtRmT0U+MxHCB8E/Q5UiazG5H99Ecv2xcvoU2Oetxsq8Q/C6k2o1ed/BkyxfIw4/suqj
3IBsJed/qhooOc+OauRkWyXTayY5UMGzVFn6/3FySTE6sIpVCYTQH07vaf7GO8T+bPHplAhviXg3
26yY1T1h+oxX8IJhehC3bRcqGUuEKUp5aY7GorsrNwpHR24PRplUyG4bFCOu1bw7xrkF0C7N+kN/
PvGxaKJt8+PfMM4WZMYl8UbzMVPj/G8tPnPP556bc3JT2KMQ1F58/f2kveenDXZPtGP0KIRn80VA
kJCi2pWyBXyFoNEAqkg9S0XqG2QrTbR71St1a9OmpEiQuZ+Ez7KDBY/bX59QVrSebuZgoGNeD2Ah
kORk5AXV+sAIaRg+0UVAeuP02kj6IWbQZGC5nB2hM4g24a5boGWLY+2YWXDljZVxliUckS4S5XBw
tnqg4Jh1Zb6bJgvFhqBWxDWUQ62ODEgFZ+oDmWL/wzhvKwaFlL7rg/LY0hys6og5ACEvnhbNKIQy
8zzVaEisi3LTYQeWkliHoSDaZPEcFHHAaXZaPZEEAiXO+pNctwnPiKu8Otk+J+cH9TBfVrcSqc2N
A6qrnBjvFHC38PQze/q+jZ5Hg665I3X/+jWUmNfiKlzPgM/K7hPAFlYXGU6zUpm9zL6JwIxlciCO
x8/dBSYZ2cOVTniulKDDvITzQ3b01oMJ3x4nAWVbgfQdE4m7HsPryly+4Nrh8QBskhuPrAVCFWkC
PjdpdIUAH8062Cq/TmQknHSecfKiPJYkZ5I9hGCMUMxffq1ar0lpvZ4/ettGGSF7YPkM7AIYmipx
03CAi/R1wfVbTDjVQO7Y/rfX4IwzgF4l3uQYRnCr+Y/hzLZlAANgMkRhQnKv1zgVEiwc2NUm1BcB
BjSiSo2wrhnBfGy1zUfjA5EVSY9BwC6BrQw3Isuv7HkUcK5Eor1YNEB2zKG7cD16Cx0h3L7wMQ3w
ALHtscKu6s2wXZHppnX4AK6MNuCsaZ8hhr2kjD58yELbVh625Jn68kavPEUUaLtNjiVuW2WfoJG+
C5IXkNsy/FZhQTdQeHEUJvAZUvZxa9TqPha3/KhVFOTz0FSvtS0hOqQTsVjceJcMRhQI+C4J44mV
XJqv7pGcJ58Yhn935/9qlekzfzYl6sq5LinkH1VFsSIe0ZZykNelCXSy3X6yu/25gU0bWEZ91Yl5
iOM45TQdJhsk6YX2BqzO/h46rmEPT5RRqkQUhTg07txytzHl9igLm5pDyV5+gAUGOb3pRerz3FsO
kyBjUWf+QnnSN2YKxFybpnp2xOapO0klQxhs+Bw0qaetdp9PvZ8/T1ID7cYY7YbtyJckpgzBmPWp
guTcxtQwfGpVizV38VGmEokEdSYIM8R2sF4sbYbqsa6x9u/5Goy94ZPA8fftvDlno8o1+QaTQCI5
ss0KiciABNSdeUza1PLVYSkSi9Km9nbGOMbol39khb0VjxFCdSyKMNS40p0OpSI/yCMt9CQiMoI8
h0MrKRC8ulZiXMHQtn1HDmx1Vm6h9GmWhV/GG1ceRKRcNrizoaueKZxD8wDAuAuI8XCo/7dwz+e8
BwZ0Z66jCWStHxx5gHVMWZajkytO7/rbKTToAvnOnnmXEBbYSv23piGuP2GGS3KBkCJDE0I7APUm
01ewxyCAIu8E3EbgYaB5QTMFMilzmWtD5F5FFmVudIfpSEtydbTxnqUx/3Q6442B4sMfomrulj0A
kYz4TyP1PlAOfsUfZdQXo4vcR/EDBG4W94UjQh5ggS6GgMYhUfMtGQZsCBt7NqIEExLMVlvgBWZA
2HeBqb3yshpZVMr+Cl8In9BfDhctA3OMxJRcoaE29nOHworRFn8P6weS56ASfbzpLG6gDw0Cabqv
vu3KJkLkXSay8qqahnwRr1j6Nm6TYsjvNhGAhokmKNZ/MVlhYg2YMXu/qaLPAXp4uRVUYAjxY0lC
RHe8YkeyUYWtZiNKQKZhqFBnE23YZFwx4u+ZMZpzFrTggax5+8KNsk/66qe3dcB7m7HKwUr1CMSc
J802V8EnQNENJvI3I+jrW4zdwTvfF2cR4ZOM1QL+uKCJ8HxB6I3SRe4bSoPqigppa8M7QBuPTSNc
yEjEnHxWhe3XbwPliYrW7YCRyqvoIENR0r2e2jiVzqznLyPtMz8cGE31a6Ofacf6NLzpUasgbfr7
kL9XzyS4ckU4KriMyLqV5ZUEx+9LA2Gvi4wMWkX6w8vVUAM/kLULzck0reRzCKp3MyjqZF7Cqf+0
x1JgW7LgZO280G7ldCJK29gIeqRGDWzEEg2Elxte/BDzDU1Oqtq9LanTFmbiz8FkWSKt4YbbpFJ3
x+aMLF1Oe75cjwxM7LNH3gKefrc+S7L2yZnUggfpO9qDRtiBS7kCCFN5wYC6IGBdQ3oYK2tVOpOI
u3rOxEgEBrMZrFwkan0N3g/lAuwUy9fkotw94AJZsPo6XjtB9Sn64zRWw/8teYASr6t36SaeT9Cs
MWcEjyqUzVVXPOxVOFAD2hScvDJdaOacIr61lY1fyW0M1tcWxSUvYJr1RLpA0RdBhSIHE33kDY+7
YB/05LPBcutwRVgXbV4LNbE0+kFPg9XG1d3DFITdGDhP9q6oK5ELHEaA1sQK/Yhl81tO4KmH9xH6
8mXvaqLpOFteBk3Ubs5ansva6VgrXoZb5B+ixWj+kFW5YGYZYLkjBLC8vh+os3d6Bzrbpn/DccFz
77H15QHXKcuOVrxrd4C2KhhLu3Ms4/Zh8v0Ro7sqYYb8+QaxwgylyH5y/nlZVo75BAlrMzvzidnA
M0j7KPqrHjrF4plyHomcVPicD/MTxvlWdST8C8ZR4UbHDfxyLGzPy42MzkzgF6QxMwRgGxOeTnu5
uZmiPhCYeAJqQyqp8+Idbt8iNhtAXTxcq7fq6fUEYiXNiGEjRB9iy6tpksLIYda8wFJthGujV+bC
hDNsOCT/AgqiU3Scq3sR3DVkegaPBm0jQL/u3d0RCZ1GmFYuaOeOW2yG9NQugnU1wZRQWArNSxPl
0ygRAeRbOsqmet3ePcUIAc0ASWHkLXXrCKZmlf/bXNNZCRiPxskl59PUh1DPP53uMKtVL4lTL7fE
wC2ENN3fhzjlZqilFvxJrK9zzDje2xc/XU/yUmiK32zVAAMFw1IPmbhrbMXyZhm6qoXpxUZNbGab
JSTH9n3PK1LBpwa6Gqk8CFoLkcBiTXjlIZ0/49AxAg+IfVKmeh6kfQHjwsZqlVCRZ30RAJLgHD5k
wvDeznPkn8FsY433TewDuCyvVWSXYh23uQN6REI9leLQBcYAOELTi7G2luONJHNLX2LzYOuQ4bu7
m3IBzmwiN0K7njhpBnHRNGaNjuDdSDIeCTrSkWADNSxUTj3uh9RXyi0oTbkEch0GGeyz8KfgeZtr
+lZ8qrw4PHEz3UPoXjRqigI3WCJnL/NIOWiRpOcvAO9KHEc3qsEmL1YMx1l3u82DaaSr0R1KReng
SznAVHvNHy1Yd9r7XshJ42a+rdEWXVg6bMw132rkPRUiJXYCduvzmw5NIzU2Jvw4xyXdFTJrWx6g
25CGCKw3CN8Kr2NtKZkpuZnbyZkcgbbS0p7xLtpKBuHJGoDe7md2A08+L1taEYQnGDvFrPIZ7HUn
nubVcOcbdZPindM/YwAGaLP6R4ARSgG3cwuhHnm15loN7jbzt6sESgiuz1FjMALVDIWSOdywjWZJ
5ZbB8ufXBLxG+mrW2D7EgmB3h3muV/Z84dt39Xzd7PJWf3tAFAevRj0zmjbWA6Dl5VphMWtRs2KN
9ENfhHINuIvOYCaOemu4Oe7WRROt6+9RCAcSEE545lGKtgVzyk3SJ/2yOl9eaN8uEzIFR6i1m1k7
fFIeJYAKDaHdatTWp6P99yekP5hMe4y8/cmFmqRga7jINC0D5QcO8spVbOkoDXLC3BkxcTn19vp/
9WzER5Ygpsfy4aeCgM3V9eTGOrIQGnn+JycqSZFzjExC3GVDUv+ITpvfwNNcGaXWgP6j0VIBibRH
0xeY3a5TC2vFsRuP0FzUk7AxoQkANUS6gycMP983xptRN35EtuIH3SSvTpITu/padjr/fSs5iCB6
bEaoiIZeOVWMgF3qVP8fL//ziKYW5HT3+G70phUS1qb08acFPMjJniYpSwT7cAFDApEyo01ovk1V
Uv6pgZBWAxA3KBD52fNj9gNlvBq8Rt4L1u6ySEuBVu99Lavpmsbv1u2186bqT5/ba++W7oxW29oY
7WnlurKLQJDpRQbC+YG6TC7RqHT5RndwCdjH+5FTriDEo1U4g/mvCpRODtV/cRLYgn36YwouJrp+
y9S9OdPwqa2BuzXvwerrH3LMjOf9lMZjSUcZ0AFdSPOEsdN4ljGNlhAn7NjNBmLyIEsz2YRDrF55
Q1/ztNmvKYMyCB/XCfpBHnYwVy2FIJXTI92GKS5i04b/ZGJJIe6bHVYJkTZcWrNdiNDeblHAA8pK
PcwWc3jbUCE6kebk6oou7NZcHu9/beahiPgnfHF9qPIkuznOz+nSpdnQBjwwhhHWHgJrlZnTgtt3
k4iOwi6EP6/oc8le1MhrvxBsow/vpjNwMDZL7yA1Bx4JfZ0c4AIzerGcv8RH9pjn2OFuWKErlQUQ
g1IYz7PXsiNQcmOLYfkLZyJJwOxbn9pn7Ly1VxOv82UHpkc0q3IlGMTHSS1A0yL41T/UkPsHGqhW
aZkLWcLtyR49VD1QRJtsW/hwrb7oqI5OG4dOfo2eKbu+k84jNq2w/rcY113E5dmd3FY21tQNDmPJ
Gimev1f/J2rfs7F166eSrLyvE7UJ1ahIHWxMpKYmJIrp9Q7WjjExZOxxZW+IZNqmEkr+jlZwHzrL
Cf+1g6fNEvmLnUowxY2us8MTjQ5jksXXDk37LPdyVGWWBWQelyhjrQ4geNktMVoOGhLNC/sdKlCf
bpaNQZ0W9W27R6cidUsfAmuvzj1DN0jZ6JnFJ4+em+Z9S/e3Bzt/LC+rxHcwonm2bvuWYhU7v/33
OMNadVn5+iB6tn4/QAWTV4sWPb6aybcgZdgy9Oktc0kJt7EvWbYQv+CgYfZPr1Gzq4nEv7pP6wk9
cpX/oYRgg/d75cSn7t3VvrIBGDbbBGQKAeKtLfHa9MttniyF8junh6gUTNrmBKm67eLugSjAbnFT
Bi8WHFPYdXUZRjKsYQIJTP6oKcqL4ED+yKjzj2TyQy1oZi2hfJ6PcEsb7vdT+J3iQvYmDmqeJb9B
OzgYeR1qpqZVKwAkHWMJgl9I7W7uAYSwnOPW8CaKz5zK7z94pPDlHkdBCMBmjPX2ad4KiDCsckIh
ZSOZTysFu+dewGkAxqQ0GgBEa33kL8KZsFhZBhwE+nPOSsza5cAKkNKOUWGaOQ85epBK+rI4PAuR
Go8qtdmF6lNsxsn5UOk7a/Tnt5tEjXUBcPK4bm/TZVE2JpORHy7q/Yl6AWH+L7wHkPxJhSl+9O2P
NtmNhoI2BtnCbfefkLpOTjl09X0PqOB69D6dYndT6xKP4WAP18O6LUmiC3cQimrxnoVdo9CFJzuw
xwSXI1bXou5IxIj3pGZcwxTtRZZg/yhFOI+19a9NbHAmfxyGuGszSiw9p75z+9J8X8Lylb3eCSa/
jrp0Aev5qlt/MD/gMLXrMQhK0nmLguOkp21nlSLzmBgH3bobFa8zdd3aQuIQHkpulbPIoJX00Q/O
qBkEdbsKRbVahSwCZX9BMsFXpozVVLM0slWLuFc5/Y4a8T5L0d4pmIJpbEf4Xm+UvfoVaTvmPip/
nQ4qGpiRmMPupziMm3zzxnfdGe9YGighObxCx81VY67aKKWHBbzaRXQEvyT585y/co6FxO3LS9bH
Gb0EnY670dt4qhhNnUBvtyU+B/qZm3Qnm76/bAaOY0RxfTIZeswzmrzAWgbtStfjTu4JIJeyQ4c9
0f581fkMy4fmOh5Le3CRVUgK7EXbe1v8ZmICmPldFhPD8ztYRugVHtottSASL/Imi16fEAyx3U23
dbWQkjTgnwP7I+oCKv+h21Gt3jxaiw3ASez0wDklO8mydQJwaaM48eNVzedeJ7g+tr9J4YL/yRjR
L5mEIF7K8GUNGxFjHhBQuKLJI/xY7vN8ZcKhJk34iZ70GwP31WexIHs53WGwlG7+wjqO2gd4PPvg
HqKfqaSLV6iPNmyoo5Eq1esJqbXD6ACyy/yM6FZ0UNMyKL0pw4JDmRkSrXmHEHHOJ+GvX9ugmTRY
YXENmYMBFodh/pVNIt5bjkV149bgkAqmqEWXlT2ixIDzccjWGEYtqCWuUckophk9A3hQMMRzV5vk
sXM6iUMx+10bxn9XW2E3s8Hwp98DrSBA1v3QMpoLrFTpT3lD61A4IezAxy7kA1M3jO1LJPR1+go8
TnWXhpXIziELIt0vYD0G9vm3ruern4ZtCl9gvLkJSvTYcbdG/fUvDR8XWmJ8Ak4Q7LuHi5uhzygk
sakV5KrdDNernPnkpl6w/2khuDed74qaQ2q9WybaOmGIrYQil6iEzERSkmSirIqkDVmd4C0TXjq/
s6TUkFEBZC8AXHl/y5ZMKvkr+yclyWhSAvi5h7zPqB7WetLDTrRdSedif5E4M1YFuK6pYIw+rY58
2Y51ZWG4NXTlC+lc4N/KnrNW50aE95T+W9hRKwUI+WbFOcat9Yl25anyL3MxcpsT0nSwY7CTsUaS
gJcQl/tK6zJMKKuzq/JT7s02cu88ACFF7RX2va6EZcD6/5LvHL6qIedwzikIqaAK2/zOSko8nIuw
62GGgEfRxpg6vchSosYxqMz5Rb7qdPmqMMd8q5B60+z7eTki7Uvfw8yXxgoXYIk9tBHJDVkNZje9
LbmNTZzRMRR0hHmdrqhIOAkUG6pOE+N993AGbYg/Lv3fg1uOJMvHS3KaYJ1rFf8fokz1UGtMkP8v
xcw0sJPmBUjlGW4ugesLQ8sAts7rYAJl6pvEGNHRIbzMqiV2kFqVdfz4z2PAn39FXOI+rYphs7d4
k5QXsBIoqlHBmhMSdxC+3hW8xla0oQN+1RcUwtdSs4IAJcbdZyA9VF0w9dNHXiNiB7O5EoGdG8XE
+OfMW6dF90csiUI3Z1UE41dWSxBF6YttKn3p2ShI/AsZ5Btq2w5rqklcjGQzLSacLarDY6frU5vN
37Y+h719+xteONm81BrhTuj9bMYjAcJW37uqs0GjPwLaxlvv8o4EATwLscpj+pBxGYiZfK12UAgq
HbXenonkSLooglnQsDdcDas7Zom4/hM17UEOOB5ybCYTuluDIAgtWv4w6oOXv07+UGCJ7o7uhX8w
3wXNSOAkTH1otNxisCba/Jdl5PI1CzhEAZVT+pDhfD1GsZsKBmFWnjm8DofpQNk1pliOnke5EQ8s
Bvv/K74orZOLkU7OlNbf76akxLkXLmEJddJsGBnI2b9mKR33yvUBeneD6JGyxoWscrWuwUyYYCqw
JN48QNGBaVfQd/3zM4KaBsffQeurp7vYL9pEHEathKD/mUFiChgihRRjfId9F7lLWsl4gDN5K0QV
BXlVtfKcN2Nywkf2gQrb4N3E4NuEE879Kd7DjL+JliLzeSUWxUh8iF2Xi6eT+ZLnRw26eeQHzv0D
lpeZU3YSkW9peNqyUm36Hdmwe2aGYB50mozxu9oSiJ2Uqlq2uY4yIzneBoYL8UeFtgKoQmA1XFDP
V4SXaAZ396SLqPidRmqvjSOcrOOB1QbQCBEHOErFLRbeaTdNHFW+d8RPU4oea1lgk9NXSjhcuqrN
mBusgcnptyEWQh6erhFrmaPjGMBUwNzb3Sarsif8ELnGB/YW/m3BmiGAJ0Vrv7W7r3LshsBWFF1r
01+501ToW28N4uQ2mEczvp1QCGN3yguAmhpCNHQs/gVSYU8fr+qmppaUehEMKw2Bu3Wwge8x1avP
B2GA48EM0zTi5iGX30C+o9xphb/hYm6XinxS+cLfkp6wLzBZfFVZRiMEUdo/LKyub1nOqNjzFoN3
nAo2RMoSSRn3kgwEq75SlmgQEDNewV+rRyhldVNh4jKfa1ZQfemxOZ1+r/gBf8V92AZlmOGhMj66
OKZlpk/znswrVbT3RstBsaL9ZvuXeCTNfzAr9qiQ5LbDCPsbw9VtKxxl00b7XlQc68/UGZCgR9sM
Cr7GlUJJQDtJlgI2IKR6xawbluAXxKbquSi+XE2mlxIugVqQ1OCi8yRqE48PbDe388nZGZfm3sN4
lh5mbtXhS3ujmOalREjIXEQVjhvzYtPHfFxrnWMWdxx1lYpyuZYUQ3GYBQF78bFRAMHsCOIJ4h09
GZRsWIWWELa0tAKhipkoTH5PopU/G7npaXGsfc2ieLddYuc6cJI4f88Voh/kme4ZobA8eMQe++12
5wiIafa3dVDjVq504L8Pm36Y80Ltc+6F5DijBTZINipC5FcTERqGckaNpg9kEZ8hyXJzy/z4/Skg
whekLeuw0MDyWBC/+VtNpw4kOWPZcmTsIM/dZNVf2Jqe0c9wr2ykWIO4RfGnDKxg1wxVw6q0hgpU
aCzIzzqvPyYKKMZ5H2Spv4aoHkscl3BHDbK8C+4Cr6QdtsiP55bWTWg3D86dthOfeaBbYMUy10mK
4TCKnw35xWjpNE3cuTfbSpsUi6ZX3CzMsVdoYeRmEtPULMG8f160uLZR548AwRO+Ym2vIJUrcXdC
3UyJ6bclKPzz2Yflil4SVdpBDH+X0st9/nwOe24dB71ADVJ8lwwkVl9a7uxDTgMychjVHdVk26+4
GDnlKd/DhDW/Z6K4rrahaTGozYUC9ZOv+/91q6ySF+tpw4sS7ahqTkMTYoEBDA6Cs10X2tU/iHkY
SfjTMw0JvSjSs+3LKN5DkSQjks2BUQeiXMB74CheHkrSEnENeAqnvZ5NfigS4scX5KaFXvGUGdbu
mUgAq4LJMiUu6UYw1h+AdMsQtwyR8Xy3JFe+xoicdk2Y4FLieudEswojdD5Hc6485OFUL368BnLB
+Yrowp1P5FcUb8/qzTnEI6yYg3FhfpewRAaJPh2H42/T59YjumZ/5wss9GUTFhsAWbZe2Cv1wrlo
bwtq3CiTqaq61H1vswzIM7PfDDO+ZlXZHZbYamFHMv6r/231dw0xobcOO4LfwXAx47Qf+H1XZhZL
eiOKrawPB7kfA0ga9XuG9bunXGXI+Sa8ra0SaYJwN0pcyhId9fZwemySC85EIfsKcRnQGTyhhs1b
SP9QFXw5Rbqb6SBCK7UIWXNF8+SeVqZ9RlVH83mtZv8iinuqD2InIxFhF9fdxvYq1pXydGFR3SL5
31eMAP4xG0xQpMeK4b87b3SUxI7+LYnuJ7PRHtvCS50RWhk5bVXJ0ufSAHxlEslLIk+n9bXOKuFX
jIzfsJSuXVU4votIW4faRj1ayf1+BGzknPWRXIXOxlo77lJ7MAJJh9PXITFfbzefzKVDWnO3W5m/
4esvC2NMUBBEdFCiNnru9M66Ld0mVVITw/kW+kQfI7qto36ru1K4YaPZttTG4emL8MUJsjJaM4xh
XbTM3Uig6PiSFb8JmaavkHvB0pdhOA73/XJaQ6lt49nNUf9Em6n/BAKtjFEbyBj5cNj9JlQ+v6up
laXRPE8XmAOzUlFJ4cxAtPn4uKcFGmAFoluQ8YXwmMnqjAQ7SkLmPyjtJq19Vic0NbXqI2X/0lVw
jhq6mRPwjPUTZFHjtZNmHRt1/suxMG5Pqswk7/7KkVFzAn5GuZ7gVJb1sUFLNuwF6lBg2UDtVrVt
1gIuz93gQre2uQ7zmPOb1TbEqlZMpOR4Pn7CKjcyGQFy0E9y2PqKw+JX0rRlzATaNU3lWXuxtOCA
7zUlHkTDw7vowzeQgqseXQwbZ+A1tfANwTyBbd6IoEfNaMGA+5G3rOq/IGZzfxIV7oMDmycsoxBK
ZcyfFcl7H3GO0fRzoJoMovV+XsygJJwJ4ub23zgzqpIohuY82OEdF+GiyPKUrHuJC9mbzpytt29P
FeB8t6fmyXVDZlMXZjXaQxQjCea3w5BFWhYk/3Hx2e13D/KvnAADco0WKRwc+3CVzP2MvbtOQlND
Q/TRR7kpOTm+QIT4uk3a2oKZTCBmDkr5DR7hYVC3gg8CNEp0Y9ZSVl6hk5Y68kLvWhbMc7Baz/x+
Rv1AlvA5CfW1kogTX5a2MLk25mvQ13zuyE83Ajc03786gctBIcbVM50lT32vLNnwe1Cpnj10j71B
hRieuId9clggLnH4HVxA9WCOIUrG+lmau1VLCFeQ9wyR0J/4AQM9LW0ZQh1KZ9Ac8f8Yc8Ufohc5
FolYLes1PSPM2XV1R43bMgVy4P5xE5groTPNjimDTb6Z5lk5EEWg1Dc3DQejQBekuu6V1L57yzwY
SLhGW4AeMvMa3q1olkCCwoByGEP2qkeRmu+la0S5OoTH+ZiZtPT2Vf9sExuFl+kpR25HyGOjHJ0I
BBIdotRMeOjVTyMd2TR6A+fo6W0feqCkZLXDb3cSO8lQc8LxDeQ+WfZK7NogRJLp+efpjXkf+Xqt
UuG3GKO976Cb7c6hWUHJkBQz0Nz6GEDBumdikQLF8hRAV0dKxynURuKBfFqQgTOXFFVzR+J26YxQ
l658PTk9ChIzebSxmY4w/wEZJsbDp1gDX7GzsobhFQzpsQthNY9+nKyKxQ17ROb4MKKCdSkygIbM
mW1xjb+KBODnWO5ZSORnI7Ynj1IXh2IDZzsb68zAjvuQK6nEaNcp4Z+btGlwdLtm9QNOoSkJEDGh
CQqrnfa8ze4X6NZtS+aZIiUj+q39GBx7HuldzaMMDMkGaCMcV0LoQ+ZmklOtMStoCSHl4B23pcdS
D6p0lOlwxNIhis9aoF9NtEEq4dU/OzjiZ3va3p4OnoXoTzrvIbh8Ns/hrJFQ8PnZVkbx+IoPLEfy
shk5uuXjW4jQHIthnPXGwcU+vhm4c7J/QbEJHzo8PBY+uuoxFyr4LWiQxIHcrFtRZbbLJRBjCj5G
1/ysKi5KYuuvRRXNTmVKjBCmruvKIZThnnmWXMyoVSWvGO0NYffL9XRJmQVtppZ6tuQBLQqcd4Cd
3BLzXJNySKPexy9kDYgxXrqIXkn+jJ42xgpHi7jWmsG1ekhjCt8+6crWdeO+gf6Y8nAlIrxTaJHE
05MLZvJDP++lyiU5lM3l5a7GeRc4lQKdXLaITdDzMzWdHyP/BdVzrI4HDjX7zYT71P5979NhVWAr
jgF6wpZoEXrwT6wqhu0TF3WuFcnvnt6U85cM9fmVIICpoZk0fdl3SPSX4fOTxkarOEPu1u++6bmA
TU2nLK3SUPqg5jHE1jmy35Zq4q+MhiiFYMrFpVJQ42OB4TKrJGjmx5xpOf+MRjCwyODtq6i9+Dks
b/K9zx2D+XAm4O199vdlhGy4ZwQxoqSuznJIc+ECo8xdXGotC0eRkKM+kMWenI5t/NxhWfm4t9hh
jcTFHJHfAKbw4wW4nE83gcqVwAkZHlU0P4lB06q1IorMLSXRWGs4zpizXA31GHrJ2I699EWUAN6r
msEnLEGi+lpwP7SMKPo/AYCAqGBbJ4y7ryQpgcNG7zozZxKcviRQSKVgbWijr6m2gvWBa+Hg8JYZ
Ba1AOsnKTuWRYvScZNK2Tej1raxyk0QAY6JrO0dhRfIgkDAeqOiNGeL0rhAPcwmk88downK6+3Z3
MZW3kjRPYn5uGPb1lDBezdrFjPo8L6nV7EtvN1d/h2Wij2rdEP2bqMIdVJiMqBECExiKYsQ4dL8V
T6csjhzanfHIsUxu9miSNAQjI6DKEM38VE2jttRTN1ydHz5IX4tGUFE0BkJcTlD8zhnisbzfVaL9
cT8UQXBmtpiFI2lc2e8ndZO3dJmBli3TNun574YROeXV5yKOcKULMoJB1rgRq5QRCUcYnqfzg2Km
MJr5wLLL0gMvWCEebkOOAkI4bFo58bMtlHLO2A9mOwuQAzyg9aEoJ5xswghnh6IRkXKL9ByfTul0
hw2IyxwuBvBOohaD8fGd2Kvwk/MUY2RrUvyLuxi2XaU9p7UOIlCJkfLg/cymxlafcCuM4w58Tuuw
Q3rBeiPgGp44JrKpXTfVa4GsIxceKP78tX5dYPZdYYqs/uN9+qEPoLEO5KzhCF9G96qyZZy/yQWh
+oPMg35lBN4/npBK2GQRYU+d3L2ZgzhBBhJYyoQ0Oh1kSrM3sm2TGVzLMzF07SizRCraBKKzgPv8
fwYo64WOYort84AJj3kq7VYGzwP5yH8WBcxoc9H4Btm6Ld1OM2qYHm3XL267abgUdPJERa0r2fRU
/daRoXOrV7WpSCDTWidJRSD+J3IVpvzczXj014qnRMYJrFcIXVWYNOJnVKo+BmvIrPV54/q0oues
LhttsR2TOlnivcgr74kYCaevJNkMs0uKO/mshXiJ7vWAhrL9t0dO+ksUN+4lZgaUj/j9N9PbqSoA
9D01x81aVVaZHSyUf1v2/G0+wKt+3t5rP/XTBgC7Pt9xc+70BbxddsIH0MJgGn001bA/CJfzJmhr
32Y3TmOY4L2MXJYe7KRTET/yA1VeX/4p908Xm2lNtNAx5FSFlc6fLBYFfb4jVxXMHPHHAPz4j2Ux
Gfy3w8K4ENpwhu1MEmH3eirc4yQJ0ak8bnTbJdR/bUOHiV+nKcXaYt88CwVRkW9/ET+F0GI1vO61
1cGyEWBz3a/AqKRxJVXHRQoo2/aKjFmj7TfbPMH/vZhbhJO4KoGUfNEm91qMOh6lk1Ehk7OyVkuZ
or8scUTK3i3q7sxr++Eir2z7McP3KGujajSZdShEJRtE/e/ioBF6bU+40guOy228RsjLdiXqAnfA
r+AgNEPIjkY8x3UU3NLVBFwm8S0cTXFi8NGxGEsRiZlhlr7yH/QUPjsP1sxquyynhUGplpisP5ZO
M/1hZsHS3bDWDx3SzE4ljXQqxBIhI4/q9EQtyXrTDLYrgGs5kArpYO4ENg/drWSvROABpDS9D83s
NfdAQauqxaAq/qx5BWXdYQahGhZG0/yVXM15IW1VSDGldeRoWFTx9t6ZMSTG8AnNexTkCPontrmp
+nALc5ipBAhjbjviUCNW5ZlL3nA+s+c1+UgfPynkpyBo28JbYmmIabcPzLhvK2CwP5HYKMWjbCD/
BeUMelR9sRcOfGwPFZ5LCIzk2VBo6TTPbzuwm5AClrb6sBgxb+VE+GMNEvHO/cE80e/+MstLUXPK
aW68t6bklidV7DV3yOyDQrZVhL2FeV+e0x3wlSMKPfHJPpzm3BMbBPc4dUmM4TK6+1vghdhQoc08
RkaJgjiYQPez5ECjQ14BpzKLhk+MiHIE6MDflFgdy5lmx1HaPprQ786hrjjrKluTudvNkL351mOT
gotVh9ihK/Hv4rOMvIkMC7nFrUalooqjsuE4R6yz5ABL5ZTiH+0OykTBV9mW/nHbEsRrKxdomZPJ
Gy8Ku7yWF5BWLw3xdrFQjb/N9A6z2caB7s5RQk+XnT9cm8eiO+N6a+OIU8FD7Rd/chK+xpdVeqOz
1ik9pG0PMuDJJfRGb2J6FUucME6259ZXAJRvPyJVtTBdDObDL33tm7RkOjAlgCvQDm9c0KppZFSC
qKW0Q22qIxVRGLbGtZY2VjZOK9HECy9nz2AbNKWXdyNGPADSEqp8OaoIHYq+6tNi3cOg/7dJV4Pr
BqXB/xlMzj67G5ZonHtpS3dStcRwMP1c6cXD6gUDBd+IVIdDXu+Czq1w1ywH0EXrR1AprdAHmZhM
ysqXlHWR2vNlIpRnL3XviEocKeXK6HmCBF1+X+WElm/VmJBozqME887aI17bycPBJihfypYGh32r
CW3v9GMq4szneJVfguwWwJI2QXclByejbUfTcV3Atsa4cDZDzhq2Pz4T7EQnWKzBD9dpyS+oO5FY
c2NycWGnuzK3qm4IT1soAb/1rznZzI1RvrwP3jBvBR64KOfZmemyZteAMorI6yCCqJ0TqHDr23Oe
5pdnOPr8pRf4dPnnV6ZUfiIObNZXyUpViBXCPA7Igc4qn2+s4BsMHxS2UNLhDcrsp9mtpkaFWMgR
/PFHldpgBJiAm7OjuNbJv95k9nc8C8ZAgKW/DfYyw/KxkdPrgTPONGWv1ds08BB0m2TD+sQ1GhZY
aoQ8O8gGhSmSmZFFfFqvAjfXQb7+F9ECDe7H5hXUDvKVxtQR5WYUgdUkAIzi7o/GbqebW2zJe6wM
SevBfabbuEz9API+Gytg0mfODSWEhzx6vtdoBsfkY5e20eD5w0oon4ym9Nug+3i0PYqpy+7oA6TJ
T0JSkk39KVHpSNTa8e760pEA927sXKuzRB5ZySmkZowekJM2vrvM0ONkwgMu9czPI9XHH0Z+6OqF
d5ounCgRvqTQHExa/J7luS08SDSw63L8VWoJ7S8Uyks7FRYrH/y7NRzLXopW1lKg5zarvptUdRLW
RP0nXRk7+kcPG4Lc7c8x9Da4jPpxAiLecgWzQdROxStZwP91rPpnT9jupR5o0VxUFvig5cPd85yp
uMP6LdH96oqKJ4LYZqvAqtwKMtSum5tgN6dDZxZVs4eAgk/6+VNSNWF3Q9R06PS3aFB9DfIMKrsD
+lHJki8NXu7nTLGOPCRStlUHeH59w30tdmhwfET406oG5/d7kmBHwLQ5SCIBAPfdJsn2tELLbWxA
+o7nCOhy2kpiLxSQrJ9JTcBAp/uShyv97W98JTGZkvFFnAbqh3wEdbXypcsjDSdxP9RYJdM4Kjfq
iOeCtwiScRK/8XPnfxom93rv62INy9qp/njzCwex+3AeWrPBSXUU2KI695Vo57k0fxmstC/ljzkq
AcES48o+UBIRKCKCcgfXADGU5Urzy1ADmGW8YZA5w0PHal5EqJKBO6ZdNH6GhfV0UBc6lTL+qrPb
jbSbAH56JldlcLUcS2aKCY91g3v/4G6avHU1qyjQ96dpYlbXsXNy3LK5sIXOwda8p1bZgxv90OeA
r4JClQ7UknwolU1YyMH8rbAVNzXK+95KTPW+mDg7PRxrTX27wZ0cL/49rDHGVxvZwGQxTEREDRTR
ElVMG0VMTuL2Pxp/V/ivJFM2rNqZmODcvjc3fvkH2q3WtTpuy/4sLCjJBMvC514KnFc/kTkRgfb/
7v4e62WHwgn5STfmsZpJ7w5T1aJhImao/NRDPxmTbR9sU47Q2r6qtTZILu9yqIKY5FCpuPVyiJwq
RUg8QORZLhPCfghlplnUFXu4+VJayYCndVp7E2cbO3Qsa9M1q4waxvto89uQvOvR5SlJ1q1zHRAh
7L37c1pxpi0MCDlWwsQHxKHHhiXDXGOVJUadn3U6XsGkLmwIvQOifgTYD5gOFzt0sao8VmIK1rQT
gBhTW7LchddeJE1XO1N9GcqOObcJhVMQKDDvevEeYimVO4FxxT0KAhqm1EZPS95hXXusoLAEtEO8
C8l+4R9zQUrlLkdc3Z5SrkNMNMIT1HClQasgO+VEYhXXF40sDBB9hbAjeiAPsMF+Oa/+A6A5i1L1
DRovbWiFxHm0XGW2+m6gFR8s6DeiwJT1Z3ClUB7ay1au+W21woOzGCRwzPun9U4HLPvTNsNn6ovf
qD0RsZAgnTAZeVuej4tvnprF6/LpNPyDa3svRruavH0NCdC/kPWFAGRhjXt0W/D9bINfrfH+uW7P
te9mC600CBTVJnZjAAWu8XfiTt4NcvjMv6rwwLdy7fqgY2DUxi8oZX0BWDbgDfoNU10Cj3fI0b2p
GYIXdqeaQnHoWCQN3scVOwB9pmPTUMIQtt6jZeSk+Qb549be5Wih7CdwqtALIKz2saQCjfCgH7YE
mTKWSVyNzklmi9jrLIodkaRuRdBwcGg57YJvV82cddoobxEY6kTiAo/QX4iMVvUJt0fUPBy0MTcL
/A4UIZSnecytyvxGwuoTHlrmbJ5zusQSuQZrVVUkKhpQ7Tzz1qn695Ju9qbr4jQ7AyKp2GRpglOu
+G4Hal0Wz0gH9qjjFtywF1CKsz5W7FGUz6wQa7KTd6rGD5tTgKJ7eku2SeV7oEZYRSUWo6ky5Okt
5DAHvTOwLFjjPzSgNpnPbvm0H2czMIJLVE4j0IKktEXSWqLuhvenU+5lEw3xWoEvHiPk7A9zMW5M
hnmJfGcH4w6WWNVLhb6Q7c5liUFIW05GGS42L6DIGhoTLGKZvIXCmbOXd0HrrcbXhXLCKISX5P4D
tNfhGf2dtF29RttAZh6plpqAAY9a/p7t6D+fuuoYqwaN8p0IYms+UGGp9huupVysuzH78zovIC1/
/MW49JRWU0Gve0DQr3omL2Ujz9jDnpElzp7OwdZuDmOhIfYNY4SKz3BRgTs6++wpi6J4plaZKwJs
LelM+8DUbvZHuG4FXvHMjiDlbqqT3hRVmKx8DMdPOfpFSokIUaYcUU59s4EbLL6+skmUjszi3jH6
bMOvd997xv0VyPUToCPAUSMU0ZlpD4cfVRz3elOY4gDE6N8YL27DdWVJviGnRWrvy/LJV69bBkuV
Zt325reiGtHSIG4C8es2J/ASh6S32EjDi3vimiqU23/E67hncbPuuud2fPjEzO1Dwg4EPFHk82N+
vAN3oAk6M/FzH+Yagvy9keDAliRxZHRRakv8hBA6CclrAOuSPPvTS7sYLWZjTtpREcNVOV+pDloq
bNVDgHjVLpUtjN4ajfuYH5Xg8xmuJ7j5kl0BofWGkYDNJGRRndFkI9C1dnRIi4Z/M36VPUCAa21S
pRBpudLU9jvcE8/8T1fD2F0yxU+o5oSGQmvHkuhg+k67DikYTafxVtNA4Uei9t/6KxZt0kcVs27d
ShtI5HVsW3lCz6YRP/5joimSdeEvy9lTIy5pei1R9897DVDNjJFUZLTeqQY736XcXB3Mmw2FlBhV
AP7sDzI1RpOZBqnDWyc0MR9TIhZEcyA7Z+L/FSq+JC2BSrtAvO2azkuyLIfYsg12zucxkgN05iEn
qV4YnQDjdXD/+ZYiLycA9ukgFajDF+XYka2+sd+SYyhqSdbnFzIAhBj4QwklfjkDg72Wa81o/ygx
lRVCM6rUxWt7BPOBRQnSp05pHSeWEkG1LWx3nG4W0nOZWn+ev1gijf/gKy/ekxvGcItSzsOvoDz7
mf11FM8+spJocUAv7p1tlo3Cb0HsXpAhBXdny+pBSHyjf4Ne2A2c8vQrntMsSYaufPa0I4MVUWew
fP2Adta19YbTD6nJjD2BtB20pu6yx46EmBM7nwBZpW/K9HAawPsBW4LludQ2WZ3YuEj0WVDSSQi7
47KIPBp7AsGfAvi8xl9RvZfFK4nF/BHN1T9CTdNh8U0aXYYKsAvj9rNZlXj1Z9/YKPPpcPjjIeq3
1RGcLtfKigonRX+l8uuqkl9NQRluXzq6kMsPECSDAq0yQ4DKfuJ1E64hmGbAd1KK92RYBiR//hqq
jH827a4qobKqAPNAhlJMrtRpN5whUYt27yv+bzRVLS9XENmHL/qAKBboazUPf+UUI6joSLdQfgqC
qK8vu0gkWJJPwTz5Exh6lF2AwuOEPOCnAINoWx0JoXG4XwwF3j68RkHRiclKOu62JwH0nD8UI06q
1P6RgMt6uNOQH47NkxkuuLKE5mX8rnV6FDj+OOLL9UEqy51CH+VNU385I3+ckFbSZCdO/RZcoB9G
kQxfNxrRLY3Zq9us8+HVLscYzHR8zqWbKy72fjXpXfyFqOGuBqlifg+tQAYzmiuksysFKyUjPAnu
2W7nmmXshGnRwsK7xM41rdnkB2TiYYgHEHb9CDSEXNnildG9RIAruTT+qyAemSzwOKlkT9F/EB/A
/2Ni4IP92YEBHsXI3gKQiWTfXkTWYGNqTsDLlmMgjLNNEv0elVgvP2HlwC6Dx6nWwFHjUlDVZxbH
aza1MAaVbQjJrKMxk2zKGjz6s+pXcNaqOL3Xzsjbo9jtIfMLJMy0km/QI7NJal8haOH6bnq3julp
pBx9x6jlqP9CWRZ6tAXLnzI3FxEiPfXzwt829jWcB5okPsycZhdiCEwS4W+r+ozRKE2bEOVMqifb
UjWhPNMUcNyF55x9umaKFebTuCcCenpqoqd56Lv0weTRMxA69rnT3dXujJ3p7d85GxK4Vp2fI8h/
HeTgsvdNlLwnfixaMKJKh1t9YI81iSljHk+m6+RToTYvxx7XPL1sj2gryDjpdhvWDrmGSCetxj/L
IHHBMF8ZCi0drOTvuxyQdV1MqmvAHnomUbHznmvGzMEx9qnl3NWgsh4qryyuZGPXSWIA2QfC3Dgz
C1VQ4CPEV5Ih/fQyYaIsVL3b8VlqHCHQ9J9Kz9AePrZ4y4ysfu7uSeaXy0HyyPQXtSzlVNTGM5HC
0zVWsZBAmVZbP+DGtwg8qKCTTJn89gp1P5tZFUwpN6yunse5Ob3C9iYj1HhyaMq6/DO0ZXCOwoM9
CS5zHvggoZlo2ejJAZ9/icLMdCfCDYdQ0vigcLvSeax5oxVwy0i5do5zlTx8KpnaxkNqLMcEULeD
fg3uVAYsB/jrQi/Yu/lbdQ7w+83+giTuM1Mlyje5x4ODMjugfgNfnWVXb0AGsy7PDJq61g9s9sxy
KauwsFYhy/UDRLk6JRIsgJZVMsTP3YEwfiUAhM/Mv0GPoSWyXcrYGCp30KxSD3+1rTXBrXhnM290
CmYLgUrQywDTXR990zPXykQJvEcZ9qqCLv3AnVW4uRwKQlA5HG4a6RLq+d7hzXiwwxLPPNFfEl+u
wucD2TKWgZEORHqa3tXExEo6NoVApT/CtrS0FfNzHrLxG8Waa6TuCCAs7zc9mo70b/pq13AUxKI4
h0ymd8jnzQbSYtg5wByEYVZkg95Rbi9m54Lk6DD3BnBHe/0oFutvAkrqzFm6B+nduc0QJViwcsf1
8oZdOlQMVptW67XVh4mPDXSwReExNiKDq/NeN+VrPp+EmU2DdyM9gzEBXo9QnYEmuZ93tbsDIsDe
dGL7mVu+bN9fpkgPMDa4yl9zumMfR5APw0W5orBqQ0XrWMMoCDwiMosxm/tlj5Oe0Z5zC4gprdXX
fuTFgLCG73xUvECz936UYtiZItNlzSHwrXNKWdBXt9u+dfVovFJ9UXGZK94+nDKhLGKTmcTrdt8I
cnkkwiPFgYp6rVZVUEMtjQs9i1kOz+Eo2uk17qWHB+eiwjT5TrNJCP7IKe6Ubr2NoNqp3Bx1AedW
3lswx5V3t5DNe7cmsR3rAJjYNbX0X/qFf7Ixaiwe2lyN9Y8xFO/hCEde7bAF/ReDUagwGbsaB4B1
NCm/7ByzitGVPysLOhPSTNc9qohNF9E+DVlC5ohKcS7nPBlfb2gKsDUyAAFpEPnbK6/DXb8P9ekd
ad4xwZwlh0dkeq53BPIT3ZHJC+tz/aXZbvF+wW3P3m1nXltLvnzuaFQ7+u2mpvZJZUqE9vZis+/K
JnkmOIKI4cVhaad2eHou9bLcLLv4MmXQGrBNUdk5og8J6bEN40wy543c82EI0/kSYCwFB9vbR8+D
8S9A5w89O0o5NN7hNGSuecQ8/KrqMZtZggnxw4pitRjtv2QyLSFiXrgXlsBwfiNsvnmwVXzYjPTW
sOkiot/FZBkvi+9zNr1h+eC+kJ9Pb1hhvFMA0+G3AQaV7P+g00Lk9JkfSCPvnC4o/h0RwFJNsQVS
yiN7E1mvHriQHDOMgoGJBph3GGqCCLISfcbw/u9+FlJc+3oxnrFYeu4fTQjYw8S6MfXmGy0ekh0C
7kiZYKypMZcB84yWkTy5r5aJxDClbPxI99fMkia6Ve2hQLw1rJVMf+/K9TksUxMyfwF2Kwa2lbTc
g8GhQlZqR92TzOf0Bt6kj0cjMXZsWctjuvPi3lgCAxgcdRt0GZkvfN0fYUKSB15Z1TcsHzNGgqR4
bPbXYuqc27iR8UuAUpWt8kANYzeFaNeFSF/NSeR3AYr9GO0AjkaPW3S21Gkjtdcpqp2AamI1ne0V
qaAmG90c/KU9yfXP9IIKTMiwCMTjPp/1Od3Xh+C5QurzCv8Wbt6Rch0CagCXO8PJKv8+GVzdRlHr
fnXVIDsXahmUxYtbyBCnak4A0aFEEH3lF8N0raL3hrsvYgywTccVgUHmiWfXdPsQPig8Zjq4RU1N
5m0aLD2a8s8gmJ6WAVSmojeykk+f9yQ+P/HfJOCUAAf2dWC0xrkbQzRDdZ7mopefWxSm7XKGY1id
vXD/+HF+5cFUyQYLXViVe8s6iElG7oCRgizKDsTQTrTqAPKcFYFaI2JNtok/qvUTqGh7Ca2ZQyrm
YOyQJltJTVgsVAHENCHP02Cnp5qP0PzyPyUSrmO4FUtybiVqSELvhCjQUzJr0Tj/7b2ml7OQAV23
wdxyLpp+J9wOG1F5gx0JuB8XTY2pXijiNc5yUv1SXaMSBezeXcXwj35OWadWx3EMj9nmF5yDT+ba
i6xrCLTdAASGniUmiOjUFCewqIPsER/XxeyJbl+HJZkk7wPkiS3Nyj89RMVo1ysNOpcYZn4TW0N4
FLMtpm5mlVSq6u2DaS7grQK1ZYmk5HBLuEsjXfZ2TW15FFW4g/q1MNZzlut+yTdT+o34ZlawnQEB
5wI1fFFKIAqQO94991o2Q9i4vjoYxJDOiWllcDNDWLi2w/ipo7GnHcrtWAVpFpZ7XnoFm5S9y2be
rcFyuUfgPmwVVTMm8vkaB6gaLzBOvPTgyV9c63XXB+Qm7NwzSjHsX4fOX+GGl5g0xJ6YmrCSiIQX
0+Oz7o5aC5I8CAaEiPsxin4vzITGFVHB2lXSPpvmOfpIKea+NmjHU5eGbrg7y7Wtx8FX5SWv11IU
CHqVpYOuQl1Xtqyh72qHISnE5u+Pk5TWMaEyqfa8mV7Q5GW6HJZwjvMFp8Ngtf6t65dTWnSBdu2k
yDkgUMG6QCzruVRiVnUGmBficmsVhqN+z6RG2zhOM8QaY8PhpL7Yz48mgdWr+iuZOixMsutH5Giv
v35XMABibjMZ8eCAPsLAByqAevR9L1BpD62mKKDOeXwEYdwu/v86qXB+85yfwgfwC3nU+VHhjEuW
7ID0ymQNf5Dv7eyKr1Kgcw5JsXq4VLg9drQ3dA37a9NlL3X0Gml8LjVD3qxRVewQ270U67CTh/n5
SpEavAy9COeSZxlASc7rMhpVXYNRH0GTvMAEx2Cl7W3Y+R/ijFIDx7u7xGTnNXgwsbIdjpgUyo3q
zrYYkrlnzFDzdRpC1U4cp7nnr8CjzGUurTQZ0OUFvtm7aWCRFLX3bngPc/ZMrZ+1Plb0UaaoSb1h
7SaKU45jQHk7xktUh/iBbNsniGCBld9S9WfXopA26S/jL9SVg0gBsaT56QR3J4kD4ZTJKi8WLGYP
pyhqeSJJYL/0CBZv17CcH7fYGhDbBTvr3xZDydPk8zN2xu7RjSGp/A9kwTtGq4cB2yu18aj/aaH9
fEyJ8iKzsjt57R/r7M5TpxnSj1N/7s+JS3u9D91GkTZcDxLlQWVIZF607WYEsOKqsARmHIVLnEzB
PjuBsPkiK3HpiiNBiMznT3wzXVtq/bKqaWlA/H+P06zzJe5NDliWyzGU39d9RQzDK4Y4d5+nikI3
xG2xlmiPlBdpQsjRpV3OAYUb7fWWTseEv8eyDSDldHK4+Tf0th6xW1EvFwy5Syi5hF7TN9xzySTc
jUaF1a8oTPgIDFIwYvrSDplfDdA3OIioB1yEtZzEQtWopgaN+hp+Hbc0e65B08kWq1xdnr1WB/Rm
fx74exLL11O2yQ+JVA+H4hkq/y/ZYHMxVwQFQDozruHmolKaTcwZCMmAPtnbi/EtnV4nl6IgIB2i
uOYG2rK8YJbsQPDBN1s7APS6dcaoYgeyTALeMzoEvEVyiqhoxeDyPp8uZAFAjKiwZPedw8oS1HPE
cACAmewKu2UiSlHk3upes+ss+MOh9wI/bhbMgTPZ0JtTF9o3oFYIAehoe+Xw6ZojLdtNJh5kG79j
4954DfD7CxTliYHXlWWME7Y5F0KsBR5xjIR+Zbu9PXzqr7c2lOSmCn6JGBjouQPY9yS2PkYPiu1w
s18iyMrXlArNKsrvx2vq6PopnALUFWMF+YSwn4tIyinZCarU3bCViBa7FldJZLLP2utsuJuseLI1
bGneEqk4CxqHmu67sRpPB7j2qpHV7QCJOTtx4wJaendS1Umn9j/3MXbhbVqdX4Ffu44W0SysCpXD
SDEIDgKNaGFPKoSYhQKfa/i0PvJgJ0+aHNotW0mloa+eWAXtQkZ4vpAJzcdr29x3rjMPBfHII4g1
0ZL3649qqNoaqoobCqedNF+ES/F08gxBRMcHp0Vpn6Q0E9Y2x62Qs0dBFmiPRc+1RQudL7a5fhte
859lmTPqHw8muxpVEJjv5+ZE4hkao63MFY9WGrwavw55g40bi2H9Lh799zvV139nqDyZ3WybFkFu
N85co9BS83+WKOJY7Dd+ZP6ypto9hhWToYXJWG766D/SrKDAjD0qMv5RLplziw8bHvfp4UZZFCxM
WudpDoTU/zAW886y9ok7MA1ZGEbZ2PS+0Vyu0FarIPfN2QRREpW4Ct3Wb3khqyJw5PWrVKFlzWap
WaLJuA4zcn8WKNb3fEV7XyBxV2Fs786++wQMfs8ku7Ddn1max7v03HLgzdVra8QHBer8eplS456c
ZTApOPWN1F2ZwU/fwHb0pDTPtzHl85+G1Su5wS3COgGRZurFJgo6lsLydvAZNVUmsli161sLYNxl
MeGScuGx4pe9Ip9Al9bsWcidUu+sfzu63/gDt4iCDCmdlMl/ZYfLmyN1P/DljRAhXQIsODpbFqcL
Xr1Tp7/HgmeuxAIJNThJpytvbONt8bR3bOFK6W0Pq+01Lfc7hoYQNB/i9YuucttMFDo1/suZslAA
ebHtwi+WjMMaQ7yrxpkQT0Q4bD0KPQloDYRa8lMzQgUh8IPAVJ7JRzfa7Dyj0NgYKxOtP0YaAHPC
7130JJYCtej3HGnp9bIAzq57GGtb2/u0DRVT1i3XLzcQEcVUdZ2JuQuC5fQAkAouCLLEeoQ6Iukz
MuwswZKOZwjNIkeHZIdjm8NgUzUKO12SanX7HFkvO/uuo+j52HM3y4kqkGGuTLLFs550TzSyVErW
jVCbe6yPFgixGxYnoHAbkmEJl0ubzlJTIMI4wjHFNA8EWKPHsNuTJIzD+A967hT0CNse028IA0/I
fnW5CpV4yvf7fy4XBW3GoIfmsg99sTRuWGbBmSFOkY1le0Y6sPl/to89NPxyQqDbRYVzJ4hb5mEf
f+V6ege0+xcRHSukU9kU6EBFpF9DyVWlBTkmGKiwfhWsmrrOGH6Zc6BVnpbJYDgHKl2BIfhTwSJO
eyUEtzoeTy4goi2Emyow/aSZlB4i23IYrQZjr56BZ5Qsg6U7m4xk7VhiKDJBg8vhR7HahStQYH4Y
yWwcDh5+9muSsVIfBKoR2c3mwPJdTUQQxz5E9n6+29cnR7HlJyJwlecChETPtlN43mXgZ1MRExIY
NrVa4t/3n538bY2zeqSgqIfaxgh5G9HPnhK9MqySqf+eEeiG7RtNNjN2UMu70PXhGhv0NmRH8ecl
YcszOkPMFhI3EEdDp6MLYeilQ+DZbRqf5MFFjpEOIv3ZK/RUlalzKZwHzlG/o0VNB7WCGcuHjBg4
4j2YxqoyGhTntLsereBC4uJSbKPfoxe4VurgBuc5aqXQnvjGFMq5GqKM6pHlTVXCH0OOpISDwNfg
D9lNNvdYI8ORG/e7Iau0HEQ8PW7hDdyKYc3bLQipds5theVs5cpeCVzOovP5T1IieORHlmZkQAwj
iKO7TMV6kLVj7NN4gCOGnA7rP3oWykGNYLH+YAqtUDbkteXuS3fKSSPhFuZHkeS/pclBq9mlanaz
+H3eE42Cd+sK2H2AZdxXSi1rJ48F0VsPKt5vNQlbQoyCR5uy3rQn3pSngr+uEBpq2FW0VNNcKW1W
H7ogdV65Eb4HbcikJLamcjxRdDoR8B594NrHi9TdbntZIC6vUlgSuwm17VWOpLUP7EmijBW4eXyW
lC8L58aERLrSBFptzhWciSl/7FqpvfTa8NkJYaTQ4F38weLKHKgz1NqNoW95pq3CvpFUKp25ACc6
K2exGFAqZG/5J0dzYO/pkYyA0wOz18B8TjfTV+D8yievT351H2aaf4tzOiE8wuRNX2aFU7rgwths
f9bA4XrckjmTi1IQR/MnRDISJMDHLVrYBd67CFuWoJdfdv1/JVufvaAdtwzjz4kmfvrU7rdA9LQs
qQuWm9Vx2+NZ/QvQcqvIXCBWBVeFg6wHG0rp4Ha0bBY57lhGU7TDhOxPuynuIPxl6ysLgVybHu68
OF5nF5QIW69ALxaIlsliHrYMWO+YpORwCHtV7tpt1WRmKJn5+IiF/OmCmJNjrkUJaFzBl2zLXoLj
mz9VrY84sqeQa1CI8iSZaG//INxc6eFP0aUg4MgztZyqUtDjmWb0t6EF7DaODXs2s0/t6rmz8rk3
DArnCpM3i8yOsbqrpd7YNIsYlKl0oGu0dZYtueGcy4IT5xIfvBH0+Xi0jsxxqfFBWZiKojxEqpCT
fJoJ7LPdFNMGvv/9W9aedgsz4e9ijWuPtrke4HKS1SCWiQpzDGTuqjZzFT3QpdpsFfVjkCzOhi3r
9RD3tnbbtOpROnUiRdAJmlm07tr5jg2m2CDxrefajol7AGdI5+G6qDT+7apbBlLMQD0O0yUeCvFm
n1zmG5fiK0ErymanKx4iwNLDtrkmonZb7HtdAIzC48aFWhT6tFnCd5jh2ZZ5V0xV5YQAkTtYyIzj
TcyuD8ctmYecJeKt38CGmyAhOdhVumF1Dc5sLjqHxgNZt8c4KxMysTUH1XIOgsiAygd1UzMw9JPX
dB+vbXDWRfgogI1FngAcpSCzwi/ENPcFnfwUnul94KZI7LAyghysjTmJfvvn3J56Soc908o0/GDl
pTlPO+QbQ05JFRzsUlDpBuy45p2pfIk5VpTt7nziLxs5GeaK0LzSp3gg84Tuqb5FCNdsLFxgFikY
nMq9HOS1iKebG6rDU/MJxYCSfo0VWIxkJgly+lAqWm1JUMS9NFABuccAK36JKImlBjRGHquPhfii
97Chtiq3TNw5YaU/KERwp3MbjmJGmi0YTYtL1kZ32CuXUfBTZqTUIVhb3uXNw1ozEk9lfQKownDD
4wh25XeQ3k0m9OzY+Uu1Q70bwflQIU5W9YMpDHNZNU4T6NqTrPCnnFNqpeN7uwlutMgk1R/ytJ1l
k/pU9KcKumFIpFlT/aI9S5+lAm5xcBxtF8qkCkfrg3b4A0k3tPec+F31xoC2Guyw2kfRKx+2WiPQ
DoQePbIFM/+35j+B2TJ6JjR2d+4h2NcWayMuowso34koulgWkpRdZQPq6q15q5dHBr1yK020JX9I
dLCUxrlOJdGT9Xyh3ZaaXZs7sKfVUE0qwJriAHG1lSJvc4X7TWsRbBdUVa2LPWT0b9HxJhbnR/nq
ic7amqUdqplJZ73AX340QJgZFpgNbN7I/gMeU/1oISQlNzmLvGB1yJbMRgx0N7oZ86B6Pf2owZwW
mTWrA1PryQ3cI1K6ezYsG58YKJdpganRLMGFcYBONdCpU+aneT/ojZX0N8EEHfTVZAvY0appf7Fv
HYzfzhxcTfL+nCUHHB/lt5W619YuYj5oCslkAt6H0uuE8BMyQBtC09BDWWBgHUcysUeYV3LGlSwR
162mQOSKuF7Nqs7hbNFLT4EnUFH4Aj2Uic8/qGvw3StoPrZjs27kULIHNyo8x5UoZs8gXRVKBgnF
nLcVyrWOljPJVRXQ7saP7ocY4zpHOSd8083nwk2MGU1HAzpibS0jsRJAFsyuUMY2huFfyVaw7jTx
r0j5l7/Lh9NlbzGSEonL+J3COLlP2X5Bm0TOXMZfWdhdGukepvAsQ3nrIUo/pGl2CPf0mpHjb/5Z
v3p2BvhfIy5OlrYy+X1Fi+dNJr5G3VyP5Fr31fgMKWGVFvvulT9IHXe++jLtlTEVajowuFtx+q3s
GAtbuWSDLuVcJRNvvZBqxzJrAFiIO9VGhUNlrdbW+fo0PL5bBDS6fpT+Qu4wjZp4zRLke9WWPhKt
DuiO4mhsB8m7swPc781XVG3R1ld7LSqAzDLmb7d25FlL/480vj5cgDMyeB3j3UVv0gWH11nS5BBM
veSCUMmONBtFUl4pGJydlWhyncs0sDaV/I3nLuMjO4XzHepLevEP2ZNp7h21ecSzL9V5ijqS1dal
NvkFhgwC3KuM4fzq+T0y/dH66uY50nMEqKz3uAPgraMnPKKkjUD7+4QLCwi+9BhtDKU98zY2ttJJ
vnUnDn9TvL/+64ISa/wV3vhJGG8GDYXYxzF1YJX37THlkUB3i+VxgmKeIuI5W2IEp+VrMoxPU6KI
wj/P9cqP+PrtwcF1wrwzI7aNO7NWu7MIzntLTdEgyymn6Tn6090mVAteMoRv8St7ehm1dMEQtS0G
6jqH1zeD1QU22ntaT+9iA3dReFe6qnYPDYVd6iRccU7g6MwfAgAgGPEZw3eZ7PAne83k3HOevRIx
YE2jC2j2XjSL0RtV8QuENxvUQLxmUYzZLM6QZMcK7vraiNR+1cvCNJ19s0ovpeAD4G3etFdpeCuJ
8YKnmbanpGd2cHoLwwyLxg1yLkkUtLbk49tDKnmlsiFgd/IjJ1LkfgGfT0JcACpb5rf7APNiBY6n
jzA/pI4QxEwFVClech9fq6c4xPSXrZd5R7sVxhSapElHOMGhU1vPtxk2jREiNNmOrucG6qRmfQTm
OiYEOApOKqRfbqGIfZBMwggaIhiLolN4WYie/g2bRkknwAe6ilckCNCD7rfgqPOahacFpQ9rXU2v
d2esUwSv0E3rEv1OJPtwfput3xBTiIVizklsA7DfDV+pzGF4h9xacYP1Vsjvsg5sTIWju8vC28gv
A7HlJM9tWLotYONRSb6UUxSev61ep62mJ8kK24aDiBNuvNwAdBm/bixo0Bukxa7E+2ehDFLIBWPK
ugLi7+m5d4cw9mwyhoiXxA188OBTtFZi+wtG2J1WsiDA2pgnpy+jmd460Naco7VFFgTtwoXHbxVn
Ii4Ff6i0NK3NjGL0ezpPaNmcIBYCX4J741j8LSYoItOr7JvqDjqqG5Lzn64cyaKqjWXXvE9Uuaqy
4MvH79b/JiHoL5hCmiVcwjz9z18pYS5Nl2Z+z3cUiIETVK8NCU+0J2Lp/e4fBjj3VRjkHaZru2RU
Li9++RfGwtg/Z4tuib/p3/DEYY+J/tG1ytb3I1kObbVkFgzFfWsAVbA0Vod5Jp39xssblgX5fA1p
3kAl4voIKq9CCXASvBjlnI0y5HlP0U+g6Tg6AoEirKMRj0gIx1twcsx+p2/pwkyh4mHNWlaw3nhS
WwLi3mqPGz+A6Mt1YAbs0wyp8nbbTRwzQsf3mnutwJANo65LkeuyJoZkKojjFo/ppQJEr+e9lfhG
cxxZHmzoImMPdc3b0z+v6DxSTXUuvpGgBuq0aNMX71IH+6IgyJIKPLQ97uXoImkRmaSSuLOdKjY5
IphUBdy0oTKQ4TsiXlPayNOoEQz2KHQ9eoCcdLZFiblVfTdT5AqW8Uz59do+A7fHzMYwkHXXkypl
7yGTg/LJTfpjAFqOG7V2QeE1oSywaEAiZszgmrfvW+PzHhOBQJvqaSKoEjhIrhiRlKsi9bWVrQOL
QbMYUxF3uUwNS8Xs4oW13K3XR79Ilk5QXsNhsfopmsg3ft0+ByvTWsg5N4SQYv06ru//V9/96pMZ
xhaNGlVmayai8l31Avj1CH+/hk+OiDsMZvcCKQr6wiW9I1OGzN6JFIHEISKobtwaaBhQkZdahLoa
pU8F1fX8HoivaZ4Mij5SnfQQEriUUXEgWMiREwZ/jIP47AJzdqhWfTcyL55LE7O48MkHCxeDnbwa
CD5NW/TAQ1+BxucL41df/OUA9UhL0VMGzYMRbei+KBEHYmf7wQDJQQB4O8dA8rxetN4gsMi8kvpo
grrR3Se4moLrkvHRWuY2MiWgQNSUZE5W+6g2w93hPj4PGK6NoXQGeFAlz8zIZCXvlm5Yo1p0Xcwa
iIcJ/muuWWXUjlbviNBK6rMDOnUkRjZEYo8zJm2+AyeyGkTziCeE0x/oFGfxWS428K8wNnam6Qz6
vwhwFAngnrtJVRGWBFarj8Sr4wv9P8AO8tulLSsJTO6eJtFRLKR6ySLjMAClRsXPc4Hi/pOVMHuf
2SUQ4oxn3tXvMW/kCz+tuhYv57h7oxTMiz5TqouURz7KVH6jmxUxhXciRvXa7xiWQlIsy9g6xdkj
vW74z2z4wwJIT32JT0E48c1Zj06hbgMWy9MR9n76PeGZFzLXlnJ2yA3/sS/ocK49tzTRVHHUKNP7
E+U65XUFlxfTeb0P2FyC+KxTIh1zua6+CPxpz0jfKEUw6KUG17jqqZNZ+yIbZSi+jfXF1350ljAK
+v1pa34cBX1B0Brw+jGg0ZBuznYnEO+m4VP28VqP0je/J/M8vItUBnjECFyjvWEDbG/agWOjL+0r
MflFUqR1tvIbVxmhlZqvYAjCjCEXNTmY03qoWSY/EJyih/KLWSvMzPpxqzqhkzRolZXjzAw5nWrI
b/ub8E4AGBgoeqVE4/J5Ltj21enAnLb29j4stQHHk5a1Bmm71XwhSwoxZsX8mGPp3JL5k9iQdXL/
cLHKF5A7p4Bv3p2N2ixa//iRhntBgbjXk4dry9xZRTUEbftib5ONBS9oMsC3af4OH7MRcyGw0Ncu
sWweJLqHGMrPas/huMNFRbF8R2UG7ioNOJuhUZtguGIj8vHCrvxkzMs/+wrYRBmMYln437oOuXv6
xtodT4HCIOiuUJQPqpuJDbTLMQ3LEZqcFkghgrn9lk5bbsEFL+76NKcvqKo39v0NlICyO6XiEtV1
lKfBIviEhE+mIQ4kE+L6UnVuHiUmX6fZyoYfCblvtxGQM7HDR+SqjyegtdyK08zeUbEvsg1hpEA/
nU7h12EXm4kShCHYWLtx8JjkJYP/fkGRgsDQFYDjvIw5wZb8wnzc3jU3TDCCFWN+Enk0NI1PaDQH
qNGrzpquiOYk31YsA6ZXUjbExQqs9HWGuvd79Jtd7yYd5QLUCOjEF0bGjFBHoSvfDeZuOnvnAQYJ
lZO/gz0A631R5USi8phv86Guc2C8zrMnzudu7LAe28z2tkatVFSB1ikpACWUzzXeg0WxBG3IHnIC
Whd4+1Cyqvzlcpp9e1DN6ebpbHUSKb9CrZK6OitfaQiUOWrQA6poC76bu0NXwP0s7BRw+ncikoLP
mNtvbheYqzXEpSi2e4qHToQHAEc1z5CzHlP7t2bk/IDVYQquVaVqnr+x7Bh2UShETMBPrlZjSKoD
MTFL0XAQsaa5iVPma8Tzq9WrVx9KOCLvdbYMMp0uk04SPyWOEmEOqWpo6ZQ+FN4KoGJKY/Y5bHDZ
CnkN3bid8iiQJkY1kkYwRmTVKL5rfdxMyEb9R9Zu/29NfvF5ryk2vesEbVTVyEdp+kYi28yFn9Bb
zenAU3MIIxiL7wrqOV9QYUXdrnhHTx9S8QzXRQffiGB5lwRNNgxb4bG5kUa9vyUhDmGpj0tL9zC7
VHTlAI74fAOtHXSsd5mMtv36/jqmicutfJA3/CSfTTcSaIx3eNq51w0fkRccPTOCUPNGTYbR81Hb
1n2OYnw+DcJkVP9RS1dclX+kMJgQxsy5zzlNrOabPxq2JXbtrqVGWN68/dJcEKgsNM0SJjJYBGTd
A1+LbBjDaO+97C0WuxvXRCGupB78n6CJCSZY3x+2wsp1ciK+R1DWHTkUInD/OvV0Hvm8FM9LBADz
9W/VecNuchygumJPJ6U7lbDx3d+obml3Dxvy5QmwqY0vHjGlw0AN8vl0YvShymZiyGGGRmbgmcy5
+2YAFMYmj+pzzImN1DtiWG080WQRR7En8m9ClVb4YbGJkpmHmxR9B0to6iMFEtWb4dL/V9GQjFgv
iJR1FkAYPmunrY/v3hHwJrbQiLmbdnPSoPMYohKXeNYufxV+i8rtry54gNnTXk2+/VmwHBqZ47WZ
SGRatiWJ/NZGfcoGupcSinUah/w6UVugIEJrz/hEvJaARw065Z/KyoPQ8/ZavLp8TrbD8kDxExlH
s2kxoKQqDT9+J2J09eGQcm0mgbdlLJeDsmuxeg0n3Bhm0xasGOyFJglLmWq29atJwp+6yoOA+GKT
0YJ/3OS+w9F5Txg+ZGhoMRsAy55LS+pEzSJS9d4DJ2/DMh9dYAYNn0l5HPYKwQopdZEQ8Pr2WKIH
TI+ppOSIDKgtcVsbRQKf63/BBfHOWfl8r80vHQJjTj1XPWp42clT6u1dQoMomZoaa3xoUx1i3oZF
ilokqI2jjcI0VDp6b7YP6JslQrbfFtu4K/X5+JHIm3q4rnaAYTlgodugivZSLjE8lLR5/clo6bsR
vePIafTkAT+eAByCVLsQjU+S7/xDaO16tya2gEDlkMOlf+auuVwaQ6Ym49JHMIHyQ5Fhs7bdjD1H
zkya0LYhDbdrpClRQ7vP8xqGCne+VwUgSbpmcF4NsRg1VJWIIO4pxFMzyuTI22vIQ2cskYpsgeYP
ec5WiGX9Hg5LvJZJCFEwDvsUlMgSNh1WFyB4WsKQDklSj2xCDuIk6lnMb33tLftuEHDebsvCM2Un
GPZ9PlEHNQjRm4UzTrbu0tV/7jenFyidxlhFuDrOZmdMtsVkbpavl3SgilZ2F+U4GTtzgFP9e4vQ
/ECWbXHJkFHe6MIZHiJUzVtvmG/CnpsKXYhj+nPhNwJm/CE61K5/hJliWFmO1zFUwpDXPcVGMmUe
2jPydBtsp9kH4upovJ2hrjKNXB8Wtpd8IU8uf6ZxKB9VO1LftzfU/sxm54LoHYdfMOvut+pWiH50
XZUJ4HyMtnLjm5G2Ci/FvfI5jU18AYMcCZ8LHOiV+JDpPygC4SS7auF0Qc+EJFMcK0VePyIXf1SM
BjP2/i/wBhlYoMG9RH0bKvoTUhBou3el6c1O75dnMkL0rG0d6cCY0ToQY56NBnbYuy9+45nbpHOL
2RWM/1b37BprgKh4+pMzokq02hIHYhjjQHPGWUy+80Tpk1dlN4XIHRQ8yCoPT7/Ow63YkeuZokpL
WiQwXed6C6eVZtJ3P7OvdXcgIofzHiAe5548LV3sa6kfoLyfEKM8XDgPSt/JvU86jLDHUdBG2QAY
X2NqJtbEWgcbWu4ZiT+FtF6EaRh/je/KN9xuwDuKOycPw17il03dIheMgomnrS2skyZ0T0N8hLG/
F8RqrUn2j4MKz7EuJvVR7afDjkEU1LvMI9RFhWbUk6mrbA997ZuLBOiWSSlzRm2PcR2JYOfyS85D
T+m1TIhzLetw1r2ACcnmGJ2wo2CzVWp3eyascDx4u7Cn80/Cw09ji4ahpT+JRm2x6E0/tkJCxXPZ
cBcpnAc+OOlboSxS6UyTFJ8hW1kHDXVYrgSsK0eErFfdXgDd9KAVio7BpDh5fZCnygXVK2H1RYlw
dCNAER3rx2d1UhKi6fFHof+oXyYRR4K9JX6vNRcN4yK74+LQGYAz71Bi/flhzh/fKOxBP40N6Ski
+6IviwvxBG07hjrgx0qyJ9OT/RdCN4hNLrnbWEjX6ZuF2rwKRVYJ83e0RyPl5khzhpOpfq+nnF1O
YowCcPLIQFT3IqowkS7f8h59knXNuvYu6cPDTu/mgULi/b5aKipvOwohoXIkr6ttRJUxqeAYov7M
++/DpJdPSBkRR1T30nTmxOxwprbP6ehg7d1aK4op93phK20wuXk5CA2ijKSl/vPK9GcKCYbqaBq/
CODguRj6ZtuB+7mmme/EO8YieHWBaCEzwDs7fkPEzcXH1dmonYbCiAJpWIUd8KkJuOtbVLJgTLzg
BPgwXC8S64mDPYugXtPLK/cHxjGXh9h2HCoUKtorlk6ylbozB/lCQjSst1i+u5irIa+KchTxh4T0
zFjt+AfBVN4aG+S+LG8UAgfWLFb2QqSFNsyo41pG0qUmmlUhSGnPVVwYsE8/Qio/yWhzKrQlEThh
dMtskItmiUB4oRPGEoBnpHNTPf0aZsHKITBGHXdlOpvKwZtY8LFIOR1R6k54rejVGTZtVvrQi8/v
VdMAmSudKoCQ6eWFMspvLZiC8S6p/n7inVNOfFYvK7aLqXk6qIjfDq1CychxWR3kT9FbZJxiWBDH
/4v0rYTh5CCQt2MP8sJAAqsAI/gkaMx4OHt/DktRfTnsLs2u0mZ6A4YAX2BvlNkwsMiXRdNctB3K
hfusWZVwHPRLpJKgIT+09g7pI/jN5RLnVCaeZ519CetVPxqjmrSHi93DietZ3I0WNXjfitaEWmEP
CfVBAqf6LP/73FB63kSDm4IFIKTZ2bfbOT0x0kPswoeUCHuR34c7pJGcOtjbfmb5OXEL1ssq8pg2
d0bObbzFiPmq5uNwK9+4mg4fghphznJM9/q4acDpyuJoNx+g3iy/eITsguqmZvVzjVj0o17wxFDW
Tjq2tWa7TlTwoJsOSSYF1949yARi6t57bB+gIMBmO8RHpUYhlPxaHxNqAp50s415mftsWq7rVa0S
JT4wMKb0LKK6pqR2Asj53FmmqlEL83GPujf41y9q7qZYL0QEQwEeKt9GYC0DFAezvd1asIIOXiCY
ecw/VEfdgxNIPYiAdY37JyCty+FwaBGFcgCPWZw2EgX1gmLVWlnL22Y7fVohUD/yb178fJnQF1AP
bFVPm4k+SVzRGHrYI/sVgfZbeccw7myZL9aZFfu6Cgpab0YuJ/ZPZXf+6f1VifiB3pTYIR4NVPaf
hP/Y2jbuNo+z7lxQioecncK4nuHhoBFq49wvF5Ringd+K5VrDP3tGaPAWrUGyDRXDvSbyV3V8iXH
uKa5QQeVdMW92T17rznuB88L72/5xZQgrOUqIyrL9ziGE9VBicjwOfCwJOtOoCnNQd86i60F2At1
ug8pd4tnCCxt77gkVIzLbEV/TYEkBir4X4XepqS/fXtz2zyi8WNxAEg6ovMMdMCMAVLJv/MYGzlC
sEW15ijMatfPZTDkmgXNAz2FBvLQICWb6hs2WrjGLbYSzSWZ/rQS9TkKt6aKW7aX5eYOlVHhQK/q
/7oQlB/OUEueOQO7hYevulO750VkiOM+knDVxqs8EZM3V1KeT+N/2Yh/TZOI8s5Cw3nBjmsX90J2
zVA5ZxrmSCAK2RoUjFyUa7fHi5XW40fF3bVma9Tb+/xgRgYqfVX01Q3vFSRf9vLlpbTCD28GAXZE
rSdeuyZ1UDgBaSOBMTbZHkvWwt6wm8YAW3xKHJDLRw9Y0o7SouP7svsZQU7hCvMxOgQmx2BizcYX
9gnsjnA8nC0ax8pMOD3Px6cweEbskF5E479eDX8EBOU2VV63OBZs2sNT+04FXUKDjRqErX9WEkGb
lX2wAf6anfbuV96gkBcJ7PDj5icDuLe1AXD5MpZyW0wXMzP57VdGp60Tkk7LnXa/zOY5taEHAURv
cmofqEWnAJMk6Pwl+HpU+yBXlgVeYbTuhzfSeyM7Z3PgQNM+FV8JbnBaLVM71MJxBcX1oPBGbX3M
daYv3cojhPc6cNxf2dguXHxauHd78GxOjhkfDsN0fnI+4zMDZadn9lnKHiaZNucti8hMIBYEON2G
rjRc5InIgjj1Gl+eVPGhyPKDtTcQIijSdVkfPL32fNFgW26JRS6qd/f6FJ1XGJOV+9BRHe2YnPpw
S4y3K7HkHCn/I2z3tt0R3aTV1tL6rpqsNTJJRWIFXFA68ay60q8VvXJouPJFlwvN/4XZV4cJb3uC
xwOniPP3XISr2L6cAzdKAyPNKC9POKqUZor+A3rpqeVlWuxNvu5HzxH/MRs91d3sUvkgIl+xJ9/3
5sYmiRi6riHJTkIbcAZYfKJjtketDRMqQA+rAEZ8EDWzjjWZa1A/m+/PPHaSY/w2XFLRZ5zazrZK
fmwg9DHH37a3bIR/0djbJF0adxgE0eIYbeACA/ZSAakVs+m6Dyrw+oA+dfPYXMA5F4nXbepOCNZ6
kmFQn6at5AkZ1whbRFAAaX9Y5eC4yWbcI/jemuVI1Jg0J9GxGdiARDN3qY5tKHSAmBajWcCkZMS/
yAFFIbSurMFBIYl/MSZwtPphC1zeCQtgJUsMlTr45ntBwNpCvgRJv7xTmE8UUwKj6pbxAaWzVql7
LXBR2fUtiajrNX3FG63rzdmdfpTTMW+YD1dlsyMU3gr20sHKYC+jJZAaoZFpz76gVPwGem0DK6kY
YRZ1R2l/1bQiLcJqUHTivQpN1R6dRVYNfdziB1vHnnmQ+w7euTQJHBQ0WnGVGSetVUt6PNSB+Eai
GP3XlB1AYkCRlXCoDyMTmSB5trWVybm5ChmA3miou/CflfnZzrEK/zk5/B9lLJbdFa47cEvz26u3
DGbf2W6yHm0Y9tgfKDoF3t8tnKpAygAsthCG1dlZaOunc5Ra+8WgmIzNXN9KBxISEuMZRD/1d/hc
ivCowRPLg3zOeSy9Twxp2Yzoc0Qx8kYWgpIpgDvC7Fs2+BYwxwzimUeC9G6xKNYYjVusEmV/wOmK
GwuA63KDgy0wSBOs/WbFfW803P52b1G1Ko/wHlLFiK5+a2Gsp+o5FZfT9RwjTptq8tro55Mdox2V
kI6idEd9VsZDHhB+mjnCnilbg37dYtqOzbXRdIdxaDG2BWBjuBa1WC/wjFJWggU/twEJJ8LVzL5X
xBh9TZTYL9FxLc3yA+FQqK/WfLGSCEWxAMh3ORlQpzmoVP3NnTrBHGuybLw19xwGEZRD2MDMB6qJ
tItt6K1/xwIguBM76p3RHE/sebD2wn2a4GyHuIR6LYMgI3SP0SQJ/O4tGtPbZKnuPY9K7jkZunmr
I8VU0EF1LQJPhjmwlM8Ih+s9EAZQYjenhM91JRPZ1b0OnOAL0z3dzJvRRRRT4d83ysTkYjqgsvx6
CHgXT9fUiQNnHYFJdAVuQjaCBJ1ccmiz20tF5FR/CVao5uCY9a/C3Md3c/P3NTZU8E2mAOZk+jc9
qUhULdInWhZbw48SwkANk0avXfk5eCziy4hKJnwzodtVpPa7WOl5Rdm8TlYi1XrRaldkZEu9o25S
8+DFWYw0GuXnkkelc83oWSM5naai3WFc4JMC5XeLE+N3lD5sW9rG2+6fhSKf8Y2MSRyw7yycISMn
FzUxh4kyQ8lZ1EgtlcoUGkcQ2KnNU4qXHWmYxpxKFrPZhCCcEXVdYt4MFjvT+JIP8FiaAcg4BkZk
6P6QJnQVdb3oKUwx1IBSebxT95A1x4bYgBefbneZSUDoeLSdlI5HGYjXGvVTcXvcWxBdq1MwKiZV
2l9ikV2CoRMcsXuc3nq0pS/O1+tHX1vVqkCdhmHC+zlA5M7peQhl1n9OiL4+CL2aco0+0KQedYcz
tCvTVODuegysWvnXCaBGy0GI7YLpTTekEgxkQ8c0pCTkzDSLOG7C5LrQh+Urddobh0vJ+gmlQl05
6iiBrghHxSPHkxjBSlimZEu/RJnYaprNNW+PSjeAfYdLkgpp8/J1yY0ScORIL3E3ixQ1DeffV2IY
P0BenHcztfYHxLxocR6dMihCvoR96aCPbOEhBDQsCMrlF0xS+7jroJ3/kVasKhsNcTzj1giq1IK0
2zwFJ2PuvZBP3Iqgfdfyt4P56qIgkFroZBO/DTvSkTQiNgBXuIBoKdHnb5zzCLKkxiUPer4gySlv
iUXWGrOyqjs0JyViYnRalvxcMJ6ThyWcrProTiryFoQvhqenTi1DYLLVVFnzkbf+N14rRsxjilgV
JBfcbNgmANtTndzCmWC042zlL3eWLcS10GUtbDit7z9z2R+SoeB22B9z8AwYK7u8aMexNRktBa9l
7ygUmQCHjHmcqZ7fJqK7u3sBYt99JscxCWMtPLyaC0//s7Cff29j8nJOHL3epQHjR8pH/YJOTYX2
kSwWxiehWBdVi5nEzErGYR2auUkQJQhC5LWZVkDQ6th1wOyR2TMNAM3/H90mbpygf5p/lJEovecf
XLNw1mhghbIayaIg956EP8vv6WnOPMBmghXtc8bCyTHjN1sJj3Sjpx7Ah9jyG8VRtRElfQjjamWV
Xcj1B+RT7fkMexSUOz3hwM/jyJU2CLRTH3WBGChKm4Q4pAtNiGwmxe9H7wAugwAXgGEx0cK6SFvI
JxEWqiWhW9X1F+TQsBmJ3bHF0kTgZBc20yza7hXGFF8FGzFssdarw3HZYY0ANqYQdxgSbz6hZ4n3
+X9IinNCZwYkOh2qXhQL7u8y1lvMB3S1XaHaJGFBxyICEoUPgDHiYX/w+HTqmNmMtcSFEs6TI1BJ
+5IX23qFcu9naGd6rRsUBHX+qYZ722NzpLYuZjMsTX+ZbgSN+y/kreffEodFnMykX5/4Yf+MDgT2
+Yo4Ygvqzt1l7VNfeDKOddcpZstvNjElen3hlRoa2S467cTIc4DZejfD2nIgAVvbhE0QpZ4I3qc+
Gu6ns0Ftt6p2RDZBJdZfp80xibIyR4dVI2/ZeAdp7/0feK9luRtQ9Y5+gw1UizCo+9/UPgjUIt0p
bxuMSvDSFL1RRpjbdnFt7iDxAY0loQqV54qtIyadUFc076z8mPirgXgTYAgOprWmnHVNQ1jsPZjM
Oew6T3jssKHa28/1zDSl9nJVJCv/hu3F736XOO9/8cKUOeSPzv/K5xJLPwMwXPqGGIlY+BqNRHOV
x6Yovw8bJMox6ZOKAXyhUy5e4jdcz0hek84ZX4YmleTrZli+Y5LshfBypHiZN0Z8wjDGfpFJAdY2
iBf1KAcyox3m2Yw3cxd/omUJTvJeIpNFvk4RjBRO7H1LKxghmEjkQ3KKEZdzOEb5vzZrnjketJ+Y
xSE7VoZ+zI6lM3hxkjk7MT80SyK6/krssgrAcInbHQXvJYZEV5oFPF9FUInqzvmO3c0aol64rC2j
IDP7fzeX4aidtT9xLVa5E8kobzdpj77zxjrPa0WbsmYpV1+DU3wY08hm6dBeaC+q2HOAyGEBNQjU
wlMHTdXZJqvIr3k+bPVqyvpmZStjNyK2eFbJ91Ko+fA0+sQkDYZ/hn1V8VnlorRvYjl5grryHiJk
qvkwUzo94mcdDMTMambm7/IGMhILoNxsD3g8qLZdeAoeKi7vYjfiYuqDNITgGYy11GI8uHUBI7Fb
2uEIhQPigupGeihzdcrpJbvgpzH5TfCQXbC7X5+h6llT2E57+hL/yUgt2PZTV01agpvyVcujoMik
VxJEDW8/6iTZ1fupqzhRk7yTty2mDofDFOAP4kmnD/UqEHaydCM8SWyIawd+XX1QIxaVmXJ4WKtE
66Vap0Mh029YZ5BSYFHqFmWKqnOkC453Pc4tKmxG0ggT23K/MUpQTDCB32M67PID5pRplxcIsvKq
+KN4ULDMsOwLsuPj30U/o0LxQA8bO3PCKt1NZgEq0mjHMCxWkOTbSr9/HRdGBYCnhyS2Z6wpD0LF
xNAiUCX6mLkQZ2TojCS6UkAnqe48l2cOINr48Zrxb2gFstxxqE9ufjSSjgTm1JtFbKVcy0UiCCXU
S3Aw1u9Hh1S76Xf+/SL5NF74HvrkZJPEwzs9RjyNMiHc2MfQKKj8iCG8VXCeco8HMtKRwWqxGVC7
R8Jpj8TTdkbLz1nV7aUNz1NzN/l688crH2h4fhvTjBbsQdBmpS1PiW5GL5ipC3ObQuB11VwHZEAk
qo0N3QP5xIksTkqdHXfD/NsHVucrY+VpNUvT5NsPBS6ybCArguX5ZEhHlh7s7zth+qq6AW25jM40
bwkZjhwgP+hHO5DRYx7dUbz5uaUAmEBMQ9TqXOelo0WeN3p1lX6DZBGSSIZOkg1WleFf98eVU6+q
B3QaoQRL6Rg0F+fcNqFwFb737pbMkxTtnA7mV512cNMWMnjQx/9sER8vl/0g03ZGevoejaV9CB+s
54/RTRmS4mVQCMywrQKXi+QwBGjMnYRR/IYQM3B3Ns5kPZz8Ct5rOxU2MERsI+FKQ/jhoXNjnNXG
OI3tDdjGrtcrKWmXfSNn2UuktEEInJV7u5FRIAAHNXC7cfNfNbwlll5ulYku1+Xol5/B8kLGlceO
JaF1wK82vTvtBOGfBnShvz9WE013MPFN8W8L6EIWrRkpEWmKB2fSY0VCyZ+pZU6Txo3JbplTLiPT
cQe1bDOpjozLYMb9cO41F9czOQDHuOlR0IpM5gQ2aI6jNukwraOcNN8ImI0v1qRwS6NFKb+voPjg
UXoCMP4P4VJmQMx1Wo/fMB+STYrKRPrXQqCLm2o2JQCQmwv5jxoNS8s5+x09xKtN0BHI0QXGhnnR
FFgVDQ/5cI/MNsjHJBX5SXjyMj70+MSUaD2rsUvgVLZmYQgX0uTE6B2AcgvBRyMBRq8kKEMP+p0o
uPykpybI9MkzFmTKTdxWBlRozN+u4tsSDPkMg4Cn6qbVObVaPZD1MjTUqdLbfSmt4w/emefoSYj8
7k6H7aJ7TQKse21UpHhxSjH2WOmQNk9ElQruRjay08LzU2HJAZAKfagTqYr9WfVdNLFizyPa3no3
2Iyp92Q5ejeSnsM5x/pI54/q6qaOSyLSUS4p7vAhYdJypzb1laYqroiHXNTAjJbcAdliGOXAM2/x
BrgMqQsHxV/duYyNZ3yo9tJXJ9SRA78CFX2uzTDCDalzV5bL1LCjLP6P87f/sJTwfIgSWWSKMCl1
vOg3jVUU24y9ceS+kHJFePJUyMhlejC9uv0ngcu21maiGby0YX+5xsZkvGrirs+xUyx0ozxQGWYu
1tNIBxLKNNxeErnNGNNIfpo2V7+zTPKZNwKrs2wIibIlfLWijPWwrqZLr6tIedVKt/LTYxI1qHmS
OiBTDFLqYe0CxF2UKp1CbLDyhmKKwkx/FUAqSVkDYD0tApV7TH8WHhleKPqgTIRt0miuH+JlSTVY
I7AzAH+HMKh6woCK9yuY8wt2ut5UBjy8tPhap/MI80ZvCGMYHl7jT7zdPLmHTdHvtZMuqIr+Ftbp
5G4ABFqgXWYxzP1SqbiGjg3wTd2b8ZAthdF/fTNS2PMex8WtrDxDbS9v4fFc5A0z7fnf4nuuv9gh
9S7DMwZ3n0xTNEf+nMsWtlyY7vp+R4g+xLTJlu9YaeoWvQ7v7M7TivEBo+VF2ebo+AEn7R+oidSY
alS4EcUKaXJcyMfA8n/9Je1Jch2IwGyWWixaNR39x21BjKrAjWSWcs6szg0E8mhSWNiSC//Rycpm
Yu+/UcuYK0XowZDxv6f8gyWRrm4C8jNI3BYQXkMxUskXQt+JFlumnEUhTM2R68JhpVtB2yk/XFRd
+uCLZaxC3n/dbsOViqsCeKoMT3AElQz+rApLpFwM8meZaI5CWpC+KL8x9xFr5LKKGXd0uBqI1Qrk
YJn7QXzYlhec763T5ox9xXxQzqm/558/d+5jjadWtT1rfgYpyxKR8LTseTiqMYEff2MwQNzN8WlY
Gm3+Q3nu10pEoQqRwOrt9Ycoq+9yw6Xza0ao76Wrf/HPjjCVDcB95JAP/wy6jREBAkKVTUr069P7
LMaNGt267mqW026suXUifujjjw4ryt8QLw9cbGF5ipWAz0EIikK3lQkxx+83cncqFVpdiofo13I7
YUuwo7ZDccE8h0uZ0zdYjX/B4Y9G0mx4H7YtH5ZLr+YFvPFrswyW78M2GGivcZnG/hcl2yFGpUEj
U81Af3uK24rypf2u8oAKDJniZlg3stxBOeIiu3b9jskE6JtOuixXVDAUKYheMedXNBzQoLgL/EMK
Pnl/JlJ/JwG+1CrJW9PQ0GIdD4+WGiicxl+xFBdOvAbCJdXLp+a2bDwgoBI4lkdGdxHra/8H9Pbf
EpQTDg2ynAIwtItEV0pmMK2ke14iRTyB1v+ArhiBXropca9kFaOzPtw6PUXVyhS2pjcWAq2LRT7T
+jpjSkhpjwkyr+Rv6ja6yPDfftY4qd+dmVuTJz3VCq66o868VKg/9isdls0P0kzHSb2DNLV3kcoy
MecKK1TUoKd/CCATvRgtxBOD9mq2/KSPEdYQAfadhpLgOmfvHxMrKniUMNyKlhFB4zhhmz02oOyD
va+tWGcBXrv/4nCWCvzcWIpgARBMeL7+2M7iQcDmp1ap4lu6dRjodI9oU8sASuHZ1Gf7oCCw7xI9
5Vz+0FJGb3AohU1fXu4tpuTdLlJCot8PajsmRi2K52mlsPxjmieCKat1xnHcqoy3H/jGejUwmjeg
TVtDLPipQj0vmuEd0AgAI5h51+IzDrphwHsMlrDXL1Q+V00FAJ2BLRDqhfmVgtRRoR60XBnfCyej
KqDLd4gi+yH7C++REPnxZARLnqGlwRo7zntXjNsFj8BTjnQYV/ul5s+dRRdkmNlu8d+33fAHdjx4
AqgCgHAT7WDjkeG/rzH5marIXPzmKKCerm6PFI4JHTU/QgvwXGfdCoMHgFMcpHDpTrDNlDp+iNkz
mfqcE1V62f4SP2eIKcBmybuJ32p5p5hsSSLprnxSAtZKvMzTAdMAlVhPN1vKD3aF4YUYzMMY5X2T
VlZDi0EfkBspzC6DldgtmCUrEed9I0J4aX8AGtIv5oewq7FsrJMbCBsPzVfiYePS9ae/+YWmK623
e9fBiImnGUMK/ae3mHdjSPFYK/ANudAPw8p8mLfl6cBUMsSZ3eyKV2VChsatAWS3DKieu7M9v5Ow
fSI/Zkpp+/wX/T7h+Cl/b7JiaeN4IvS0vCYYEiPbE+RmYZtCRO1Rvqu5MKWWbV/aNYSA4MS2F2Lb
vDnbqnfyVeuMIoezuOmIP7exj7UriQ+4Kj/wWHaZF0g7/S1ISRYp2Mlp0SAArjs0bt6RwADekH+C
cUDqVOK6MEbno3TpRPzH1UBstclRlRyKYgfDpgaUAhTJo+tdsDPtSGl+S3mWL230KxPGwRhr7Bhv
nRstlzqoR6AnEs+VFk3j+GtCX2PLLFMjPIB8vVxsA6JyUmvOkvl9kwBnGDlYn7xMK9CD94MIp+JQ
sPi9+twSQsZuM9MqHtw13D3wVauswPRmP/7g23BsLP3aI/jFK7p02yytLKOzb0OtMUJbN8/YhAOC
wfziqxNgVMd2klHHN4l+dFOLYFYyyC692XkQR270L0gMF8JYqFZc346UyhuGdoOrol5A4AIq6oxR
yfwd/yTlijKfuOGE4F6OW1tdTCD7EWLqUuaKJLV+DBrDgj+kXFPXTKOskgtkEdr9uPu4NQoflsv3
OyhYAgbRbdWMikVBeTBUaLqUYpMMWqCzX6RTS3Cqelx6S9dwGkDHPa/y8faJU2aalIgYnOB1BdJP
CvNOPdxgMV6KD9CkyS4KbdEodDRTve+Q7+7C4pAHNhT0X/YmNorOfESjWmZZ50c1WsLnJdwpVbGL
fmSKhPjryIqMajQeHQrqYgG6XJSI1kuDyxY+vjeghozGrgDBBDzepdO59E1BZ00zl0sML3cWJz/r
536uPKMeycyRnR2o2PGGkJH6XBGPM5Qjecasz3Jdneq0j5g8zpd6Sawdf+jATFP545/oRclekrTv
+iJri2ilLDmDEnrkXTTDPAGvyE8Ocyu4lvvCwBA2hOIZhaMvo8S34be5v+X8iTCUyf6W4VMkFbYx
AWZOCES5yu/9oFIDq474I018x96q9zT1iXCd8lmKv7iiz9GB9aCB5Y4mibpqx9QIUyalsfuAi0u6
rgarDe5HBIz8XrlN2NpbmdxUjN1RnahID7LtITj8vwToO6e0dYbSi/wC9zZAkEzqBsu5KoqTnyC7
rn7nykKoiu5vNQ+oOkbpQCkc5HDAXjiw4qHASrlo3VWqlJQsZ/z4eGLk+gSqIPXEtCE7HSAePZp2
tmz+6tWj53R0TnVQvD9hjw1o5D2GuED0o13LSRoe0hf1jw1twwACGE0mDp0spHgWy6HUdcLhXaHi
LyiA1q4ujLjZC06o1dSV3PGjRpNnbimoqJDQ2Kz3SA85BX7EvxPZy3xBA3LgCuH8ikNZSjAgPnP3
8EV+iE6AYCIh0eD/SfoHbw28Fso0Snq/gdYZEOegxPZEmvlfa+h2xagxaPNza2qMyjmgdqWggpcI
6CGmBjnt7VvNfBoAM0vIrSED6rTxcCYBiJWg28CKHsM/ud4Q7OTJ0AGF7RGXcOZzeJIL+1hcET9D
2kSAF8U+yrmUys2wIJtLwNear0vhzn1+ni+BS6MXw9vW0Jm2fVaL00fch4U48Cz6vVCnL8P311iO
AaL8fa/ba1D4b0CQ3eI4HDBkhe6E9UfdVwnu3biEu29wib/Lc5+NYPlfBwx842oTvW3H6mjCUfmA
PSinPSkndSHm6ipmV04KzYZKnVUPWJl3vOcdoaDJlheGJCeb9ACBKHMBERFFEUdC8g8QV10Q7Xl3
q4E0AoHrmXE7IdO0sKDGPyZK54WMcMUxa1MnlnncuOy3UQJdHTgl9gYtmMx8Y1wG1a52HCQ6d4V0
NlZjH2RUrzq4fQeFAET079wq2ftTTsb8OMkEr3FTOpibjUAV465PX+yAsdvvQ4jrQSwf5ao5rjI2
V+ojwyAZ/MJWP4uxbW/Qt/SDqkqmd4yTvQePZkX1Yi64rFPB9gKSUeObOHyxFpBZ8U4Ha69f/YKx
Yhw1dFci4RZ9Vm+I/JArjI6xCB/svrK2NGHH02cd7Or3A1+2VkBsbqcN9o/Fr0X1eEmIIkWDO2Z8
aQXBCOTQmyv8TaXOmRvLPb0Vofv6SmATNRvrc5D/Rai0tdzZkz9Xa4JMcG0m3Kqk0lhQsNYHnW9k
3PuMew27MKNhDYAYBAqowXbMdT5cYqRTWFiMGNu6H0Pe48at1VvvTbazorfTYIpzSZE+gs3zoGeG
8UYaTnGEWPZej48DHTZBQ93C7tvsOtLhrWYzy/NeumnD+QNivFuBD6uPhdkPxxB/Iw4VczNZ7tJ8
vpSk9Hz0XXP+ELw/s3M2OC72bcrBoIr43F90935GjhunAtxvfPqokfl6/sICRDopS1ycQGAlnUog
lprKD3lTEIL11J5yO8NEs4UeeAbNplaTfEosMRkB+4eRqofw9loNGY3soTKxaN99uWPQ1rW9OF+t
S/nwqPnCHAIpl9V2vIEp5NsVgpeyA9BcQc/hJFs1rJIOOXLlJn3cfTWX5XyAIk0nZeCW8zQfgZFS
s8w8VZUObGVTem+I6S8avdomtpBoU3VP/KJcWY5MiXcj3Rm+Rl8xaokfiYL37GuLcZEBS8h8+MqJ
7thNHB0niH79D7o5MWLEDsMlvyog2mvhfYW5Vf8unv7JcqVD63wA/Tcjd3YnGy3+aK3Iw3cwcBCm
jwbuMw8Eb6IAGgO0dzvA6yGXbocF1LiUz2e7RW8OSMnNksYRJjDO3Ov03z1YwvJtDoWK4ZdO/nBx
X0Q9GjxKV9oRClcVs206wY5L8PQH8CQG8jLAhrVs690P1eIHSt9qxjOO17YmQMXYHwfmPLHS0L3t
iHmp3Qj1+Mp73olNRpOfs5ha7MalPOUd/CT3Xx7nE9ulGVF5LLF2axuOGWBd/eRGXiS7ungKo+0i
33FfI4xa/72236wycbQyhhC8+HS0GCwQrOkgoWHe6zh+abxkiBc0jtMPPneXMX9Ldip4qADrnfpO
/2RKwef2ps635QeUNZaj1RCZwW9M2uSVL+mkVf/PKnZer5ddDYhhJY76X/f8980d95MIjIcmDza8
pKMjFzqQn5YygLzvRsznGceCCfHrnTybkhAb/lUKm8AL9LLn2BfPdv93b0GNYdvSEnNv9Jq//JAS
UdKvaieADekZVmzLVATcGoIo+PRmM5lh48DdClXV8OgdpV0wO7jGjfhvFpk+zMLh9RC+0kx1QxlS
mSH6OCVk3lB2vzBZZjRsgWPzWMW3B/1cMm2HXev5S/jS9ue8RwAXkmySxR1ufLyrdDav7j64nKe5
9DYz67dWzwuEQ4Ia9r1uGAH2OmSVajY9ak1Uh62umLC7serMhCDZjqawu7PtfYUFFfOkyByo4Dhm
oWotbn8RIkwBI8FRFtHL7lE0kFmwfwXAsmHzJwhZ9eo0I7D4lrDVEhIDZt+09WR7ebTgxi1FGaD1
sEa8hKgX85GYDVkcoejPQUu0nrrMijDv9mqgacx1V1BIm/kT0al4r89dMz2M7EmEgVBjEz2jJZ/Z
bJSNY/oOd58pKMZCq1WA/DvtR05c6tUKESwwiLagTknXgmhy36QUxQp6WM73kisuDC8ALyaq3OFr
pCQ0SfAn9nkHh9LhBOfVJyebG9WfIZVpN1TZ0n9bsq9lOmZHxNBz6xL3Ax9st+gNCXVMlh1hT1+A
GKV6FmkcV5gxancjCK2P+aO3tdiDvLsPLhOpfV0gXELX3EzOGvwi7A0jft4iVenSSUWMpiTzpMxu
F1sDcHgZNjjHw0FVLGUHAIARCii2OkcZo3PXDID1XOMkUvgdSjrdaI4pvo/lonSYutyZyp8L+LEd
31KsqXJJDYP/2IBuzZOFxk/qhmToF4LeLEpFiJ8PY+QNPfqdfVAzVTIT2OPVj+r45eM3o8UoekXg
N6+vucmLJtauSHTxIqgQr3ZKby/EVfy1rx5su9kjEFReyw5MMF/fThyRgfn5TrJhhgnesT3Vjjbt
I4cVxablA+yOlr5PdrWBft5yVZtYbR6MxlCbsDY8gfvlqUUDk3R+lIpY0NhAy9Jbk5YuoQUMyzNV
BcIpNp21ewO7PzZJi21m+z8gJRuMoxnWr0biuFn2x1EqvJWRaIZzW0Cb7NDUYG1J8w6sf62WNcf8
A20HaGAOX1Ps/CHkM0EIIoAU9T6u3DZURib8q2yTiIRSCewiYYw2quBxXr3NJhiAd/MHivQURDS/
ik1vJNHRdtUI5jPsiIBp8avEVOooGDaayWmfHa2cNuPQs/wPpvTXA8obKt4awGhwW5SX/FPu970V
wNNbPFbSaiGJ2fmdRHGr6Pc7vQV64Z5LRd6Cc5MvQ64pFVHkMs/nJeb8QzHfi2oVzykTI3h0Fe3U
C2wtW4GsqfJmuhJSXxCUqJBuOn+jUaHKvh8Qrftd4VDd6Z41Y+ispeWgxtfrqVj9Xgk9jHDePcyR
0WojQh/hxM36o8VaHMhbnRb2HPguXqC5ke+ZhQfUTm7J+xY0qNUzxw+PGOFyXUlJGa5ItOhgVNeS
fZBuOBc6etJTLBc7OB0k+2cjI1ln4ZKvnVrvi8sig33RLXyff7/u+IKWCP1pHQ+tX78oYHBdikkk
i0gAxEJLSIvYagfMO3aYbHOw88wLyEE3zf7ZlVwSlNm8xz12IfuvmVf2E/ycsIK69b8GcQvnDTvG
okzs0ValJpHa04zhOkpVskUI5Ox4Nn8CuDqPDfFciEd/AOD4eHOBeGNWdf735Rzie1pKwA3pgw94
OqDZ6rdHt5Co4J02xFq15DjBHISFL3q6av+N0nQyFgj9VmsPDeRQqGDSV/ZG+FH5V3ct76Zc0XQS
leWtgVUYug1RplHwDhbRM7+PlemacIT5bPxmcjvyo5ZDH9EC0IRlMckIjJbL3369GV01Sq6MdUB3
bcHie7kpTMGLjn7yR/46cY+JUlMUWSJagoL2z5lTS792WxDl1iQoMuRq6hqODyN6YVTKJuzaElcc
U96UHrfwS9AdCRs0SQzQPlf2AhWGWIxI3TnJRejMZH5CB0HpjOhQbwYPhx/z/RxtugrjkKJ2lt2I
I/tJQUQoiSH9yd2TLOJAolnmN3a/dWNBCj/QlwnjERqbfaBFkgqmRn9MocD040sWw/fYj2lAB4XN
TKCVovyAxWaXhhYjhf3ByyKeMG6G9D1FS9E9iI0gfKKvsnlEI3LyfvWbhaUu2UPe2LVQiaebJwI5
ZJDxtE4wsDHq/cmuFOUmU3KbGrGrBARjaDtBjAA5WqubR65qJdvZG4GYOBx6INdvSBK9wFjCxyzA
awT7iPK9Q2k65lIm3idfV29s7yo/iN3zva1PRHBUNmGgxTdhubAEvVuqJsXunNaOSJUKKOJPRobG
jKQyMBgFDyNMPvCId/uRcgpyLHUZa5HYF0UyENKg8LNUWwV7z1yjASIWRM+UFITXYeZhi1KbW95U
uFO3xukTJFRKR6N1XiuKu0q+Bg+ltW0qW/VtSJ2c/1Jv3Ab+BAmZ9/GzASq9Nmyfs7poO46oyxHH
8EKD294ZhN0n+p73spo8r/i+Se6lmijrImwfL6cGX8Db8r5VBWxDh26WCfCQc/6vMo3T++cEbjWT
Swlh8s73t6ucB/wdmirYdSFtNdTXxiXSpaxvgioIxqQmvxI8c2/02/T0eyBTqLY+kyQT2VN2cZFK
WoYrOPzZJbxtYhYwH8aMuMNkm/ucrKxwX88bCIEsYR8c4KxXE/iXzbAmn4qwyQfKxae6kB+io7Ab
XilJuA9Dq10Ykeh7lH3xeGfsnf9RIKlDqyW8zdH2WEK5t7fn8+E9SWbbbraQNrPabt+dhgSVfc+p
tDzOLlMgxz7b+Bmu1e10T9h86xc4HHAOhtUcN8ggScZUxRRfiw/uWJvxVx4b4vKjwUTBozfZFCKb
/kV4u+qiR9/5WpxRs5Rq1CtTe//KAas/G2rcXd9x31RBgM2+LBYm/cGOaHstVrJ87PylnTKhLx+S
a5NIWZjc+kaFfDdZWcN1HrAi+d4Fix8PFb8denQqHAtI88LgYi7qI0sjQTYhDGgVqLPtpSuvz4KA
16peZg14YJHK/ixo4cmYQgFiPvKT2Orqs5Jwz+GqIAN/cawng45ahOskBYhR9M9frokvcloSrkBf
85mId8hAUPSOhBZ/Ms/uJVJBRCiVAKotLtDmJiZBos+fS2QTc6H/9et7EDzHaVA/o9Q3cX9XD42q
mFg7i/VLgyTPMzQxJPQYpJbJ91W5/rdaT9Dca2k8AHLxuKxrtyX1etGVAwKmrVRKySEAHjDWno3A
lDAbD/zYeKjA2IRrdX74Rdc6ag7OzUOxwJ7iVDBfhRIdkuKEF4pH29z/aXeK2pSbSGcSnu56dnPo
qk9DQ6Vio4jBKOazsho4d+nO2GwFYs54pedT0zCT0Sq09PjHRYyl77NHNgbKmRamZZtT0vvn3140
yLmrWvmkoHLzp1z5ubLZopivIEgC38ic2oFv7JP/I0MlRyp4wO6yHRkTDishroxMS8iFArfXpwxm
338RLstzx7ciQgfrs5QP9TubM5fBKy4jj6LIoeqVU8rVhI232+PtIswdvHsk9RPluPtoJtEw096H
Rw++EyWKP/w8J4Z9qYd2Wg3z4+WhoqUREQdrPagAwyIi0cKkricRcueKbSU2lc4G8wrpL+e+ofJX
cjcZ3x4w2gICAdtMdMBBKI+Gp3SIHhKFfr0eViLyzqcHnwobtFAp13UFTGhFHk+qXXc9Rf3Y8YbC
8paLVS2QMB9y+GdBxNqu0in4aKQMT0p+4TgB4OAllCogYf9RM/vRqwr/Bvy2NlSlDXrODImUZFRn
B5y4Ud/qYEUo7Hjs/3g4HVI3ZoN9HHzZlu2NiREerLgOGFNXB4dc2CO5n9B6wJ7dl7dssb+c8F6/
KwqeiO4UzEPSwXRe5Ijr7++ylVXn+YQ5IK3CN+q3zzCMXDv4UHdbubc/Ni7tXsUlAcYwfZaSiMgp
lbOw5MJMIpxM0LwePCUDUMrjD9VP28JK4pQ80KHUD1AUiu6etHGSRXy70kgsLskX1e6nMWRjbL/X
i/jhIpAcpiweQYq6AIhbjOWBRQsNlj6umJVPHofEdVvz2oq5o7+5y50UTuT0QRLy442pfagnj0bI
LbiNggrd+noWuCmJNyfGz4e8BsTQsedeEjBxcRTOufRzvl12OwBs/OUHj/FOIFtJ5fFmJQCZdclo
tuw6Q1K0CBWxaHmlKgc42PWIuaAuM1w1d0U7ld8pG90r6blXaeJ0BuqfzWwBEe9t1OHliQwzkNqV
R5jIIUWT36qVRG4crq8wvCAv+4c2sbiCJcTV+IW0ojBao1iZogb+0rwldEoZ40ijja1wTF0bwQ4k
3BK1Fv2dIcbKKQY07xzwe7vOq0kCRwZ12dO/UedJgSUTauEkQms+52a2DxIOXU7XnACPsnoerhB7
kz+9Zp3nGzEPJMwUfhJxblH7yE1v8z5SFlj04T4stJsjiwVf2sO7KcwDam5/FNqqKlUxjP7Yv9zm
0QunJ3j56Y5VgM1V5RbSLp0YwrkfC5HjHczG/Soekb5DKrYMYCBjsaXS4ghfxn1rHKwJzHndmfMy
xOTZEAPdRqCwfTPQimipfqqZDyPvUekMbgia7VYIMdsiGaiV+BlWEWxO01LHaMo1l00TIWaK6Oqq
4w9yTJpjWBhPH+8Oa0rHN8eHGEJN8jCbITmAKMHnxNqamVSJFAsSrfaqVxHRCUBgetWGXdgnkTrX
8JbtNcfEnID8vwrd+Jozo2tWOC4opWRs8EtamalPxFW3G6pB9yBfnZJHpuUyKu55T7YbC5p+Gu+z
CN+he6Wm/LPTkT9NFyQY0x1LMQKxp8Eo3LYkArvjSGz/wT6liqWnl0H4gqfQqsYGTtdIMTBz4MOg
j5SsPoEFnedkPKxtDA1sJsTroy75BFgF0iTg4hgHOnO7xKU0/ikzN9La3Djz9d24RylHZoXHemAW
tg2TWSdGzxzFD8haYzrEiYxMFTqsF9dxQj4mXKPiXeLglEpDSvje6JR/urhriUCsmwroyHBJkQjJ
lfGRC1PlJAnqrdk7cfTdggdCfC2RCRbxJ2oPaX5808R7CwNrEZsWNehqmYeFb8suOl5tL00MdzYM
UgfdGcdRsAuIEovIsMJcL7AT/siIQdsIPegB8J0ojLyZC+M4zRDaFTT9deuEneZKjBWLNLo71mah
EWTF2jgmn8+dCDfZ9X2dWH3X2hJciVbOhotqTHIkosjWmq7GP/w60xKYUzeS9D1tUrMEZDu0ekx9
eaOlq/tcYuJqCMq4sb2xd/3blUX7P6IMFWrCa0eCNNuafKQhZdIMhU3IlrQASX5sEi6oWizXQmQk
cMlB3D+otlf+UyHCsgzWfitcb1URahxgOLPpCG8KQ2Wx4dXnUoB/BjSghCihJAnQCaLZEbsG4oKL
A4nKdMFJ7/dAu7/wnc56NnYo167+2MgVR3Raza3MtEcfx2/mJS+pe9B6tDtjVYiFc8UBKqZB9/cM
hKW5bxiZB9mBXsplMzaLDX74K7SaXoXjNO66af8K/xD+o/jeahxtwN5RpnXc+ABxQHacCJYjCNBZ
I6rAt4TdJAw1Co2lrHq3OAEzRqjkW8Fdn5OZcqLYob3WQ4VJ5mS8DxSpVCpMx6jjQVDDGQzzXLIN
d9LnmQIPyHL3u/GoU19O1K/5JbnXg158A5Q2Yt2I0QtYEbO4uck1b34ciE+Q1C2Zhv7Tuv9xnPUI
kqiOXBwgRU+Bwnubf/6ueS0eZmQvhtl7QB2lP8lY1a1GmklfdzS5fBbLLf45oQRS4YV7D+87Rlub
tI+5nK3xiCO9Lyxy0rmGVSythJyb+b2mBmP/iv7A6VLVtZPley10FEhAkSI9c/U5CPkm+qIfryo/
nVNJohq9gmeHXGdlhvsT8Lb0QKU34o8kPcuToJAZz8HpeXhwgep8qKNHfgDIrehV5spXtoIlcmjm
G5KYV2/huNvFWZsDF73/DyJmlAAjtVumemv4HYbfrZ1ZCkbwUHCA2+2Le4D8henlS8TBAKy1kSRb
onTKGiMRh/tgacudIve2GUgCTsZJuyepumVWxRlP6yfTl+XhOnwi/pnLhiZ9YxM/lSM8Z9826BcZ
Anwpkvz4kNt/hUoGeKx3GupqAfudcLq3NvRLNeG9/cCB4GtQx+qP6Xdt9W7u8mNcJpyTF1JK9kpW
Qe5FtMhvz/cdMafIrhhKAciMUZmwYqA1onTIgx7fOJFOA+U7FkIv67sqdo9fEZK6hcid6oS6yUfy
kL+3VyprsLYTmqqyq86u1Fr39u5mti2BFPpaXcq0AsJ9kXRqbUtJDGwuOIaGVshu006j6P9cploH
2GODmfLVvERaCGkw9f4XsC84DCAqTS2uM44I5XNCHTUzKiIOAa/VbGTBIBh0onBIwCzwed1sxTuA
E49u4elX8ArQzeBCImtppbkI6epVFkN4Xp+WJCMi+aRUCvEUAn2uPMAOeE7YoUOYIZWqD6FIlvHc
Pc67gIWvw2RJGi8hyYlwXHAVd5EBKvnZok5yM//8CTon2B7wQ5674W8lTQJ/yqxX0bq09MC5/kzL
bIstHuh4GQdHM8jrBi9BmHj7AjhUyti2eftNMcIbMps+9EwKx2DrjfgbkltOyWK5IDxtkClsEFh5
wwIMR8k3bHxpG/Q/9mM+Az4C+4uFnrLn/BT2aJO7AOJxXuJqd7h7HY19vTpxnekpBSxIDPC8ZnFE
5WjOoO73jv+r5N3YCfgUZTrBcAj2IpjaBVb2KhoCTkgriVxqvxeD8lH9IqF45bJIR6ixGfRhugtJ
DnRGPrN5OaMMi91BOT8jchZXzUpQt2vZD2wi5tr1mKviOywObe1wvOz4BD+6YDKNyoBl9ayvfjBD
PWHqxwHt2TTrensjagtJQUc+C7YAjhUKc4iM4cwODPzn7DbE1NqwknLYgaC8K2YGIDObbY5X7Sw7
LJx0pQvpiT3nDCh1AOqPWiLQpjvZXTzpCvcGt2FNnNvH+38k5t1pn1Tv229niOuHjoO1iP3gfCB3
7xMZlxXIQmEVz5V3SK+nVgQxCegdUgL/sl7JtdvohepNRYz43ja95/YNfpm9ROZV5L7YzWgJPi6R
JaHMe7M7xHZ/0fUVo7TloxPFccEK0KB9UpzqYnMvnpiz6Yrr2YgL2+0VlXO27qLLRiLcnbyCvy03
SJh4V6cgy1Bmtd6V0fRLib1wmCZzYCX4PbIH5s1DKpF8lQZ3j1oXvPE3mVfQ/hvQQ4eHO2scn3Ro
g3srpXuH92WYwwsb8nujq9N+twpXORs39MukIZhXNdlJiNQGtYNCMjbJN3woZNRZn41ZfR8ZRDdb
n0E5IlaOUcVx5yDhxuwZPM4xz1k5nngWZE3QIImZdXIUC4dTPbSvKpyEwE7JyTUXo22BJyXf+DO3
50OSEMxDxfjomwTopGfTobboeoF/qITO0/nV9HBKPSlg+QjmZ1FyRI3tKDfsbsO8xZF1NtTzZrUM
Ri/lklHIos7XtF3tOGnAbwe8qDw6G7YXZRaeMoxK+EOSyPPCvQAwT3YLaCkqEpMpxxt36lOMWg5p
RM2TYMKHjhA+HAuGKd/WxfBU3B6d2G+6Ph/AhC7RuaUy41sW4yKvApNfGhMJnL6h/bvR9UZPmvlt
Qz7FI0qQIbqmGW44D8EiKAMJ4YbgRRY7p0fnYjbv93I2VJcv7RW0QiitHodZb9FcerQ3Ahz3mvSy
z084UAlY/bVX6W03VkpeXaXt2vuwg3YYJL0Sf9/K2C6SKXCGOFndPUy+kLT/cBSnF+IdpWXyGrml
CPyadJBsAqApjsIcpOgv6acNP/sMp9wiFwVzgHoOYRnqDJG0YKhpGZAbLS17dV9ZRmjU9u9+Iazt
ijVQYOV9EudZPHyx4xywttL8AIA6epvDaVZpm1o37oOZOF+6ghd4h3sgae63cFiE0AE4jZ1gVbGW
VzJVbZcn1WTH3gTT1Lpo20R0f+Lu9vbjfqVFtV2L5oedb/f56OauXe/ZK4abCbX8L+4jOM1EArue
JdiYECfPjCip90JkSYCLaFzwgQW4W3b/Wq4xhw1dkDVNLVfj3422ltnWyJZrffdTaVUF50YBhYG5
s6q+thylsO+RdqOXNzaNXvuQNELhoTJYhVdMSakGq6P0O0Jf8oeC2nF9ZYzvFaIPAc9G59VOTBXA
0m9H3sbMp/vlcVjYC0wIPTwdT0dZr21DffSBFuChV18JeSCkIajiUjgde7gj0xQXePSQc0ALCYRu
3l8bPCY1Oth0fQ4McabZpTqCmxMA6jzwauF94CY8JXX/gSSHQnbEAEQvmii1HgyxdPCa2vkLc2B5
lYj93nwOoHiVGSqVwMfje4orZnWHfu69jpKwN7qFdQ5TKo+2s7UdEKN9CmOhnI3wyk0ZJZLRn/RT
H77aBVsxL3c/jlLI1RrlNwCzt/LSyerBdjTcM32ATNSbstFckK6Iws+b0Trir6m9veWuZE5ISG2o
p6dcy28WIN+3cPsfJSXz8uRPgGUvRWU7XBgQSJFiGJ28IN3kuP8ift1KfnJcBoPKet2y6pbNxTo+
pm9ynSHrfcprHX31D+tlnbTYTorJevqBCnJ+vu9imXzXdwODlt0k5uYqlkyqerlhPUO/FaGC+ivB
ar7XvlxF0mdGao6ylfJN/v8ohfh1731d4O7mkFJ2UmD6l6f6oNumukPA/a2OmnyxwQQiTwKmrqjr
asAc2UeJJsCKAX1RVK0gYxmaHZGq59wT/FZqPUS/ANSwy1kSMhut+sxjPqTQmwRY9wZgC2xYRfkT
TTUowpgCeSOBhZftfPTVBxzhziBtsRHSZZ9z02ZtJVOgNkq6Nv1mOEVCChfCEXYaTkidJuwrf8io
W/2bWbbvSGFn1XzrOQ/lfEHz4QOshGGjbTnJ1rwrNdkDE7KiSRLvSHPjfAFpbctQ/hdCwXpHalci
IT49c09uMHVt5+TwdWDE+yUZU+kLoEvbjr3y1jw75oz5bAL40NQVUBef/EBjWTjMZv+S9FjoTIOR
fd7AxcDIHTNUms7uv62nMWyX4OqOGqlkluUyGnsexcPX6HFnVTlt0YndMeACoVV6bWNfOjGA265B
WV9ZVmaN4aRfL6LynU6DleiLx2XVUH7DpbBhrOmVhC4IpnyPFAv8VccqOl26xnx58NyuaNaAarDp
IrlLQRZUFKObq3U5YX8U38XAFVD4s4ooyshdWTg5Ts0SLCTQnPFnauYgZHUi2QgVdwUB9oBU0yks
oJbQ3SFAU7esZZGeJ3Zkzq/k374SpJ80MVwsYU54kfEyeoEBndBwIe1d1ErDVXYqgsjMk99Fsd1E
/rWm4HxW09hpWM0f/WDxmbOmYGn3KCAuIzixeG2b2dlp1jsFoDeULG7xHUIVKdMyZxtHwAo4lra0
OIL/uBlsyyqJK81RRR1j0d39KMTuQD+egQCUXRpTkXMYvt2gq6cKzSbnwVGaEtpcpShkgmCMP73H
wOaD4KZPOYMSeMUmu8npT9kFpaZkwv8YT0UmBP3M/GUJweiBUjQpZHh8UzcAbQ6R+xEZEePPHG0E
Qug89melfVMniiFTpu8BbclNbhQH2UcwT5Y6SA/mmn2L1OwPH2MzEfb/8j4IuMn8RQYdUCcc8mQq
YvyOchDSYFksv3lcv8cQmV9WNbcPJ7q7OvBsom68ekySpPrx/vySogZE6K3QQbXs2HaMADEVPMvw
vRx3bc5vOzz6JptkleLq70tbuf4quawY4/euwoTZwZaRZpU3u7Zs87fcgc/84iRPnFxy4WNM45ST
m5Xn6PU4wztcjEkxxotO3OF3Ce5Usv583WkgLxnnRHYHrU2ky8a8QCew2UojZXhrVMdBo91iVAOD
XZnIVdEBxzvbeu3PlsmwglRgBJtdnEE3dHwtfr2C+lgkBKEBNgpyRIFrTjWLfT1MnHN5c4deE/gT
dXYVHQ/Z8vRZDzPA8r/xnAc4F3D4vSvAF86kWj9blikSXO353/ZPqLwZRf+PVAbNAVfVC3xPEewZ
5hoa5O6x4PI9Fvoikl/Zpfu6vPf0RurcyeA7hhlfeSIR82k3VH9j+GqOsYNsFPJADOkILNdRYqmK
6raYjZv2bfSdV3fplk+tKFj/HyzkqkGvo7bQ4T9Oc6jGqzw3Fff2BdcL8PXa04Gw+aKz+N1lxmjJ
3a+jeM9OIjUu0ToB17QENEdGkF0k9jaJpyOF3F4I6OFQ2hGj4Y4ydIk0VhzEsNtY1xf4o6/ixir+
RpZnJS1FSapW2RJJ7pjW6HZfANSLUNv0q5kBUAIvfCPDQWf6ITdeeOUtIT4yMZr+wTBFUSMYyh3R
YFpup9c5jsn06TjPS9rM4lnAnylG3a+xc0TMO3N/h1keNy+yry0mgN5+19ienhXEnyR+Rr1N9B+k
uRs7/V86szpEntQV6ANQAn4GdtgLHCKIk1uMXooS7m98cChqEg2PZmmy+368OnSps7kC291RD8sV
tM+c3FUq/xF8EPYbr2ZyR15n0fJqnVJhk33k8DHL65oPNYedh0DlI/7laPsBmRY4Gx4AVnv6vK2n
ePAAPDbgSXopegxmUpr1iWtYA0f2PT3NyzPj+n5Z80CLAQ3OzVitJamj+vpI3NG8u708suxC7DFb
ZIbrvxdUQsslLaEEgxOeBuxqO1ZpYigg2620P2u8Y/kZfLzoW1nY3pOTNXFDVlL+cY0yaL5RAkxd
zp/4UKKSwmXAvNvU99i5ZqJCQ/dd/phTQwGFQIYKTNmWwvvfFoXLCzX3pd+T+DXFgF/av/+r6Ac1
DopzzYAbI9kDtO/JXIKUx2lRty2ml3tH+RIwmVZJDw7YzeHCH18hox6XCS9WTqCwqi0jF+pJERv0
XvK407Y6uEskoIl9hgtjKjeCzYn+8nFS5t/uY9aH7/D/70bhS20S3y/n9IB53E4so/v3O16UCcNJ
DcfDFjYqEusi30pgGnOkObbPzWEQiSBGMyL+c0FYATNt5MXGVsvimapjrWif/PRaieeV4Ia91ON2
DW9uNd6nuy0Kd2BJ32gvg2XNeW7dqbhZT9+THj460Ej4CPzR18B6czhk9yGgru+beWQ4WIV07x6q
MXqW5LKW6JPDchBmvlcdaVYnq2rjKTyY4JEGfcODugkB9AYDzJZ8SutMhM1nReF8lN7KcEXUH/ve
l9V6Fik/Efq8yLmf9UwGPByO+5WVZxiYX+tvTKXHb96UWSI34oefK46xUa1JvVgzCsoES3Zs/LRY
vVFJgahSj+M/1bbYLB8WV6dWrSGvqcefel2DmeLkWR9L+778mmHJFRWQqOjiuIlpgEj0vrdsdHkl
nr4r31isNpKQfR3iSyyclab3t/76AgzHvpZRz+kFdNuvh3tuCW9vXwFM1EFPlBEwKW5aiFsZ1UWA
FgMGlHfe61gIHhhr7vMaslT2y0gQ2YgMZaYBGKhY1Vl25fyzNm6OnTzqSaZsNacj+GLRbBO9AjgW
yMNWUZprexRThwzwcsXFMjMxu09GCPs3+WwEb8fa/5h22dJrOBY+gwZvmPiN/6gPa/TRoMFzFw1E
X4g7E8VsEWO8+zwqCtRUyy+xmyP3mD9zdconnO05pW3NlSg7hfXAxHAcChA+U/nJWdRD7nZQi5Av
kih163cr49D/aFghFxxZrk/U4DIfM+pBvUu/ssE2/6s3exM4rQ46im/rbDdppFQTRxgCSpCw/ELr
tYUslr2bHSdahkN7OIM4pJZNnNbQ0KyumYuca+QnKS70s5g0E17HZXZjF6IIWEo+K4p/8g1zJwh5
Z1aRh0wHSvLHmvNY2cAEJLTYsxj0FfGxzfLz1AouJ4OoD8135m0ZWQTmin8mY4XMnaN2FLRxObtK
X1pWCeueBPxPa9L0J3B/Jr5Hx52Xp1aEjvNkXXY+5Iu9dAFU5F8o/kXEswAFSg0Y1tUNfNwHXUKv
GwxHlmIuCLffuVg2tONC2TeW13LYxg1jEG3zZjICH/HHJFffW+MTQJIhIqoYeV1gEEQe7v8/0xMb
SRJ7lGz2V2hLz9XKCUKTF9/qf9VO2Ztwao7PZXc4KqnUcZ2gn3Qj6Jr2CG+yMj8fr937HXfBo4GU
PAZAwzTyOfDBWfPYoJYy4dEiQMeY0IWqfO8ijz9ON92EvDFRrl6NRgOkeu5bXGfaH+pFHXwqcmKp
fN9necyQA4HkQ5nvDgbt24m2Z5xTAxtqu26NQ1ncIGlDXaIiJczYeU3+HOZUy7Rf99n7Do3xszw6
6xLm5Bz926AdR6/YNvxFvFoKsxa53q6Z2cCOY0pxK4ouNIGVx0NiAXDTA84hcF9T+9+Bf/P45pLb
EHH1Ef0FSPdTJxmVamLLRAyV3uTsOCrqbIEABf9fGl02YtLuKLoFY+zBc4fQBpRpwLPT+BApbiX8
t4Gh6Pdq9nwFawdV3AfC71lekBVW+GEFo/wuXG2A7cFBnHPfSOeyyLQ/zfOhurfKGIAEVNv8FS1f
TkP1qBrdbNVq+v0eKDD/AWzSDvatS6vlajRhvM2wzgbWFRjzaU/+TSfH5TmkL0bw5NIV65WN5SM8
rfVo388WMxIMZZf3ki7C/HBOOpaHFpJoVq55k+puJFw6TFTnLKiPrSgELVZa4Dm8CUXjN/NjGJ/J
nvmpUnDlax0EGvb1CJlWQQZ0E9UfluRrLUw=
`protect end_protected

