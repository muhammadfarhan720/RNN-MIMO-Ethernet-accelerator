

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cFLsLGMxKc33uWN5++EBJ6nM3nMjEzLyDOmVCYddEfhXxhtVdI8+aatqgtp3Ba/l/yCezshycBow
CnCejD7EBw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ETWk4SXvH4Fm2GG5jH5kM4nw+ZExM4GVvWt/h6QOdFfR6hzjEsB2QEjT7C3l2q37sLhkRQZRDPIA
VFZOs2DDVSahZbmMx6QAlcERXIJLBaHD4yetDyCopP2pbQNzFWvylwZswPiAzdXpHqDbv316qfFt
ecRCgYbecRif8TZ4CZE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jWy834UKSxvxUqFpm+r11KZ9yLbAJ1lAvL4uxx3OnSEX9mS0Ageq1xbYZyy1EpaZKyGfUkA5rggs
v/x/bT4ZizU4UAqj1DZe1iiyFvBHW4rb1N5pKTWJQT0nyxak23vI2HogsFtAcE4zEyqGgPI75D8K
JO0MgWaskqyXVNIUHcEYO8ozAOwdaYl9/R0OM+HPCsjZK9Aptm+7cbvwZi9WmvVgiF3I+DWaCBSp
cY6uH0pOJwxT5rKVl1ESfXpOAVgd+BOcgOKLqZgxV/8QqwaW7zKB2lR1WVpXS99ZJ8OJdGCfwTn1
peZF4vunUkGRN35ERausCEg1N+C+rMFtD7CEUQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SzqRiizwHNj8XiIh+k1aSfAq0u+mpl28JWOREmSGQCRWxG2UFkqkMzhl8agNwc3FIUv1AcvE7WsU
in92k2i13g/Y3RhzZn728l20laChuMuspF8OwxCQ5y9zE9b0Qjv5xeMveaFZZURlDGU9VoXyx7gH
RsoWisoDeK/JsWEyisDqO7TX0en2dPFjo+X3m4qjfUMALc1arQSapi5nSHD+Jt2VdKBnq2S1gRK4
c6bJGKcRFqKDPn7XrFcLGWYOC30NaNDF3S4b+kBUKj2A+TwFG23QPwbJos+9HsAGWkBJUGde3PD8
7EnJkWnRA+DQiBtgCPM8zJXbW10FFzLI556c/A==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
R3hRIITdekJhp3OnA/czKh4heCRUIzNSE4wxnFTxGOMLXuH8BNXL+XznRcmGZAQbvP89bejqpT9N
RGY6CpQ6DxuvUpLRXdSjd7Z3kZmWuix0Jxjifw9hiMwkQA1DUFbRucdhL7TjHx/WQ76+8rSmhxB+
Y4t58BOlYB3qUM8VBL1Rs2XKq5teda4K/AnWiO2j5+nv6by6+gUJGN3hGLxbTY2jqzEmKkwkaEoi
D8YRhOIlUp1FkmsCGH/ZNk9J4LKRZEJroOx+EG/4kEWGdv3WyxxYtuYI2yvKpC31u3anovKf+ILD
FgacNaxRB39s5Bzv8BZCZIQWzpGrhXVYFmrYQw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FLGAl2I3wwYpH5U6kXQhL9ZBuXmpyFhj3nJqITG5LW0zuaXgyQZ7nBXL/FL1ItTAnhNHQILPagts
zqnWCEqtVHTanjBKcekiLrtqa91iRZPA1L9uzcU1y5DCgPMi0WeBrZ3LC4a84QIxBHyjpYuBGqyF
/7LJG8c4svQUJwCgyt8=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nEkQJK1hPP3UKQAAiRULiqqcxrFKkfJi40YQaxV3Go2qLxwP15ZcLIN1m4vL1tjMOwxu3XZieQwM
HoEMQxlaCa9rhNgz2fJ7h0V60+r8OJNLzVX+sWyYKop7Ti/J4FeipyFlxO5pvpmMB6vNPvSoLR5q
M3due4PkKX7JdQJa7aZNTka/iG6picJK3XOVXxHqAec/j6Mws2amoJTirhIQSiIguyTbbezVK8LB
HLRKw6crlE7XR+N0wm5HJyeXcyS5TtjelO5RkcIL2p/YheqBQaqLhN905ITiRTZVS0W4NmSFTpgG
wXPS5xON8xpjJ31S6Pf9Nm8mMoO0TuN9aFLrjw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 506800)
`protect data_block
Jclb3rwQ59WRLaqXFWiueEHryIp3hjP5UIAYyu6C+l2syOIAdMrCQ6Ac4jJX3Ip7+L7E6Am2CpWZ
nrlZkMuwRPwvyW70uFYn3pgGrqAxN78EyJb8Rl3Cw8BE4nTgM9qgMuh6ZeoFJx+Lw329hcSyxwtL
wWR0/ExvXktsJnJeQI1a20erZMsMVVoMN/9+vvHt26uh5NTSWtX8K20YssUayhiJltcA+DTK6w8F
DIdbaM2LezSXdKlxiq3oowld8x7AHDKgX2XuNFpZbxdWXaiyQjakJ60fUoQJ96X+LhfaMwJP4f/q
qDGboRR0IllrifghEqlWSTe0CYm3qelNK1X9raAQ5WjYs0B8UyHbZo4mn2pRW1YPaYV7gPcjjqsE
wjcx5ixvsfUZoBpo/GJ5pzzNntIvFWI9cE/cSUWGVTBPMWU4eo+yDLkHz6oqXx0tLT3wwQ8knIi/
1ieuqYYeJsNuFbqM3TFk190yf54wIqEw+n6NBYnCNjXQC/qc+2MymxH8s2Gy6ZW0StBdWJzF5QP8
tUMWgTSA7AJTAWacEiEEtsqgKbkC0eUqR8sxmJDkDFzGi82ClppJ7WWQKzfDik/hWdNyuifSW5E1
+aBeKCQnRxKbjmQA7CoFTdLvzXwHaJYfF6peAFA/QoV6SLVw29n78ueKnTAS2aKCNIDG1tyzHk2N
45yJAScqqmuP8tvQ8GysjPEHhfwpXrUd5GVBxGVC4F+Q9SpjbbtOm/fP6lixnKJH/ZazzR2/wVVV
aqQcb46W8js5R6nGyeksz83n+T3DUE14vaDMlu1kghdf1rGZdZGumXZJHqvVobZ9tovyXk97J1UH
bA4Fm79of6brcYBU1mptVuIhcQn4ESo0HbmcewkajSeTZdXQho/GDky1T9XlKyQjeB8+PJ+TKyT0
QexXT43zxPuyREY/gOJRSTikh/oJaSotU8zEyABQQsk/crHcWjPNPxYEALGJ9GEfgTjT/ASJz5eJ
tYC3XlTjoAp/97OfNfB4IOj1BgK+hVWJmOAbIaSmUJnL2FfgnlIfgcvee3xkFK4cqF8queBNIMEI
DThNGNCUJiWJH9iWK1Guc0zI6gMXYUTPolvI4Fn2ICTVBB6nKP7zRSOs3Krsmm1aoK/U+jMsJu3B
BGox8dB7S5nxwvGxZ5fp3p6solJ/N3lgVJjO4HvJYsZ9lUP7d/lgwKgqilwYa2c58U4SAkiKtYko
mMaOE6NaFNT09jvbk1961KiVfpbIvW7Htu1G7Dbc7N0cwj4eVj206Rq/0SBB85lemwlYciE0GYEH
W/goezKnowOH+R6tgtMbyBNopZqXeOdnJj0VABnHQ4i3nCz6fNBWPymmsC6FxW1TiURzo8VwW2DO
s64vWv1hjOTTC0dgkPrZv+NNyUGywavk2rWubXPw6RZ7M4OV/Y3q0L+yR9Tfqbg6JfeBxkZXCIxm
OnpjupuiCS9rLeMouqgx/AW4P3TfSK5XhZSHk4cYIuZ5uxLMWONzZ2XTtf2ZT1FCCFHBuHiOajZL
g5pbsP6K6NeO//2UdO0UaJR4cXjT6GXzMmyMCqucXrEZslJsaTwA2gFtVQ6CtHHVZeU8X29IjB3L
10rpYwys1XdBrwNvY/AsdVHHemNi+Bi4ENAmlehfpEY4Inmqs2U2Yexll/wNDEL5vfdYTpJ+/x6n
BgnV2DlkgnlvrPKqSM78/laXS2s9RqVYsn43ImxexQESFJK4wiEEsqImvXabdwvRyc1fBqdtgA64
Zj7G9S1ODbQP/rhGSOS3oQLRcSJc6gYeZwEv+MsJmwGz5To7eIbm9i9YVdMQNvMIEyzzHXkpLrNE
qPFBYJeS1fvm5nl4X2QJJ2ophUiTyBQELvjcfPgfnIxAX0hcfRx3xW6OGHdN4ByqIi2ofxOwgOfs
goFvtEoeyyCbtroVSCOAHc9GRkQRNyOdC0DxRv+4vFPU9mLegwnT8jv7t8w0sWYDN4soq/tLq19u
C0B5IqUS3YcK/bxUDQM+dbrUOn1Z99bgRR3wb7FmmjYMs/pehNcHpqblr2ooUpWCkkHBHhcaLPHq
Ztio5VaLwYNHxIRnonShOvEPeeKj5JMHFTI9Nsz5bsg2pdwxauyqOQNB6CDmPNadNiSJ4O8hGEmA
XsxgzdHh5ZmNkarX5Tx/rvCQZDW69kQ8MKf3I7bxgdxx5/YnJErPsSGlIDHhI3s5lLFdTSPZ8/vz
G0UtcsPaNjSgKUCjSDTIARfC1TnmRTO+IWTQYg9EBoDYe0DNmlvSP05tgpdEbMulGIffK6c8QM1X
avaqvJpyzZB30srWeOZb/1buKRhjHobhveAaeE4Ssk64O3fbIAyQWe6mNcujh/hs7LKs5mnGCLXQ
R+QdBCl6GPgrgkuxX76quYeS4edzT6+VIsl92vSKou7SOg5Gw6A2j7OiwokIB/2tCC5MgQrRUz5H
f+OOz3VyA+uzjtMynC46HSEZVIHoxFZgYe4ySMr535zeX94GalbEQuwCmrgXXZ6Zqi43+w0OO/Pb
JScUSHXQQ5IL+Clo7MQVH1aCq106ClFP4+LbuvjXjWM+NGjRlmvjeYRIOeCdEGRNSmDUJlkH6Pwi
rolydwnjAx6zVJzSV6Nn7STuO6p43ErPrQUN1iV7EEwDMi5dpVWW0FxKdZe+q2QSTvneVHDWwq71
EtpRgp2alp/lqOYfogU4BX1itSv2dMo3iEDvkYNvrd61QLuA9uR3S2EFZk9brxIBh8iTufj8INVT
w/pAbNf6+tJoCBmgxv34+JvC30/yk5Mhi5ySpj9QeSigdZUxj+MV0++6f/lEbmk1NrpID2aW+GbN
GOCS+r8FG+1SUjeK92mBAaVSJ2V/ltWGJJWc6tN4AfTneUMuCSrWV731SgpoIgrLd8rA7FVFoROw
UUr1KDgo5SYq3GP+QdSoaDFat4O5zLei68cGCM6Epoh8VREPtIKP1g+L7/afr5CPoBnvlXI7oNwZ
0IAl2oHA4xaDKR0hy7rePowp0OjFs4sBOv1sdWojrZ6dUdfFNfc328oPpaILI0ZmTZSUzMF9mSJU
uA0f7tVYVgAt8KlFzJUoW2mfcmZmbCK6jgY52gqhSY/o5EM07KDguCt4tpIejOKW4gWtndsjf0l6
HZnS6hpQ2ek+PKnkYY+T1wikr0jA3/pHV8XMyUCom1VCFJ91PemneLwbZdkD5gUOGrZ0re1mwEtg
5Jf8ArtEpW+t2NdFIUnaMHF0uWoxqXsX/Up+4gqkD5W5GIy7G7yEkIB+c8z88BXxUvsGyF2oCldF
ecm3HAi5LOFQ0PSO6BK5z5/XMkr+5MxjvJRu2q5S6Etn+Oq3olmp3rnWQxsBrFSJjFu056M8KmYq
Z1o6ZZJDuUodrmtRm5b7O99jTt77pC8bLEFkt9EaDpYI4NK44fiOhjx0l3hILGMZ7HbYcJAeECpd
dgldEXXswqBgivIyTWIlWLnQt6KdxnjugE8UNIXKo8gEVk3SJpXKLqwEcRVt3HeCIhJzy61SCuD0
fWB92gjvodFkhug+ttqhRN5NgckGHfi9rUUngW7UCRHqI1K4nCmB77A+kNXWQlYb6nJrzdg9o6so
6V9lascTD0DeUksy0AGDCZfUc4C3a/h6sfnJudOGXUyvzKxBkvGyJK9PleMsuTH5rmaNJivMlmyV
6Q8wHMAlGB6mzBA+GUgicIWIGnbvVpWKlfXFvi4QZ2vz+7q4Q0WKYdh8oZ+WdWoj5sDgYUzAt0Up
H2vikdhIzmcwaQyjrtQDU3c6hjVB4lzyp1PiJWENNRSgRur+ZO0UFteem3fOrJfo2YoeBBpU+jef
UBTUx1hWmsi+0aQNQWHcBf79OtS385nWGFKqyenRgXicfisvc+duHp7vzhKTAfvZex3wcz/Z2QxD
FiN3wcYmhyWtIXJDsc9vZNWeg+j43XyDq5gDaiwz4zvkFoZnTl1cBgbNL+48jPnjO8vcVYNbvx/6
XehPw7Q9IcFPtNUbyAOP2zRFs9sc9XFo8raJTm2kHbenlMj6x8DiiERNkHdgAw+499BMSMks5Om/
ocYhXTVNO7IAb05gQdx+yPG5SXAj/1cbDvYxgWorJV/Owa1vMh0b8x8tXvblNSbBAPhm8lw8sZti
vd0IqqL/9VmmMr74wEYIxPb/Tf86uRA57VjQ5ykM6iqOqAohUM9Iz0GMSULPvdeYgepsaA+odfV7
kr/4c8KI8fur5QQIQELz3p6yx7ImuCwE5w0UT57IKBFfkpOXvZ1hCf20xqunhInUSLZMsqM5ARmt
oIUFF1EHRn7sAaUmi9hYFIu3pvHhWuuCO1wockm6Q7+V+oi1S2cll5QKbHYbEci9yuuGkyrjbyJM
wx1YoIs8DBotdb7rofQtZcQwIbPDyj5WAkdOTowiPy1MbscNHNtoV7iFMHnzpmRi/FiKXHz8IRpE
1yGL5RR/Rjxc0QeXspvp0xNLqwJNJ57v89lPBvyWZQHMoJofOtDqvY488kxI/Ef/sJSef4/3rNEQ
m/JWOWuQkNjzpsgJiUNQUR8Aikty3nWCTzIGV8nwRfizJYdxmjR84n7cxqFH07JAGgMU/sFrIgak
0JnWCAWAImpKhuto6djahExrrVIsiCf4XGkWbdfY9RNacVW+gWBlPJtL/PuqP+PFt9o2IXIxLCB5
h3BJKvvf+uriu2nzCDxfkmVzVw5UsviGgNkxOujfgVOCupbkmxfOvCzKvGZ0kUYc0eR/k7VgFfpz
/tZIvwKDfq8wp2EvezryPjH8vzMTkGNJ5bIDrAQ2KsNmuvJd01MKeZaC1+jjqmUSVfA3xvJJVcOy
LXZwFHzJ33OF0SSOsFmBbVDfdLsq/vJ6l148nRuiEOv8XK6VN2h90Qq3TdggIOeHSdZVq1L+ZKzm
xpw5dBiODijJLdgEpy2t9KPFBLbPWY71wlVx7+TB6sH2c4wfnhU+TVEi+Q7fGJSZ6GBKXHu34gBW
z4UkM5yemuSMpmK22OopDUsdsRor/ssj9zl6GYWIEKFpSUEdtMnV94vziSLIod2kOByRabs28inE
mUMh1/IJjeh4eJOvWrPJFivuubZTGJSt/7G1E76CgaAQBDhahBJbnqx+wYHuJZlO46XhK2JRC1lU
jXY9EoScuEa+u1aQ9ohfs1A9iDWte8rbm9mWiv4ibtSQN8rxC3AxRdVmLH5tLHEdfE1OfQNaeit/
kGGFXB5Yeyqmmlrz6UJ5Kr5D5IdUEV7NNcByE2y2CFbvJDhSBLo3UtVn77PhuRkszvGTVZJ1BMLr
v5y0wrxNF/X6CKCcS60EVzNDQN6TSPB06jCD1Z/dIIWREbHwuX/UkYeegFtC3ovx09d+4mv7+1/f
OsnE2ViA6zxRAui56GYQZifB3dMeceGb4TFvrv826E1OpU/wl/e1PFZ2VhkdLKrrX4XfOe1vzoLc
rrUlDU/3KzEpkkF/WstFQSueQXg9ynPgwCCq9dRVa3cVJblU2U7Hr02ZLNKskjLKgG33XNsWT7X9
15UuRmbNsGtsBwq7rvjJrly7Jq6OJ3jjpi0FJC361yjWYKnJ62/Icz/u2dDRPVTpqxhoEyfxoowh
iD4WVefg/mISgQWmAwqJ9rNe68l2lqTaMzgnBJ8XB94wZGo2ISxjUfINqpHsD9NCw43aAxBFyWBE
IVEllJ5YISHb+pNlFxWVHZrN5f+0IIZ1zuG81ZxSKneAgiizkch4d+s/ATqi+utg3WU5W6wp3DzO
CHbp9oCTqO/dod1D1vJu0jA37Ih16SYIgT599s6zSeJ7W2+rIQ3os1c9W240frhwxkU8aB6WbqQB
/HTNo2QYiY5f/e4164Roh+6VotW/3IozxwhJtgUZ9YErFeQehcoOV1AjXHaKs7YjWtf2X4gDItMp
YG4HnpwdxE8kdRvEYmHPz9M6faoDi5uEKoZZWKCVA7xARARnNRBwh8GOZuH3Pmv5UXTnnmDuGkY0
RidrlS+LjXHbKoTfBZ85fZZjKAHkfNk7PGhdVPeK4jgPA70DzGuO0vcdpkCaOYbp2+tA/PflG6HG
Xx8QKF2ml6n4AxcR+KrphNWRRxX8LfFwSjFL1XKmMwjdD48/BlqFYNRvMDzc6lX4s1C3PPNOs85Q
QTjJuV9fUeeJuF8NepdERFn08aZS9r3kofL04+Cf24NDgHsDLMY3fbrWuZ2gjk4+vj+JgSatb6rb
0CYk4A5wyBiLPYcR+2fjhgJuShhAuVcYGsKVOG4Czf2SPe8KvIpV4SAFYt8iVuadFeBdkoav85xr
Xhoqgmo3Yh7BGyZBJ3MMwqx/Jhuyxl6p0qnowLPiedXAcyI5qUMaSuJvhbIwUTbDaFk9gvU/5Uuq
8ptDlldGEgRK+52j95ba/XyBv5mDU+Ii4INOoIyMiRSJm8rr6+reuTo3kgBwTlVs0DphwjiYJujo
dSJgk9mOzsemGtKLxOf5SDdUNwKzzhE9vqr9xYayR45d5N870c8BPOjcIWpvbGYUSEaRkRRSgHF5
uOqjBWu+3MKTi9/IiFPKdERPX8Kj3gzKe12c5iK46s5y6a63RUTXR6Fgf1gFPasMmUoDsBmGRkNn
U1Ui2qldrxxOyCAgox4sIKLEXdQW95bhNkydlmGomMR2gSsiXJk2P/vkzcJi0HK2qe3hBR4T8ZRt
Jj8T6ULfNh+zsEDme8K4OR9LxfMZMr7qXWlXdp93TYbfJAifXVTqwrSR3/9/7LvlZPxf521DosBX
6iDBrpVxPHaufWQAdAXSeM2wB77W2E7ZP0rsTZ5+11fWRvg4k8WW2c+Kenv9DQLL+gJ77Jh+7yqS
ljTqUsqRnLBB9m23xz9mizafMayugtpTwNXHhRhsK4nP9Osi00RS1fWPifCBb6Z+xPScpz48IcYa
Irtr+Pmb32PmCNvlc9wdZSL6XpvCCSKum8WSWh4Y/xzp37sxMwEWl/VOCZwWvhvo62rlCt0+K1E4
p43EN14zreyEg6iHMTcq2M3gKeGkVQk1HsmftDv0GgUBuEdOyfPYXozhKk0vvf4+yZKK4qJlcFqq
AfE7pD+/ojwPZq2keRHnEPXUhGQM+xS8NdrJf98UWYql4Wq/P9FsAB1WX0o+R4IsUXdVOHYHTpgD
4xUGQP5w1zV/QViYWHY+hFELSK8ntd0UvE2XzPWXjj5ZGR0fulf03LEw0TejIyTAXc3/atd6fD+r
0UigG00ENaKC3NtSoe0QTkN12dNw3yo+3eKvqtl0F6EckWn4LAxYCIO6bhT30yj2Hfw/d/msBxX4
Kv6qDaT9JpUz9T3icXau0qpB6AT1ADPmWM19Ock5P+OCPuTcSzBFRsDJvlprfUXhtpGCJIcjF5e/
R68/gvMLdtvZstmdhCr79ph9F+jsGEEikCv9h6A98NBxCy9xpoAeN44txLQHRR9qk1rH9PdRUEZr
QVGi5LQFM9795FrF+mSuWazbrycdS/tSGF5GwGDtZh9ogx4aj67Rvqo2VoeQsxPp6DJOhw8WhcFM
HY1h9HTFPcAGMkjgzft0lVxvoF6ILVWLVFHB9bSWHo3/WNUODCUXT31Fprpvokzn4Jbp2UXIJkn9
2A0XCL8xuZ8xMu9NnYc49fuy7NwdSVQHs/11DUIw1awpQc86GP2skuycexNrW90WinPd9GAbhYEN
xKS3fP5tcp5We3DkuCsxWI1bVL11zogq95aWQUWfFoIScFDe2xruiJLfN4PbnxQaxTp+1RhlGQNH
X7VQrWaCKmHQzo9NRjywANhrfkInVTK0f+HvE0QYnEoNoltj3cZl+jPiE3cqMJDUStqYbQ5Um4a6
DNNeXeGpVxKZ0eMBihlStOvzJl+svb8FH3hOaHuuEhBR5kb72fIyoQi5uk+FqjyVGUYYaTFp1+PT
T67D6OKZXJp6n7ShpKD40drmbOK8/UfLHOUSTz9zD8wzGGCw9W8z9c6ohOIJqQajQbbsXdHmT5BV
nocOzPdqXlyWBGIFI7yrCSb/oRIIUs5Kcmzf5CAsAbXUG38na8GRlssZc6FHiml6A+rJOVa+7tV3
vJuwsdRfNEEky0fI0N4927WV2UqZyFG9a/OhZLI9M5Rs+OBayKAJKoVDK1JFgznDcwyWol9elsyT
WtpxzEKm4RlyPi2DBEYBiZPrS0MefkNLdZUb7vQoMFoTTCEVy07KDfxAe62RtoW77rKXZX9Ph0Dq
iuBDvrb150QDMBNbzl2WG3pxjxNRGFJ0WlSLuamrf7cjehLKWh/ACqqMmW10uuejJC5mQ4OCHWA6
zmha6RLWNbq5YTtHfxGDH0/PJa6Y8Rg1CW1Z2gl+LO9IPIj2a0Uffg81uB9LNnNRDTW6iEGghUNN
MapWmCULskvnYZv3E8mKjDkrrzJS0hHWFC2U6BnOK3zc7twkzf3qrroRxnF0x4Fa+aFSEOLyKXKy
9Ql9UlNKfbrhcE66YNgi3dFX/bulmyoEBogxRiLNjpGJvkEkPB1/OTio6oLu5gBb5p1HOec3BoAK
2+Vm/Qmv5Ir7C2Ufw0l4ijp9duxDhLZfFP0pPshiqrca4TA3ndW1c7VlZ7itOwxVxhHAYn/fIh7T
NQfJBxIX0QGjezBionjCH7lw1QRrqLiX65VhaKIXaYY92Xt+JC+o3q2xs+7H4QZ7Tt/h3LR8qlBs
rQ4MAuRAkAadsa5xrAZ9mc0N0u7fmmitf6fzDI0RlY4HIXcICfNe1GFloKBhq81klNIya9ZTkqyf
bn4v0EXc45qfZQMdam+zo8DkWKbe1hipiXroG6BlK4yeJie9E2Xpcgm3WM8v209P26ayEAbjPyT6
kEnHN4KnLj3eXGdJzCDoP1YVoS8M9JP2nwnZd7TFkZrYCLB62TXjUq3nnSMnKMLFFNS8PAvmpWCl
ie0Ph7X0C0R1TQU0Ro/1LvsBfHBceMp/62c4TNOIUc0sRaiJHyv7wmmLYyrVOWgoYD/YNk9Pf4om
eAzyO8vHFFTBdF/kauJXnpSsnQKkHQKp2JlifroU8jCSwIApaeymGi+4NVQzxsVrJNRKSMdGKK1Y
1y8gHyibaOhVa5jpr+mxQiinyubcBPCmNM5rp9lLXU6YCLnpk1QLBjxRimet74Ei2HqzL0mQqqMa
X78Cebc3AX7oxsWBR0tlisI3JWqmkBqI560KYujFdwl8WfpXsNmkqnsHaw9i2m8nXaLR+TKYVDk2
a4CgWqq62N+4Q46jfPHUwRb+NAjysn852VQirAv1tGRBiG/ZNey4WXk78yDnuwt1mwVFQ35Ctccj
Gb0TLZKYWkLVFKYHUpLn1KjU+wsBlQZdx9WxcYM4Ypi8BLxtV4VlY2qKy5qMLuCCYxu8dsjmmMpN
mgWvjQnZGD9H3fTK7SdkAyyVqmvRpSc51m1p7B2RiB+nqKNt+UmHfZf8nDGnT5zaxUIZj+s7zHrZ
9dQWQLgSPUrawG5PcM6nEXevA2GMz4FyN7UzTk0Vkf5BOMVwcbnHi8iEYOwXMYrrfjq8CcJZzksH
2kJddpSM1pPuYMloBK/jZwEYtVTJNNgqok0rJua6yRwANp8ETb2ZtO0wFVkTIbGhfYd2jnXk2qBU
zp8zY8mig7mUAy91Sjj9gWxuXkqTv+R5hh9wkoacYyoicTYjhth78YXuTqGhpU3F55JnOZTITsHM
ZUAjPyawqt1C0b135DGOwtHQOLfsfpYWz0Fxw3xjj/lSINwC3y2k1FpPdocHEL5DhKXi/psgQeNL
QTU0NeXEy+1jaAeuSRkQ7tu9bReqq7rV16/BMhsFjeS3ExfrUMETJ3IAiDn6XeloouvWqczpCE9Z
QG7qQTyO/0VcfPScjJgf6vkiuI+/OnkdSr2m0L65Yc5UjpC5A+SEfHndpC6NmAqcVuLXysyKSQIq
skX7rcUC229V+/HpEOXyC+VUNgffDWP4UE1QAYkIJEdAQyBaAznrYeEt3Lfrv27KMe6mkfIq2+Ls
qrg2CUqB3AeKoyTJCqa1RW+adxm2tbJiby2VIq+bJmDRE3QEHSmc69jv7ArS5dzBx1v8H7wPTjyE
b4Rdp7DEs27hN2S0bU6gMmWO7xwVl7UARTcLI6R46jSsNQEOJu/26JGZNwQAIuJY3LVFtTAzlNP3
CehrukFZriIOC/b5UAeEafPkbeg/JOaUocWbx63JpLzgNElhcSRvn7LbIMpun2pGncDpIhhwRg2G
eDB4PAFavtxRQ2Tw0BR3ea8zJOn+fbRmYAj6phel0P7xnq2/7oATF6ZdHs1b5COleFlK+zDlN9w5
l42nJlNwFqcjEORI5oCnvY0SmtsCtRNkKMYLHwqE31/HBu1+N81BY8i4RNnqBthA9HbaE9jMcGI0
oymix7yKcKMQpNrd6Clu3ImWmUUnq32z9ix6IQicZBHa+2lNTMCqVIEnWiWUYlBFdV7+4flJ9kXP
g0UqAfDI75a/nnGq6g11ddbWz/B8mSwCgqsgovmDJWFOruWOL0NwRHP2/88I3AntzrZWxfknEYa+
XAa4NmgW+yy0MsK7KQ+xWvmodPj675qMBSNulrQmvddR45TED/Hfcg11biajrA55roehbQ4Kb+kz
QxzNTuV3Cf226e/FFIQ1D9aW4CZpJwONQI/X9+X4gVODAjGcTHNeIFZg+D6ugJZt/1w/KToUC0aK
12DE/ufspSI5VgBkK2DBYEG/3Nz7q2g387qQzujIyWMF0X9b63O6ALa/DZ6W0V1pojWUn6MUu0xS
b/JjbrvNt6qRY2Q/PV2ZP8rB7SZjJVIzNJ0ZCWAyZJ42kb4p1Hh5UzQjq8HHX0qH3X8CQY8oUNJg
5XlkeTWMExe44dzeSG7Mn3y4c6e0ATu3g23vE+cYsQqreGnOknGi5aP+lAJSftibmd6NPNpJNh9y
mAiSKvAPuSQYp2l5xpjWFjxPFtqS65rqNAjZa6EBz17oa1gWWpo77ucRc7jyGL+DyZ9HdQYUr/iQ
nRxZs75jQ5+xob/ozOERcW/UKWFnOp+l7jI0qJv4ZTpJLErC9f1ApPjUIES/8Wjpl6Te5IX/xNoj
OZV8+v/rU8uU0dRr5HDPOTTzcp8I9q0duHe0GWDjZS2Zrpw0lsMNdQD1nDsBMYE2AYjTOxDyS5l9
yQZ4En0pKLE6ssobazKDVJBkp4auXJLXx2z00bskaSvguMG3ww6+8l6cNrriyVf3HeFTujxgq6ld
Nuy6XaqEmdeofqMnRZm3aBXQGQZQitSSdu3QwZ+j7PjTzd0yRmF3n5v9L1M7G/khJ85KeEKMbzhY
zDvDwBGgVIj6eHew3iZ8EbDCKqI0Obkw2wfyNFq5SUBf9wHpZViR4v8C5blVO1J2j/vsjqQlhclH
jrkY4/3xcgyavQGTfxFsUoK9q01Kmfj/aghQbONsR06uj1tVq7V5c3mWYYU694cTJ5gLunf4VL19
32fLH1rNxFyjPfrbCF76a24NmV+ObXUaGZ6Z8NqiE26WYJU1RJy2tHS1WRy8Io9fAS5UJM5Sh0iK
avUxh6kkXXOd/uIeRqoyGKOZgZO26rxKBH/m3X+qRaUebLmnEk6CwcOn27PsTX8yAUu05lPqLwd+
ap5DYAci+QgNOV914ORCiWL4dN2t0S2zUW6ssyzVd78xoP0oNqBprk7SmXee/cs9xF1v8F31WXxV
uJNmVnmmxpewq5+ml3C05Rte4zSE/RyHKmVe/sbVK0YWzlG8MWsW9pmRd/ocEemuEr8jiGbnuEqY
vDAiBKN0HJN8ObNLoluBure/fBivaQkspZlvpnqoELikmBefs6Tjc4IjZtQ4zy6+A0nDuRhmA7Wp
Xg0MXrE735GJOekBGPrGtlm056T2Pjn5rqMLBlFlzMxV+cUPYqdMpfPVv51+Tf4aARLKyxbi0Zgo
qW8nd+ww945K29TFtSfHjZWyxYTZLpBQxzFSSM+n9cyV0GFVY4JlEHAQAKGeVejJqYTqGHciqaDx
xfW1ygwm2oSXzc17glvWbmUsHt7UqA7jq5O32mKKwLhEWfQ7ZeJ2vxqjWdjua63vXH62bz09Tj3K
KEKIX+lYtVCuxEzk23SQ1n/MlrcNxdbmlzO9OtkEq0d3mbMId8qKSrV8JHmcjsuh5h7bfytyskNj
ZB2XzXAgDJOLy3NHTuzGc9NBTES2xVXGT7Q7B0Eixy4XNER2XGl9AUK+JbTUQnQDjj8eBx9PLuZG
MGJu1wn5NWoXSwzBzy/J63MrdpviaDPSd18m0gPx71o+6Sk1/GrlzGheD5R4Iae1CgsNo8mlobiq
fMju5ZjVc4YfWhEUzLWrS0PAPznBs2qQEsusTdkV/ggantFS5qQgD+YWPNs+uFi3mgZa4zvnSyFw
9vKgMk7+4CrDrHpu+EMgAIxtBVLyM3Tpp8qadulNG2Pfq1uE6Y6sdIx36W2SSOxvVTNtpcKsE/68
BfzBJolIhbRuXGCQ1ZFstgIc5oSDa9hy0+QQJewVNXhCRzZhvRVEBgNuwZamU2PiJJ8L1WXkeEX/
KkK/9AwaQHeDkTT7XPdZB0WadFnhcxBv9q7c7/uqzKC7EB2pyo/MZukRPK93QUGq+GkIjFJ30qZM
mX136k65U0bly8/YcsmqxkjmwJMzHD82W/7me23DT9jlphH1uTaTaWzvEODEZu8jaOVK7D1ggdIV
Z9BWlKI1264FxWQKlOeXmSsPYMeINxv13IetEGMA3OsZbeGeFg0DcYkj1xl6OOkIddX0MqEQCiO7
jxPfGys5Pb/5dvI5wrnAFGZfVt4WcWyEIwdESTDkjmqakPkLAI1yjMyPUTXHagncwIdsXwPkMAlK
rxNhM4HKZ6WHoHKl/x9uZqgVTZ7i8BiukdznMQvmdXWI+N4FLVBj4Ds/5t8vAxvodE5pAYN/frX3
3XRnsO/+XefgE+Oi4C7nJXPEv+qtPfs3rPOhJB8XwMG+6JYYXHfG8Yi3o4Kvy+EZ9NAzGW+TmYi6
NOwsuLJqngGk6Ym8ns8Ybt7z3qOwpBV42iTaks/oHZ/LExq9yXfFss4aS3t5ayjyBkuMa9NZZatZ
mYbJ71oNKyyzk8NiO0VnvxVmUh1fh73Rx6C2D/V2vGHchMlvRibV7ZPv925p7LJ7W+2P/QwIPn5h
+fEVNZ6D8NMLk5Gu1d3N05lFR8yxJWkfJ9nAsX7B6KCfFvpb8alb8vO1kmk6rkJco2iBtcOIZIA1
nfkSdogxbZlA/DxXFd67ENPT7r+tpLI5pGc2fBFI7oHHnRmHSWBoyu+zHBK6k/O2DEs2agPitF77
Zo3DU4inIXacwZtbmXUkmxXqKKuNDTiSOcZSdkR5Mn3paGQ9F58OCSpgucwLLrTichs08lVJJucS
3JKLXLINDMRXmKsdhcUgeYDnNNcdJWj1VwbHtwYvUEunYVAFr1N3b7QdeJEVHp5bL3LMHNKvbhaF
iaHeGEviFi87VRzy1/EAvbALMtB6FldR9tvo/eKr07bUvHU+cH24ICYciP8eWuHev4U36TBXSGft
V/lGENJ9kUx9t/h/x2xTq4i31AadaHL6YRlnL8JOPHClp7FdwwqOSsz57JAiH9aE7OKsbInJ4071
68p+60EB7ONoXQlAYWOEZQlDt/+xZskmnFr9co1Hcfj2GZDzu7mvRNKGsXYqNCDC1G5J+SOPvxzS
vZUg38/UKCQliZwmJfSy2623Osj3xjl6cJ2fS0lFIFmJX66XycU2uQC138pjDXtTmZo9ZeTEHDhJ
SCN3n1p2VQVXkdJ8hqilApnEpOobJdocr4JFZFnqgH1AKsxi7yKYSQ3WVFrGwXxDA+Y8fVOe4iA6
/OQJLhbQD+9JNyJI1QJavSt6Y/HT0ksx9q+pHPFfdAknrrPXfvl/4NkKUARED9g6uy6CoAcQQTxL
W1uw0TLS2JDQO8Pu5jASuFZDQgMy0HLN3yTlC+tmTj4npRcufLxbbfSdEehyKvIO5D6jMAjTjRMj
XVpYBWSFqrGSmgs6Xj/9VeN4CmG0tonDHXYLQHU+vzDpfsxMoOqxTuVwjWS3lS/zjAY2N5Lr+Ayh
doph3NrLFyjzXc/wV5VA6ZA8lkJMNe8L/4dgmYQeNfytLjE73GGoMM3c8pVFhy5OgrcebC56OXhC
9hOx0vnlm4IOtcIYL14aKhLN9Sf8E9kBk3WuI7FLkNZNN04QxU5ZNv7kwzFXgYg7a6MbdjJJxLYh
pfqUC2iq+CI2lbOByQ3fkplzlzEcHhwCGzRJUcd/HCr6MdS6jBFZekgbRqf/+wOJT2n4hIMuO7Nj
ippFj5ujfm2/v/qajAa7NklFzi6OZv63Yruw43wKtlvNzXe+QSyya4AXpBC7QPW0n6ozg/eBqSWL
oVQQNBKVDy2EKP05tpNaAHUtDwAFrn9d225XvK/IBRIA403TWXNTxZkdJuBCKDFER6f7OOZzOhMI
+YEa07ZBUkIYXThNv8DVnNeKIafjoABCFiS2nHg0ZHS9qKTgfR4af03QU+C924/Qy5Rh+8XXRaUi
T8QoF6R1ZpCefDnhq1aB+thA2mnBR7kRMuzD+sq9I1whDuS9zx2xlAvqikdeoR4Pwy1OG083RxdG
i/Wm4YrUTdibGnoi2vE+RMACiLdE7zkacqzsMWGbPUNix2WeuPikuugCPWYkmUHmn2HKqR+UTq5Z
r91QR7NRJXs5LGFgxZxHkM6WvnYXw3llvPPmEfesMmlJSGyMvGHkKt6su8WZ4Xxe7d7gbE683TbS
5yZNm02JsqClZNdfaLNEs3j7ube5T++PMtfet1Lhl3uGwz/n3rwlQQlEbtNFwuo7Op4d7lj+08Mw
yr2Ab8S6czkhkjC0tb55NBBjN4iRcVZ9pUqsxaljAP478ItCGhQ2iN0xGNUZPwHMua75ahjVdmRW
RTFW7snNyNhOAnYi65Ubc4ZvxoSjv0hHg6jGlhjniJnXxuRZfiz77MGevP4mU3AxysbYZurDgkbc
wU8KCLsS0tTxLJgjCL6QoS1WofMC1KYGYlrt29Uy/gG+pJxofpo8QefGhi5IvWJxhTBcffJu/c2B
WRHWl/zldTH341Vn9/Jb6eshf54jlgrdm+PG9QZn9nkTd5NmMuT3RW8WPomnEd/5OUXACQsshwKm
/Eglb2jT0v+IyOIQOJAxbOpQuAr1kGM5DjpuaQaCTJXUwBIL3TJ1p9cQsWZYFS8MVhaHyO4T6iBv
BiHv+C38VesL7N3jkaRt77z5mI5fTLxCzWHfyq6gzLHKT04PsUj85bzrB3VHTkb5NYHJjNupcOCp
H2i2Y9TuTcrK09NYKH0kqTT/aMSOccUYOLUEvt41UEN+F3rJMDrH23SMqsKjApkNXNxg3GaSRkeA
sF7nYyxrNfEt7NRJzPhYZH8fAxhpiT+AWGSeIAiA37fPng5LWm8UV0fvNewQQmT07GlajUvesziv
3OdrIgVEJFIT7Z4ziueeaqBFcuF9/UK7QOyCP4H1u279LU5DTCyU2d6SiOhNdxxHR6UbF0ByCkZ9
OjQ9q2OhSxUxmsh/VtVoRaiDTvFTt31GaJijOet6yRtSb+tM+xGaDek3AYfeKjmkaQ3RNwnYDQAL
gxxW3vNa/jWGV+7P0OZD/omsn83vWldur/TrhreTdu38tKdW48LdffRjn78E2wwm82obmJ9LhStb
QzHy2EMixYTdbUwQLWvTAwAL0rGPbJIZ3IoYKHdjsj0HJmWOsLic3R2UHlvGpCGnmDEkGTrQpVFc
g3wy4u5w0AZPJFdd0JKG1MG0AnYSGd/4HY+P+xPwwkKK9cp+fmcx+YG+uttEBxMU+EGk7rup+/GH
VfX3++J0xUpEV4myO+g0H59OdcOaFr4NMFWcoS2tPcd0pruvbHCbJdV8FUeOas0XOTqaYvgeZK6e
EEJTj1fVDmrw8AMKjVnku8atMoXxLU7qpIxWfFXEW9a7Oci5Ntbs6cgIYnL98JqnokrlFo3ZYG0u
260XpL7sEnDTHJ6UdY5PH8Q84k5WjWgnrHMxfFsDOieGnncCwcDZPjK7pCfz37ow+1Z9fsGZ9TLA
gzB+0wdWt0w0eASIf02DCyF9wc9Zci5eJSYZ/yG8gerBQw5qM6yuOsFATRbyZQ7T/UlABeh4MOi1
k2UwwMfQf8COw+eDT9mXPiIh4kH2q5iEZU0v2IBrC6SjmER/Ltksny7eCkG9k3xyGnPc/tB6W53y
UccOMkxGmzwVwNrNUOEthNJbCY+ON2GqIkJxN4L9NskK4cZaYe8E7cuUDHmaQ5LHfoCuUtyrfvkD
afewBiilQ0wERnlMWowLFhcGDfIn/70ci9cxRLD2GecRm0RZtdruser6KsT1iRDdAQlWFTkAC82y
OXhDSpkNOkYAwI+3iAQDGZwI2vMuUmVsFjzJ3FBgR5gfyLDLKWpoKAGH3gChwMPGl24icHrG8yeo
oGRuyYhsCsTaseaQSNANqTeiuzKzRd1tv7xkJOe5hb+TRySsqJRl67vcyGfHEnoBF9I0ONrV50/6
btq7eaWJQgoCzt3kQ60ajeZjkTY/WMG0fsMajrpEZct5ZG3tw4trf9JiuzqdUPbeQenA6Lzf5Hpk
Ec1OKBiPee9O0wodLW4sevb1pUATwQ/hmbWoQByVfM59MGcYw8p+hgsYZscFgF9BIrShZxmSJ0Lu
WE9fheKUFNj0RtJV4AufKcQ/LN11d+ZATVkMeCwqlkCn7jYD0iuoyVQHCSL3w+MCbAXx1iLomXmq
/qQrT27n5oNRzs8uOz0qO5HMIhz6MRS37U0NFWt49fx7HY31fwarHanZx2KxmL8ybKPKw9kjWnPy
I4BAuxg6Fvu9dc0cgcArOuZWcFXzvZAQzxES6wNiXuC20IlA2P3ieHp0aNpyhUcH33l1szqlQ4I3
ahwencE9voZmR7Aamce7QSPg/4rgS0xSTIc87pMqqLgH0MAyl9kzgNE4BxcMcR7m7Dm40FlLRXbY
jOkdY4TiW/7Lur42l7uQZtKNipDJ4ZWPvMQmIr0Y3zcOjco56KG6Inn2u3Ga1NPR0lcrJsWR5y8C
i94XD28xVUngL5MKVOqYKKnOUu7hL7JDJWtAiuPsJTfAlGnKD7u1p9OXJNLaukOl/bEyph3I+vrc
4Ag858B+p1MqT39qa68eM6ZBsLQVjeWeEEEWrV2Mmc2MoZ2j5nmb6ByItlrdwxW7dMI8BTCBVPzA
e7jMQGZhVT7U9GB+7vSeS98wZkSqSzoYVFA9J3mRRzxdNHR0Fo26PwS5TXqJEn8Nv5oPnmcRpZDW
xpoQX8r3/UYSfwjNNy8yt3EZzwGNodyBVhhGUlXP0fGL4CL+VzgYdvEVHtsq81GjYa/jG5nxDDHR
zdJpk94IZzi+wAKTkxd774yPpffGH6l5yJGd8Ygaan83W8JaxJAQu0yzOwK5vDD5SWPiqsbWNnei
hRIt0EDc+lfytKaPayh01y9WVoXmXyxP+C0MYyocUEMpmaFqpsXgnWPA4rOLs92J5Nwz1vTOw0kx
mDoXDZMTnU/G3rcDfAVzoEDRUXR336wjdVInWepNMkeoxvWIHexO5P/AWBnauW+TR22XdD25pCFP
4b4RgnBsfETZpqXuCJgvvO+2pNn0c9akj4kvv9+v/rICnRHwlPH3fKXeHexWgicmcLvfGaykFuDt
bwAl9MpN1FYg3dhF1bECm0oGE1zYwkAKFotC2VuXcA5+ttPPPLqBb5nnVpXdpG4klaw6HTerx05y
RNH++aYdydSQyZewVJLAfwZNvjQyP5LNMpsApIpdCBX1jfoqcTy52IcBDVFvmI4VfcsskqsIvxy5
PdEgtll6PC6O/Dt11Z6hYB9QReKimgVtJ1pYQfOZ/rzXqJjVGFbzLJarp/PJU2ZwMCOblKzm9U3r
Nnx6D2UOCLXzYYis6DzumfOP56VjtjAqGFoFJ8VP6l3zR2OcMAC7drp51Y9dO1nzi5gv7vQB2c7c
mrwS+bsGxtk8L3QdJfwuUlGNT8wzx1JTgzVu1pSJ/6iN37Hv3J0WQgX5b6AuI9tnOlh5XssIpf+v
y/cLZL48Ki1hYUrigxq+oFY+tWdqHpzuHuzE8nHE3C8rEhmbthHpLhlHDtq3zahrM9wDll8YrAqR
Rd4NsvwozbgbILT7NbSoZLuPbzSQfMxcvLmGLKb+L5XJ5zwSYJij6ii1LClZkSQP2f5TzAgdDUK8
0/2nA888uhtdjagHb7rV57KMeLkhLaHqiMT8hSBF+bDNY/XqG2qlQLeinMI9Oj+LQE5aN4pGrLQq
VPi64+YvMkSNbUKVHJfiVE7Y91KJcXwFh0cTmdDGZZMLKfW10Pf3VdW9i5BFQQ7TLBszSzFmCthQ
hyrCRI+rkuWuVUcQltIDGuhsTp0LJGnoyXQlbp07bm/BG6DajvXbKG/+ZknWWZQPZoe8MjJ8zg2Q
ECI/abOjxY30+dBcqGJJneNDVJ8Iz/mEdsUAVTtFGa12g0ArJFzXSnlT0AjmN+lWrqcYliwW+/lC
3J7TZnduPj16pnGmVntcc7zcvVaLmZ3CK9Mw67TwBKPm7jGqa3FMEp+kLfQfwPDIjxwbCI0/xHl7
qUO372r8abDVMXnZUos3x8t1P482S1i/702SXdPLvqL0QMvwwtKFR5rUG22f+a7+Ks4YHlUqammh
+0QT5UxE+SMRctRwfNIgltg2IVSVzn7ZKGfiqehjB2j26XsBcqbFwa76jOqsufJX2mhImr3XNDg5
f9RC7XfY/1NhN3ZTqJawCVmy48MXsZq4rVI+bZzQ8efMYU0sW65DCfYHEs3yny783TAqpFuk4DmF
KUC83vg2nlgqifAImKgPC0VTIvYP5rAZTOnna+1xT1KYomsR9tSU6KYZtCKiQXm01DVeP3RqmHVT
oXBWilsXeEPK/x2e9DY6FsO8Mqgz6Blvgfg2OfclOVpIL2/joBHjQorreZ0lUA8YHUEHII8fohVD
7q/94WEYi15pcB4CSXsFOUQpeu9xFyv9evA+Cp4oozNdTIWEZjOmMAL1t0jcgzZ7o1CZl9A4MR5a
ASMQPOpI0eRL41a6EmjaaUHlz82kKWuioSV6X8/i+Tw3ZG6YBSqKF/RoocS+wjv5POoEQ9SBp+fB
WGa98oCcfE+b+mgooaQU3x65dndRQe4EN56yDqRfZzoeQTccRK9V+7U1Amg0T//AQ4mM4rKEJF7S
vjZAp7geoKPpZjF0doZ2MynBkOsvXbNjirGvY2SNUNG0i1g9ryM1/aE7r+bi8HgbJzOzuxNJ6bm/
ZTdESi0thQBVhkKeTpL9+pAI2zi8b1qd/M8LLRHbly6x65ccFnE6k9pdJTtNfy7HhhBAeHPAryf7
XlJHKyb5RB3qh8OhpMLPoi4ZUrQgxmosKlLQcT5G2gBH7es4AIX2hW2ZGMpAGIGmGmUN9Ec73Tpi
9+yph2oWNF/haxZzNu7f9GnW0/3wB8+O5o2pIiXEaquZohB11r1Npbt7ApbtiEV4rvJIiiwYT/U8
AVrAnvk/lonYezGIuCyravUEwceSSi0yz65QRxQk7aKZfe9Y/JetBylBNgYjMNgcE0lq+bXuk2xk
GpIMiFioCYhU4/M7b09XuHZ4fDOLjF+mAkz76TCwOIPReq/6eyjf/U484I+gddQ6+Z/s6Hytwk2k
3wYP7A6vWmM0ZrDDaDP4QAh+2gSGGOsIN9/eaurlhzAk3qno2bLPBfXZUkr8dPYtelpgTOxjWRSZ
qvVOJ7x52nvGvKQyxGxQkj7KxBZt0nZd2MYr5npnTwSJ6gcoKGzzheSSqBf/6KhMT+AvpUv+P0oT
SI4vSGjqQHyZqIrFx27gkQaloPCg8F/n5yc72wmp7BUMyHeEBSy5y5VTX40VXtakRuLRG5RcUqXE
TVUEr/aS8kho+e/Rmc9qo+tksamY49XAM7A3IcNb9kSBe3lfOWRiUaxVg+yIdlu5FxOmuMvkOKlG
8N6ZsaMQION+yj0Cp4eYPGHKPlZCBRPolXeiAL9z4WJiYnIQLAH0N8Z+vCIeqm4RZjiVLrbRG0m9
jVXwstd7nwrrsAHWVc30GWalhHurjUawPNEYJPcb32anYtFQa9O/+pP8w6mMcI6sa73CsAdd7KYu
YKKXFOK43ou+eMQFyscmWgUXXoj6ZYFhFT2o49ATuy4q1vbdGFRRcsn6oUK7jBGx2QEOR0Qzk05g
+bONlEL5PdDddCRJRv6zmU81sF6JZF2MP9NO7gpdytk4HR4xAGFJJZZkfn57hh8deL25K0kfQ0K2
x/NHl+EicQLfFTcibYCp+M/jm5prt60ksJWRr0YAcRDKRakN8Ufc9zofERuVmTW+oYdVLA7gpsmT
neTVaOPMXDb0+eySVo6Q+RtQhjz7x6562dvHtXxaako59oU99Gxji5ywSv+AGQiOrj6CrbKzccEC
1Yz1x7vNBWKAy3OQuLUDjMZ6soFFrpKJsnLqrxcjheph5WiyJLJhF+OwV1Zq/BIDd9nvNXd7TBxw
5nLICvnWs24epT8OFarygxswcTPHYNngJnaU9lxawTqistaoCoQnyz39c1leKyO5Yi96EHKsVBNK
avUYnhZ3t9+M2DPqi1wGOiMxheIyNqpU5t29AEDrdaPlkCxEIKPFiZbBZdT+QZiqMD2nlERt1YfW
F9yOSpxgQYHTUXdSM8mnTE+SYWbH9LSa8hQudGodYLT4nzwZTRqcQE00cg3T7V65saiflzjmbB7V
CfM7o/3hF1V80oWroLeHLEiDXXbRLPBCOxLCoWoYZ2AQfCLFpXeCpvUvypRFzhjkzXbtaOv7w7ep
wZ+5qXHrcOSIGXbK09lpjFyaY1mlcC3NTNmZXgGt74SEm2yHb3h59N8bidxk8SR5e+ZRo37F7xCT
8P3Q2iznoaEsoQnlXy5T6wzCcww+R63IJnnnaK+9OKXMI4lAgSxyzGy3KmdsIJ9phmSghNFah48q
849FJIONo19zPzM8QKrZPXyY4pANIMtQ1c2cSUJ4U/cGbt/w2j+MUrXf0BC2sf2FGG4JhAX+rzm4
bvIWOiUOPLDf2xkTeANiNYOr8AxFbSJmrOrcYl00FN9dRgecT7MXjHkpIg4rzxoD/qzRgyGKRBCu
dH94vb0OO4iO830hB8kU5Dd7T0eCWFm9P7FNitEBVqRxNEuihM/YpNOi25MSq1uO3YkRSJnHr64k
5TwG47fDi6sglv0/NGN6DatdEJRfvklHrI7JJsyioSOWgXVoTkC4M7BHVQ7goQ10vbko6pvGLcL2
tZLwKdWRIy3QM81tG5uxsOPCFfOhtXOCwwzw+LGfntdbcLW2EXSLHEGjVJAzJtbjlaIKXYyYdnv/
/EEdxD+zx4dOmai297zJ0mslpFFQ0mzdq4f0XZIEYA27ESdoDQKosvM9GMbVD9XSl+HPicpgFZI3
W3lfhm79QHa3vii0gdkZ81/8TNT1eBkw1kObSC466fqzUZtIWph67W3CGmtI130Ztj4xg6ghIG3j
9trMGkDb8YBoDuQ2XkNI1V3osQLZeFb+/Gu6hMOKn6PkmFfZAhLdsK3pO/iGlvhrWeyPWOMXA26o
lq8JLwp0XdhfsPw/1YEGmvm6wd+DxMEkPcCcJ2qu6hnSaiNLarHYtOn5b0Jou2MWmZtgt1vLIWU1
IURL5+uee0UNeANIUb4F4zY+Od6NmRqfUrZpKuu4k2otbYMi7OMsDDyPUkyLEGMHpN6pyJaTSKCo
tQu/5dtSJ/HgZjizl5tdW4XzsAyH2Si8/5NLh4o9mGjg+n/++VFeTMqDDfIAGswwX5aPtKQ4ff/q
e07XEzf8Jc4nI1o8S0Cj6eNUBZbhz7uYXN5Zd2XaFZms+CrIHQJq6NczYZ/hJeYA34UEaJO4AKHJ
v4WDENWdCXgq49Vp1uww8DEXFRPkQAC29+vh28gfZaha2ElW2oHxffAmfDVJECYowcHzS66OjNiI
jKo/1DRjHX2sTrEVjy7pzLYRJFiLEEc8tZaKwas9bOmJ0mJji395J41mHTbzdhkR2yGVfO+kcUzo
h24fze5I7ry9/nN+amyp8y+YSMc8TVF4TVvVWvwzifGCYI9d3pJd2R/xgtiDZeoplBV1ucyy8G28
nz/WTX15vbk/8tglh3xm86yUz1NkdlOvRKZm+++t7N9vf3jjY8eEp/VXD3xTG3mf0De0phuBe1UL
z2AVv54Ut3P8o1uxA09xD4HDiONxiVa8nyf0j3sRdLb734tmUIzWOcG2f01LgtExlVESk5aFAPk5
f/SXFtfvhSTyiXNggNTfZtyGTyO14eFKITJGKpBMB5JjVaraXQl945JMcydEHptogP2cEfJdA7Mc
lFpj0+VAwQ/c3WJiodgaIbW/R3TeguVV6vB99iyhWQAKScNAgyjc/nVuzOmmhgGqBnJOU0fCIBTG
WnqgWpPoUwOBo7MSpbmR7Xlj+7ymjoSJABRF7/LIozEdvaMi9wnithQHEfmysHf06X4pZDBQ9K7W
0xbbqN5tZbEy23JUQER9lIAPcxGQV0vvIYCIXcKcec/Xze4QjzdPdJPeH9DNIelWctzUjFrlTuR2
YjX9ldNQozroVismFaIeIuypfRnS/I9BhQDvWK9E8QXL2/An1Uc7GGn3Aanjv4KY8vj5pbtaVbpR
SDXeyYOx6Ean3Io74ixlsFTJM+Z+00iqiFHmTvoVLmMiCBLXLQiw3DqbxAMfv2yHDtvQp2VrhOi6
Lm0Oc+8o0f0xv9zxr6YrN4WXXhYfJsZPhayoHt2wil4CQAqpOQnuEQcMjOez5UY3RYrvLwcpmh1j
s34LaIp+ozHKWL1G+DTKIdrJEdAxbKv3REEfFx+ZNBTme+Xbg87Gv09IFB7hUa9ppSzEohUHgcGZ
eBAMlONxdHD3bEXwpa2Tm6WNhb7jQ46g5fcfnQVce3c29LuOf1mDq9q6QSXiGuNSK0f0bpWGowPV
QYquMyajfmdpZK3cDzw0gCFN6a5bZQxTgRt201/AXkFL2SR2ZMtm8ZLj56r5qDAyYsw8TbJngE2A
0gKP3mI3BRSnmWeDHOLNhpQzLykkvww1P3KHtun/e9EANdJXnSCO7x9t267Y6GaHg7DHLFVoLWZZ
pXVdN2TYESzZzfuXoiwAA6+FeavLVjkzFaybxz8uwY14oFn2KBKmVX9RBHM0PzhsDWXrSJ6g6AZS
fLL5Km0IYynmAj//vXK5OYZ+Hs1ytJy3dX4uO1TZHPSEf/gn2cY2BXZAwNi1gzQySXc0eS8x8Ykn
sIOGd/jvnshs4d9BwlOnC4oC2ODD66H5Uh1ugZfkhM6BepkHjcMGztqIvcsH4bOGJMk8F5ohpqcE
+p/hbveDpu5bQpUw9LP3sj0GamJ8UAwajdZKOdZlHBpsf7R7f9p8IyhXLIUCdLB6xiGY65xepTOY
IGUlY59WIA3xgiNj/DWIYdCKwW6FjUdBBqjuia1D4tq71oxnCgLCthJ5qJYN/Tz9lRXoXY9SCcTL
rvOPp7R4we4DdAC27xmfa7YQwH2l5tom1lg7xL6Gr8QRTUqMwXi2vYo6lvfeeG5X4jt2FX+6jxey
/RBSStrRV2DXsptjSErYAVdlEVYXNPruDbDMT4FYUeE4vOOs4KLV3afb3ITonvPpETy9wgI8hlAL
M5hgbbjRNqUrNNv4qnMHVcMdekD5LlUKl/Y/DExA1FbeIzaTX8EPLeEoiBSRZZKcWMTBefYsI3t6
qLkcG19vPrxh/RITODb89nMFfTB/UI6iGhwxTE6qqZrabBflrDo229TBBLRV+KmarsVYqx6UYVK2
p9fKZQB+NzXBg+kIyeqNuftL2keFUiJdyyuEVpmW3iqfk3sXbXySW+GJua/07NjHsxh+7wm6PnQh
5Yk04PP+rJx7oG1TCDg8JBpwtTkbNL5rZ38vF6vIaIg29E+G21DV8fOxjIV/v6nSe0n6QskyIHLJ
dx/0R/9WHXA3uruyTMrATB43JJCARght1u/Jcj3lHJZMAmPCRmpunwqq+Tkk3Vbsu+o7VRiMstDo
nGQuwN2xRpU2fmtxnyhMC7i9azBjUCB3+83ATl6ZaQhZllSvFm1TMZ5UUf26txoX+v9B33hLbxzY
wo2jjjuMrHWWEdZbqy0nSlxZIaI7i6Zaa2H5md7Z03/1lQHMiOYRIkf9KwsPp47XsLRb35U9pOi2
pYwVfWLKIL/13EZIO3/LNcK4FAsj426GtgGhkTDknLhQqJiOvB6cd7nWtc+vyTu/i6OeDXIvDHvA
ClrCn7XJ/rJSi1kN5OMwJ7RqQwAH283K7ODxKfmoN9PWyJuIQIWunbx9lAQvHv3n6IdEHdOK7lvU
6Wa0GQ+iQLHKoDMdWPtjgy4IBe6uVHndtpJ/Ts4EFCj9IC7AD8qr1YVyEKdMmblHY4hdR3hFoT5P
3ZlfWntYtb9g30aWlzmB60ubqWy2BLcGztajgOhlsZ7IJ86CkdbrPbfRvviUYq3XimwhZ8f+XlWF
mSf3DiRN6ZQL83cUFBSsMZM1oPbZgeYF8i1bktMUVolVXb1wMsmZlopOxrCiIIGkSa8rJPh3ZC8E
eQUk+ompc7FutJpqnx9TorePMTrBsaCoR83KhR4/1HQeAfshc4e9cjD6qQbw8twLAaN4btZZhXWs
iCIrXJuEVQM+4InCmECh9Aw1Vo9pERgt+GXlpyDifz84dsXgt3FFi15QGgQXqSwGYmwkEdkBYfM8
5NthEZCkv8HTTLj4j7ea+pyir5kWTsqcwX5JRJeKX6pyFqbymK9cRa7Oz+dJ8ENChbPAHe+wfVEC
XKuE/+WFotPdi2z1Qj40CEQpoRm6iJr7la7Poer0Tkk+pdKVvdfCFt5ZUCRoYZEiJ7CmDa1MaKrs
3O6dBaMjjSdWS+uw528Zo9R4DUwdx6mobrWVvE9SJ5WrVFsNzOSNl1P1ePIuQyYWynNEnntafPjv
fG71T2oFSHeV34i/sF2/g8b5AtszjwmSFPgAJ2hN4VpnvjV2rg4yfT+9GAE94DX2SRx2ib7PLo8H
/VaTLewIhqZ9Tbje3cJO6BwMefUPErVtN8CFAjqYswhXWCTxsLXracPz6o4Egw80Her/KdEnxBQO
/DzmALFnWK7lvbhXMaTEut3KcbeWqF60iGyUbTPMW+q7JMTrBmxZVBxbxeROSCVxaVoBVOx5RFtv
6gUBzzhZBEjIY5nIQgKvXkAIpT6fHSqA49QOde4Osmj0Qlnb4OuGZO2NmyDM/+0B2cUxNrzWKgkr
Aqzeb7pqUHaLktBHVZtrMWrJf2AE8HEEcXPjIhXaqup+mo8LBcesA3b5C+4x4UdMRtWrKZ86es4W
DqCrtLI6dabMb3yqjcXbuyHVi90mOaP1CDJJB/63KZP1qKFNN9r22goHiLc/K3bYAFhdr37YTbZQ
3IBZIFfphZFUY5tbNqObM8kbNL4CGwhDlpRbvXowdv3p+hr8DeR/jcETg89QgCwSxe3wJUB/NjTe
RLG+K/uJiVri5V9JSDCMwIthp0LmekS6yO05Pq1IMQstrj8Y+PNJoxkr9OKxZki0uUx8UZZK04Hy
YQEXe8QqbmXa0jwnFfvSgxjpEJj3w2LFfvIOpNWx6/tKfggx6FCBdkXIrtv7KBMs3pQ8nE+qouG1
y8Oc25WYYibWBU41Ll66Hdj5bN0yBDe1am4txIza61TvrL7N9GQIkTxoxKcf/hzZq0DaPGW7R87Y
/5rYDq/KKqbQO8GAa/1yHz9/WR+GrjpBrcHoMoZlT/uOqePBBjrTUbsMaPdpsSssEAxJOCSb5nSJ
Sd12aD5p2N0oEIAG7APMSQ960Hre9QoHi0luz2N7mYd70znQX6UtXKktI6eo6tDRR1rjQpHR24oj
q1oUhXm6Yp9dwF7oOWIlFVsHkckrpUHhLbV6uLxw9zYOKtqLykrrBTAujFdOwIqvQdyVO5oH3MvZ
3n037QqwtqXvrqqujTr1v4N1B0YKpJ4fvoYKjm+P7T+IfzPF19QYltidjrqWK/xPGvxBbwcE3iX8
TOm2nACgt/qAdWqFwkwuhD4LZ1+pH3CRS3x9tQo5lF+iau39ycJ6h5/gFoKl54dtiDORwT6EANv0
2KTIahktrsuseMJri1+e+UlsJHI4vzUuVe5OuK8ll4k5eD+gKIeR4oM4M4ju3jx/KvQvU+bDG9dO
zzvPQGCkPotqilwFLGOR43KnnT5s/txWnC3CYHBJVv1dz+lOzDl6w3qe4vd+oku36poR+PWdtdKE
rDhFTxw74yHIyCwSyA2AdoIowtMo08j4aEkjUEVf8J8vueD570Sy3E0Ua28hsLjhfc6R57cUFssL
i077wFkTQo/2ddrLK0QHUnpSV6rDpXxGIS/wUW45/fV7AeRloh6V9RAIUCH/DArztpEVVFf4bF1k
6Fj2BRnoj7QUlqV8JM5zffRVPEsga7sed4WJX5FqJNu2R0urgcX1neETLgCbP879W91x4ammNuSF
MGSPVYP00vjF/EtFtXFLAqeWVR9PfoiJL3wnaXFYkR0wy8sr0TzOjVcoxkscQ/uDblF2AyYCCZNF
ke0ComC0HYWNG+U5xX4V26jRU38KJACNPCAJLpt/Kv8OdjBbgjYH3HmucIvRF7roum4la0SmNDJI
LveHlNnV4biKMYLHeZtktWDkMHFAHmJyYDkyo4gQMNkBLn4QDCnCkYopvOwFfh3qHQKss42CjWGI
LeybAAqQ5dRkO/m6iD3Hd6qemZWEw9UwqegJcCE7xDgRtUPCGONjCcPOE1ah9GOxBOWtVHqvEHT3
PGMnz/G+qdcMuAGj/IDYQq1SZsvDu+fR3MZFigvcJNEJNUp/2yp/0V/2zOz5sHhLAke26K/7qLoD
IQigIMVINuPK2pws/9p/+wtFfxr4cDUSTAMai8V8x7IfelCcsl2XwhEFib9AO3K5O2WSrEq0b67D
HHYMfN8r7p/K/6bIKaDYkrOgoElhB7whfRpkra8dxCtcRGO2R7a9xnVs2H73W9Zuips1myaAvgf9
/zfi7ehyoNmzLwq5KzAiuSLXtcQ+hX8t4JsVY0LB1RDBH/h6GHY0+zXDX5Z3xnZc2mA/ft2d9dNW
SYK7lHCom67a5epnDevbNDpJQAjAEVFKkQ1jBIdiJhBi1IxxmdoGGRJYsYcWVAVTPq+BbWBfLXEb
jKSfIskKyNX7jjTsNaiF4w+s/CE4JBjUVtcazJk/4GJpNwZwTuIHrmyQIUZoSrzQgg/kqW/XcKYw
RhBtbOQjnQvC+qAjWyuovTB5V/mtarnZXx0XIZ95+GXEG++l4eQvZggSGP45IxJdGDwPp3pD1Ab8
V3m568srQ1rY8469cfE5CaGKEeKSjTKtObghDpcro6PS62WVFPFnEZJ506YNYGRo2HMzwXEWYPvj
dnGhFlhspMwVVPY8rkkJBo5dk5bJC/7Q/RAktQpPppoJgEfRHz8PdC97AgPkNt1o2374/q+A15P2
CYD1dTxU/u2BYb+oH6O6JdKB2dvyDuu1p9+c1zCQhCgmYfiTEuRkzGNj2G4hvibwyJof1A+FqvPx
frRJSfz2kG6jkIGXzFL5JcTo89PRY8uw21e0UgV/u7P7gcfX6ys8yW+Vy1fk6uqgH3/x9EVNV+g1
4vHoiU9r+g8zcxOoq36de+SbgKgmiJLCoQJl77x4JorVlN4A9e/blOwq/siu1E+deX8qyoZlZVGO
k9QWw4svbNCskyKQ/y3TBugLAmMqyfhovo5WiD8rizrjuUh6aQ6+nVC6tS8T3ZoLZC+rJOBckDnp
60Ju8D+idOHOMs3wRF1X8vr2/ZRDnsm/ijFJ9y02YPerHFf7s9qa4BCiGaswDeaJLB/2jZxOuW/c
tYn9VnVl39QYFDPePMr7BhpCK0/7mGhvugmJay23aT0stCzEwn5iSIAP4xl9uiNB3y0af8ZA4e5e
ieJ4ldWS1sjlrXVe1uJ7i4Yb3lMNYXDO533KfkJtgH4rh2r4qDmjXmAkuFLKW0JgXhr/nRDcjxoq
9PkiqevPfzlJkUW6Nm99kDf7yYiwIFiftIy5M25M5UBWyDjO7KH6tUWtZgvM9+ERI6BVkr/03iRq
axu9kLKY/K4GbcxqTB/WpD8o4stpYHf4c6UnkBUhPkfe3qUSbBWTJahCnfKkW7tELJ60t+mUsN0Z
jk/KIHphWanEzfooiryBCNYGAXF39I44r+6/VMK9AWBfYCO3sWb9UzEuq62gU/5ek2ZGxlQwLdkH
IlhYAFi5/JthwoPz7RR4d7pJv0hPRE8IuzekGHrjWLQNPxezm6nCM+TDiWrXotuSWHL6j0L5IVhV
cKMXkquDNCIDwZeKAndnYPbOXN3ovXJYuTl07EYcjxZ9gDMbdTrTx74a5lebVNEZcA220FGDGX68
Ze++ntZLVxk23mD7i5l9FzSKpy3+qZ85lEAQ1T78EHRT8B8Z0WHYh+JI3Rsj/WlmfOBbF+oagRu+
nLkRbNvEhqV7GGGockyciRAbD1m+QgvgiOL9BRD0MbIStUx4hGKGY839HMNVUKIrNCeszFFz2KUy
pXQeTCS4lbg/WAFf7+LLTCYJW5p9bh++keB5MCuor1nReGpBvP1tOd8zJ80FIPHL3IYNQiHG+Hsm
2uM7Hs8A++2+2pxdnDS36kr8DPxMeX12F4J7EBPoQaQLAw4esL2/ZIcdn5ApcylANumZ7PYqnRdX
U43XNx23Vjbp9/c8kv0Y2HIiM8lCYcjLkBREkcFnq4sFeZ7LzPeWhT3PyzivqfTiPs1SgEIFSXqR
Gfy7gu5x2FUsGDoeCe3/omJ0ylmCtyMVMPQHDFxUN9e5ihYgcAeu4/o1BtYToiSlst89OYj6p6FV
kMXX3AQow8CF7DLbq6VSpIPtcOpLY59JNzEv8kHQ7IamfD9+0j8kdph6ph00wiYysjGylM+x5C/S
DAZO6yqipt/wfnRvg4pM+dZYPz4XDJUNTPq6PhYaxGy9UJSN11Bsh+mQa3wyI5fdsDAMDk5BFVVd
tX0h5SoBvSJeiHPBK5ngCNm6DgHJVgTy43eWDvsMXdC950UmhTUkqRmDNNoPA7pGFsusHp1WjbJl
EtW/ekREmTbDwgc7dIoJlfnSR+eT25DFbDPOqNKMmg4l11jz3iaBPvVlUK8pjidaKvyGBQn3+wvB
e9ilPgIq72mdJ/UmsuVi52yRfOLaajTI9QfROTOP23PHXL7ldObJRZmQR4y2OxbjQ0nLxSX7rmTz
UaPLtvWErwSp9T8ENfwRjpaTyq84CvQsLB/uW2BbrOD5KiM0oIhdB+rXfkLx1g2LX8DmeRm3YGNt
m5vjYUqyypfZ8CAnVeaiX1WY9AbqzHZsNozguyHNUVVOHtmFdSltkr00iqdhkrvvAS9AxgoJ0yuX
HEZ5HR683LaBWplBqRRs6amBHQQ7ogVYE77pUr6lqx/lPHJ6rnlCKrY5dzU4X+iiWCcLFBxlaidQ
1DfijVX7FhpIZs20n7x5epJH6hS4H8aSiuX10Mw3KX6YFunkfIOJ78aUGHeqgEKobHVsGGTP0Twy
FJh8MN0uv/I9M2iG4zPRZnjUsMcnWsRKXVs+70G8/eu/syH25RyMzRWsO5VGV6LdaPg04vevhVz3
7EVt2WPVH7VXhCJbHDrxxc/GFtUdSFrvGvleuIdIIc/RHobaKNSUks58Rn4hKXwc8A9P8bxb8s+S
lrlHoHDmr7TUBc2hMmJmxFRsnjvoT9DtNxIDhSEKfzlW685nQZ3gT7BrJyBvDMzPCMSoS2hYY6U/
cS0TXSXQComTcoy8tEPboXwfvxYS0OAzdyW3mcGbZvwXXRFNYu6Eik9i2fOUugGKSyY7oimpLelB
LG1xKZhGM/ybyHhlBRFi2ucm0adtrHMnv4YeTAdVRFwdLoMikkDOO5tFQXK+MD4XrNfpGeVhvxa/
DrJamSV9RLpiqWM/o0/cQOxNbTsBJ+JG+eIXW4qjfPBj7xVMPpWFeD0QD/M6DC6leR6jU6YS3zGj
2A40k04js0rRjPCscY6K2NAtzdQg8U5uT1t38W8jvC8s0F+T78RIYJXGYnpGtb6j+gy1HSv40Pt2
T8f7Sqb7SiCjOc3VdkKP96w2gM4TSsKTW4z9UvkjZecHr8LfOAPmvGBTBfbaH2qcMWsDbZ786kja
cXxEG0uQym8ryI3Z6ejTmesJUJyDVOe+yyI8uIMFh7SgQPfGJDv8oCbS7RfwwUAeUC07yH/ifnOT
aiFzWJ+qAzEc+fiFOLzSiZaat/qxq/vj/gdRKvwip4d98w2+XxAd2c6G3lN516msC9o0kEO5k7WM
LmehVnAwmJ6zaO1yYAHXThuP3tF5HghSislp4131+MxGygaX+xwR4JdxZfByYiutDuxE7f8KWox0
mFzhMD5bOM+Yq3UHa1PLNz/acTZuRLtQpxnweLXj+gGz1osO4issBCkQL5oImLwnkihR7rVoMc2J
M2joL3pPeq5J8SLV+M8RHCLls9v9EDPLm57OcU09CmOHqxLKhdrtME6Nj0h2+TxzNPKnaltSIAC9
LlJTpp8yngr+mfziiRjqTgc95viL2foTEDwWV4xKzVQerljcaXuqZBhzOs0eiQsonjMsjQEw8FlA
yuSiAQ3L5UtJn3e5zAZbXMLbEXtb1305JdpcAHcRhfveGJ6T69MA6ckFqnsN0Mt04AyMZxHtCNvX
/r2MmPYJC+3Ary8u6xqytGPBCREQvdrWAASMQKLupBiCp5hf5uSqzJ7K+ltMgkCblMkGzPlImgcd
tqCjSkOu7KxSPzjKfnpMkzvbMJWNB0OCuEheO4Oq5Zjywow8ZXf8er8Y/pa4Z8YyVBngrh3qK0RN
hhgHlUWQ/k9WF3jJjNnmDl2HRJsQaTpUXm8WDpHlxebXmiAhlaQOoXdZS2uY6xyYpcNcbVl9T1ub
yIWzkdHgi1Fo4fEYPwUjtMkkDDRTg0h8HX7d4XIZ5HhMnykeB5Q2fEMdYhgcti+pntx/C8RHgz0c
Azm/rrv9vpPOhlywPzuLLAyxFFAD9FLbpsCTrkLsmC+KpipNuaM2i3BlEHFTTbxLbKneEEte+1y8
pYcfOJ2ZsCDdrxAv+72t5MI/kahB22XZhaB5offYSWOkZKP2dq94/WC4ou/CbyvFas2AnI9KHPdn
TCXc84Io4iZkpbn+JfSM7+ZuKJ9bPxCjWbpDg463qBnbU+8zDXdO+e4n+BQMiDxvFAYALg3QCirS
YFIaIhcgx3OhrBXNsr4A8XmkfwGY7Z79Z9xWagDIBV5lIRjkw32vzMtlrutfbhiSIli6M5wMwQsk
kkn60RqGRxPokJe4oJnN8fU1ZpKpVG1lHHy36Z0Ly/grNrNMMJg7GhzaX/AvBM3rdZVont0LNeHE
S9OxTYfp7+qPXOmvPMvWnZolTpHNAdNvoB++ZPpoFns3TL1C9a4XyCHT7Zkv7AANrxnPaH8jPusC
hJ5G7x4722up6DFcotG43//104V6WIqn/4NNyhynW+8ukeyXRpKak4/HHMY/icjoIVqU+JXmPpbW
l4aK92zyp9S27hENnKamjf56jmEWdg+7KsyoSBC/MDjnFtuTyIRE5YSlw4HkMPH+72nHKrq+Mu0E
XM+6nV8yJ17jHzb7B2K81TMOPMNAx9Vzx0tpyZECvYY26FjT7bhfdqiL7QdHDUKKLrN3BkJ71rTu
uNBr5iS1jr3XkmLcDGnT38P5dsE5dvRYaXqpcjJeq+8DiV/t+3O9O7bc3rOLK+QrjiDVMedavB67
j/wwKDfvoC6uUD1migXD1vOJzOoFR3rYb6JFAK6Wo5gYEJ05uJyT8G9B6clZL6b+6sZ0SndZtxdV
e5HAUXqwMgA81LVT27cCWF3pAD2iK5ZXrxTsp2GR4qQoGv91y69Febm5HLgkGBIzdhwBhp898qCK
1WRI3uFLlPkR3RGES5hEmJHp6Yj1J+jgPQZVuHbHGyOze8cHoXf3a1LFbJj+gkhVThrsN7a20TFh
8GgmkxvJ76Wo/4PLxxlUR4FAYcM8J/CTN9GMgW5MrtgTTWM4LVYZR+7i8p4BN6uhG7IHFKWCcZHc
05166ECyYM5DRb4GXVTApdpOzVzahkYwLUl7krBKjtju24er3ROEFW9RmkjYMvNwk9SNH3+klY7e
cvw8LupFqTVWpPwSuLYBN/SVaIe3RdRuHTfL6S4SnBf4DIIjkOAxTfOiYhVDtYmFTtREB5QJbX6e
/IT1oMJBzEexcBv2XPgE/TseWagiCYgD7eGVhSCYm7XUTRqTLn2i60iutBmyCuKa8+cTE0X+OCjI
QiaUewP/lzKkQ7/NXxnpwWCj3SxXQN+s5uoOnqSqVKcw/+Ax1953mflwmSLZxoW5MUT54ur/oZPC
v9YBhzKGmFR283S/K8X1TZkDvmDjKFQt3WvaifSOQ1tpFpQjrc4rxGFfhOC4o6E9RwpX5kYh0guB
5wnkC5FsVbfaTe23p6NbTF9Q/qnZdUW1oi2OdFjuFi93zf8BE7u1VxJGr42Dg8uSqYGg9hzPgSJ9
euFc1ItpBmpwAOG4r8dUu6ojAFNarvmmzUVOd6OwlVrfymDuhqZcuqfqsv3AKmhbdlG30eX2NI4a
6UdeyjI/3ThWJDfGfyxzQOn9NPICDhpYYEaXyNpiW3L9Gk2rrV9cY4/HIcgbFRukMjTB+Erz0HRt
ACNZL4udIoXjQpNktL8/0M7CeMqA/m38NZG6KvDp/ZaX8aAqd0QeMirgJNCcfYYLoOBKsnq4pbkv
8gE62jSzmXnFp9tRaTUIkfC/lTFssFceUCVn84EMrbGAnJ6lPceq2ix13SfJzdk7IohmK8e9NBXM
If2cGY0IAQHYTOI6I3jhmr7fqUC11P0H64SzS23I5p8GAba8CD0TfLQDyuwNjVE2EievVNUWMEHO
gGof1sZetpeal8uYJdaAAk3pn8wN1AdhZEl9uyZKF8qEsx99qiZ1BWTMn9Dl5Xil8aX8G1QF929M
qgftPResbqB0tGxT0B9W0nyax7EU4VPcdZzUVxVLDdIfybK+NwVUbA4AAvXOLGbGcn6d777/fO+W
M67p/4KGPvNd0hD+3tAevVkIaJFMVT6N5Co4Fw1CdDOeUnb0HTdQoe9C8qZWGxXB3osmWd6wCRQT
WSi9K6J2YX+0baChzB+11uMHAgPbgoh/yiS+bEp817lCDoMEjcEOJvzvg0HdkqVPgh/N0uWThhfK
f7oi7iD2eYwsS/s0CXGpq+l4OwVFYrCg4Wy9HKkaiFGu89qN+r0tbsTjUUpahsVwrdAEXGxXLWg0
gikBEp/FriH1Ujw03XZUOiatlzO1+Yvz+aCxn+bSeKCkMGzOLV6ArPBeASCYHqzhl+/9eOKS3Lii
5aBLtmYb1FK8ysGvUnLwcNs3eA1g/uXX2Wez6OayLLyimmbnS6iw8RC7sY+bcSzqwt7KRZlvz5ZN
ESQK6JphtzzWt6nFq9NHlbnKwPoPP2zm+a5FNeEfocDQxTN2CuN39gSerHAvj1sGz/dB+mPS3+B6
O9QRcXkdw9xItIFhX7QDFcOHYts9ExzOBQcNf1cyq9wieEG+OjqADkcsZu+nL7jUa3d3FYeVhenH
q7sQUs9oufOQy2tHKo+Vv3EiL5dEhBvXk42HU/9L1Wwvqp6rRoWeFeav0Ditxoy5bhAvvsnPQ1t1
rixijD/pAugZ1DOSNe2PrlewzxstGirEH+BJZ10XcpbIbPHmiFhBScfXHANb5poxvli1SsKYN5GV
uGoAf7jpY1nn+lIAnkwBwizWXwOFIbYNYl1T1t3m27Jz97Pj69nISNyYl80rSy0x1H41TCJNGrXh
JweJoDqnd59rKp8peq+1zSBBXV8u+Bn/E66LRJR42UXCLg8miX5vVllkclto8k1lGWIWy3IVRhlr
pFvkM9+JEheAr7Dcif2/XVvc2jFmiK3UK8S95fdAUyOyVfHwXSAtZG4XhAsolXcnVCfWC1fo11mn
JIUbg/Buw8zbMOQPOyo45k+lLjYf3KAX2EfpmZ3TdKdGXYC2ZHitNUxkrN3G2v/j6duzKZJE0eTp
YEwNVKDJY0T9DzQwn8xkoZpMZOyPMQPvuthGcpnaEmZ3Rq/xBHzUtnG8idyCTo2KnfLNt9bzf6m7
wcajYmtWdGetyq0KICkC5yGYuQin9P3+YfKBnM8qYl/PjVTIoQmDhF5dWazS63RaOoHmhecyJejh
rkxd4fffBFPCA+ftQkyj78fl+wGmMjZBQLy9jaF8ly0+6Prs5LlqkeFchp0K/jvI5CUrlYbkDAZN
k7M0EYbEw4N92WKwjaRA9zSkViOIzzm9SsBUUON4GcpEakUjl5im9dKjfkkrKU5VoZ6wdBL0wQfr
NEd5J6fHxgIGwzJBXYyo7Bir7dHcmovV3dCjZy2VGmjDF5GzTs848wliagUz7WQkRLM1lVosqfhR
DJB/uxf+iupsz8t9/et/+kyeIP6NscUWXU0KroN4e+ec6B4l/nk4TKwRY3qkYoc0vYRib4FAsPJC
ykm63Regqwm37AsRb9ISz1dAaCenio2OSLpmL/iGaYaOEXUJhfZhdLtSlDQZVAV/3JcufoXMnbSC
/cOMFhxESvPLv+JwaEp/d1kiQBztxbLj3bJJWmrScbzvCho2WcI0T5GF+xCAuIALPz7R6fcogVZD
HZk9Q4btRrEQanVCn2HwoywOpssb0RqB8VNDK+ceeMvEqqQx0Q2Btew2XEO8F4o0kLj+XGxqb1EN
zTV1v5ekxGYf4tFbhckxrCmFJ1zpVfrUzx4WUIhIerRLc4Z1K9t5KXUeKNs9XM9wsFYHP6geYPTs
/c2LtdzIU+SR5bJtRzQ3+II2697S7qJMNMtZujaKzfqDt2pXgHP0ym0pV+wgce4HNkV790FqPINh
L6yLO2yZrPtFHQ7ORUecuYCZ/OUZr7BnWAopnjDBu0cg2kn+YZy0Ra80iaXUMvdrB4TQNhLp6lB/
Xj37/NTbJqUh2o6IOYIqvSLMYKIDyen8rpnyOfshPLfrm5WPi5ECbjf6MUsLBRBPSFBaScLLGdT6
AkOVBN35No36n3vEtUUwLt14YaCFtBDXh3W/EbyWqWUuT7sWr5s6CmAdARFTTFkrtPczPompBp9i
jTzESHP8PwhbqS7TF1H97gFaycFU3lyBze67cBeQr0RNx4JHaE93qjHnD5dx47FMDMqQOdo5Q80t
w0xlDhov+qJWS4/l3k3lxN0ftqpLb8ulQkaS8jGiDzaVi3EzXwYDr4a/PRkRqa9ZTm5ktElFEG+Y
xEuXENp1KA2HBKJCr0Y2cVSGz7sPAOvgWyGXF+ue9s5x4s9uEtOTNUdmZHFiJjVUBdziP+EkW9rV
UppGKhfZ+vGnpZ16JqEGElNGcYnLN5PT2hxU6acTar6UbEK7xBDWSBwOGWOloUqMGG8sHhDC5FJ/
Xol14409O1td1JzaL7AIaMqWAQ9dZ59WiMtEOaI82ymOHp74elT7DCYuiMLXRLttK8IjXCxNnCKZ
SBgTYsYOS17DPURI1Qpi1Im3tbpfbM1iT/uDVPzuEGvBlc6FDhROTSIhuLao3eNcZv7b8mBX/LPk
7fywSxPN5EfX5OjxXJlhG3ZqxCK662XRChvT9vBA/7etwcEnRFgbliP+kp9HOl3xgRkXCLOj+ZYA
cqCNPjY2wEufYs1gD5LdAHftS56+ghxNscR9BAAgxpNjJTnxagviIzKEco34R6ADnKed6QZ741Fm
JVQaOymBOtR2B1pPE00nugrUmbX5cF0nyLe7/Lvs4d+WKbVBzUfG/TlP62Bu6kgg6BhgpgSkoiMz
IDKgG+5MgS9um6CPelFiV/fscFUxxsPqzs41mC+VALOE9blwPOoGGCTiiJJfryhyX+Zj2rCbzekK
xeemQc3oP1oHHsJiLzWU8suyGS2AUbzD8vq8GcwnLxXzlpjO7T/Oal4K8an2HshN7V4a8T+f03CV
+8ou3yGp3iLcfUv2bN4/nK8dt557F2mpohkAmgFEimCosuhqH3cPys2QW1hsS4jz66me/HX6PREl
aFQ5cxVy/z2+6m+mvIXJePLnarNTwjsMX+/9Xl7YRD8elCPFuDR7s9n3X5ta2orLWKOojNUqrKwD
ppqkWURc0F2rsZIbovGO9e7Xp6XZo3+se9cyIbUYDRMAByNcq9QJEpmnCYCqoCNImg3deErXWCyC
vMW4hpyP4cMv2IEaI/JkXJu0jGQA3Gwtod3iUGs/S64vC7cZFtK5Aev8entyxqnrlCquP7DLxPct
oyb4xEUHk3hH90ITO1qToHlaEmo+BkC+Hot1hLWI+iPcShsygvZZwhLuRY4ru/Gma8qsywoEgGWw
HQSVUALGMT2E3CQEEvUljFyJ1qMDbq5dkpuEKuegPZGnr9rJVo1fIrgyjd13OfHkkRk4o3R602Ap
syryLmC0pfXq+KVB/c8oAB4ft0V0+pygJIkdVPofUYDfc0lc+41iXO0yg61uZlc9Zl0NZSBIHw7h
oGB0Npy2APQ/+qJ0BAVcc1u+MBf2D463djmxrBQuMZxdp5EI3MCZQZpNuu+kQa9UoPzrvhR82zYp
/+HTkd0tAjq8FFCup3wDyWiX4wshPHuyTIucGK5kanh8lsvFZY3MkZs1FoKVjbGXpoUUQfDyQFOS
k6sg2GAJpKm9YMewmJXdvS1GRuuINM3vYEWP7zX4KA1wkc5rQBJlg0dUdoTQjnjsUMGt8M2wFQcm
e7fSZkEAQEZFOytIosNfcQWeoSKOG+2WKmoCVQmi9UXRFdxpwtK93RhoPOC5tLpHVNG3y8yc4mfj
kwLsuLEgpZsReGkr7RgNAwBAOb7ErBOPjvRR+74nscQtFAkyytHbc+w7enOIMen9UhTDINWNtvOA
RdFRPanyU98gHQQoctVNdycGMI6e94UQ8aC2XnX7hKnJ/d59bX//FL7D+FH8oUjBjZuJs9PdTzrX
eye08yDExqXis6pm+TDjtaKV6Yy/hWTjTWsZ4tdl+eq7MgqWIoAVVKXRz81Vb/IEjoVeZm49loBG
Jk6HtpMPDuOKBc9InBkjlojjj0F4DtyHSAqjS/aF9xkIeMTBuObUi3V1wNvD1/8ZfSXooZ1xC2ls
t2qQf4ys90V5GOzmsibXJjv1Gw/59VQHmkMNfKt2ZVNEZHAoc/CNyNih1qunqhlelZcZEC7zjDJG
R1SDcRNCL718DkqYRqZRLCy7Clav7NJBM7wAqQN9yvQkLN9pqc69976kKWBLfuyubB6aeCHIc2oe
pzd1a9MQ/sRNZrsIGmbtCL2oGsTJiaXGaw9ql6Ph6eZO7Oj59LrDEmp0ITOUby4f1WdKYZQVmcrK
b8dXVW62/UNo+NkwQ1lVPwixz0s44tCOFX5e5ETTtsb8cVUSnmzHpT0m1Vg4thyyfatekbszAPqN
7lUM4onByILXiNz3pVVh69FqQhZ6ozwcfc4GnSUcuKKF/7+0bP6CygS/l+3xpMMhkoL27VBzbm4/
9SLlCoA743evnRSXRZgaQvJf6/b0EuR8/iUVeYEC+j2vzdmDl/aWRWhOUMkU2/vZg2iaHPJV+W8j
ZzVJDyzRPLYj8rMcs4HFdEVHGAogXic/DGR0oHVEdoOG5X/Dm0y7HAc3aypTGbodtiv5Y6Yuwcjv
Y4/r38L20gTQ+y6asdLv4NhpRL7b9B5xX89d/bDu+yE20dmoL9jhG90jBHB9YTX2VXd78slGipmo
5AP3CGQFoJWsdeG9dzmksZ6mrUkIHFIXE6wtvSbuJo3IDf282PU1wF7NelZobHB8scBa45vGQll0
9JoQrZCCfiK/7PTvnIIRmyWnjkWDeNJ6hVUKZAs2PN1RXiL/9PKECTl3Wn2jYOWPY/rW4AL51Gmj
A6CjabNgb6c4566U9zRMWAXKYYDDQGd1w6PpY7qOg/M9PeYxOEH1HrelaN4GazQtVyP9+qze0ufG
OQhQQ42fZjAZz83FLZHAWHSHM16qrF9txepIgjGJOUN+rBvp/bQKnkE00zC+c29mnOR1sMSy38Qk
zMog/fNr4lZ5t80bkJKe2gTcT91QRR6Wfrdxg9hRYHEXokkq6GnjmXcZ4YKfoC1JRklVZsS5yAS5
q59F1AiO7ScLM1NqrM+xJlIWGqmk1SbFLODY3ZfaPYvnQSzVRZde2i3orARtXr1Miy/DzGa16SKV
GqkRebyahmMFdl76yAwA4VpG0AIA5fZ1cnloa3E+V/xCEdRvyDYFpGnYveddsU7XxDBToj9/gMUm
+wmCLr3ai3M59yUPAslzaqB/cV6ac0xegRlJHpyybf5XtaTczbkJf2YBBJyC1Pw4pcJvuD+BDWhm
/PINwaki5de9dt7XOM5+ZGVlToaRZq5Hlh8dkQMoIvzkgqjIdwdDylbJIZIe4nq4cRFGRTQoOLfB
+uyPqLdvd6W7x01Xlle1du71PWAbsXRS7RJIcBx67fWlFzsNbC7iKVOD1hE277/BNx0GDvWu+Rgd
NLvEDg4Vp51XuaYpL6Fax4241t56/IC3I2XmiXBVPeHaqXMxyWOGFOrJrOZjFU+lm58r514V+nYO
B8/Tlf9JUglyuhcTr6SEQymKAc0dhsV4p5dtvagMl+92aBQMhLj3wqSjmZ/Fu98wrc1dBMgQLc8U
jRgDUT97RmRIKkbmsrq5FKI7xKrsiWbhN0m1V0vX55A+nHVOFUBgMloxZmqBxGnnS9wTWDzabMZy
8e/73Q80OD5BM7EDU9wF9ubnPWofuR3jozs9C3Wl+ZXutjyfR9zPacn3Pn4OWGPauYeMD9Ul+HKS
lzPQVeYr4zn5VdxZn6FSYQ85B3bmW7G4qs5kfAxjQQVX3DcUJ9cV2uqqLVaH/5cgdTzOdunNv4dG
qtYzWviIDdA1sNaXQtw7oaWe14cXYx9Jt2aZBnImo75BRv3IukA5BymbuR+HWj1vfNiwXD/AJyQZ
7JIpditmrDBHt6zm6O3M7AMBLYmCNsYN+rea7YJCTPvmvhT+OB8f+fZYLzQlZKfgLi4cT/nBUK51
UtqDcmOk2yqUuNVqUdPR1N3C8GUTR78bCdALABjQlGxI374mGr+NcuMM5Nwu/pkOMpd1C/lnb2Mo
bCeWfBzvDvUtE4QjjgScghWktfYZtP02cz55juEpfF+44fpv7q24xTW2GcRwBOf9tUnXkBmsExTX
Ja2y4fKWL/Cm7iOYGq8fbU2EZISjvYaFy5yIO5apnQer8D9Nip9mbbc+tlxy5nXeRZyhtm+cYQOp
0ulEvyCQb+9cE9qQnp7ZdbjQew0kPJZMlx/trw77gGjPiaLEBfc+HQceO9Ib7jmtaofNDgcYD9NI
Xra5VtUH7bcHO2OkI6ngSV0lduG29c3qI8erfdwOLRuFzWk7uQ2VYRMZIwzBxrAiuqExvXcQD+Uk
u7cQUQvqR5jhOrJRsmznoQ5WMBL2J0PWuky+49P3D1huseKzbtq21yL/Uk+CQHdJLNF67APF9OwF
ADw0Uv1N2ubObNpdb3kZmLcwW/VDJ2ZBbSjBLrr7uxew3TT+Ar760BVCIlKs+d1updEniZMa3nz/
HTHFaNC45bAZiAfKxJPvYyO0AleS+WK5UJ0cql/k+MsDvEqY/tWpi8IGEk/A/zmBsrql1uGCitEI
6TFAW7qKN2JWndbc2oSKgOKH43/2UPqM2imUjsJ6skr2/L6ITNpLJBb1jhpjlgelAM6t2CO730GK
mfsLM5cZrRzlOVVovqreBsFApbJHTzfHVqWL7id9qOif4Reh6GAnSSJBp3rHY7Kovh4fn2kcPuuN
L3LcrHM+P2Pg/bDwl8M0ZsS68Ai2otkio4h/HsKvg77G3aUT6xcMHtomTkNUCE8Ps/QDm3wENLgn
+KZ7QOIGyT8eHDfbGWO0vZyvSi5U1zHexO5gy1Fn9SjUQzSbSFwL0I0IilvhusZ+pEj6cU6+ZYXY
9Bq4r1x18dH+aKrIspsyay9pM4jRuozG42cLsxMUru/eCjB5laPEqC+2J75yRi/j9YLiCvWtjOhj
4kAFfg5xw53Iyaanj6OH10BKHAt9rV/wUlV8m+Tk0GrUNdtRng0W+t+BIc0LKgtYo6GdYDBf8Fze
c2bIivw9e+uLzwLWuiRN1Wunz2VjcnOhxaktNyV/99beecntypbd7ULKtVnNNQrNWWRvPv1OMYFV
DbvP1MOiCi7Y1G2ixVSTDFejHeo2z9eBCEsDpfdiQ2gTGHnLH4nz8TqJ2BBZTpwtYrEjmpMR4SXT
FYjOdOj0YB7dJMxXXIyVnv7xlnadmJIbGrTtDQP8eI9ODkeYuPcfVB7viN+eRlq3Isj7rWndnRh2
pbkbvlRFzl7rKHBRatP1fBLqWZBVJsU8QGxveSOlDTOnykBpJz77Ci9N+RW6uyycfeTsnTKVIzFM
wtLDiJoMFL/novkUn+iWtUVB1btE+MiZ+r7vQ9nb6jZEviIpzg1LpKL26TDvKYjehBPwLXERxN+E
a5RPmOIiHFpxpTxlcP0CfQ8KPZDp34AGpUoVi++JX3YjACq0HhLhGMj9lIku79We1rRLMGLJCSmw
hZp3I3+eco7Kz5ZyiwTXDBNJsuk7ILK1o2CjNwCsJKlf0ldfBhWEN+SjOUKHtMuvjGajB78JIz6I
8Q0gG3ZVb3Y8gV4Y/S7SeHGrdUd4LCXRZX5U/vxemrxF7+yQjUFWKjrJAOO6cgpuhycuG8U1p5kT
jblEKi3Y0ne7wDuC9wEECjJBujFXj0i1pTUHINnQu9MnDlXHD/7dVCOvliPa50+6NJO/z/q6+Xr5
vL1cYut4/yAHVQ27+yrbpKcZjHUFEljRJArjPoFY7vNv2i8pM4uOuub5EnkkzQTqT3Dp23wwCevb
csT2rO2ggQK37NgnD5goalbLlF3NSAdz61neI39aRIB7oU14RT5mVeO9aozWZfVXT+/9aHEMPUeY
2PIn46afJ5hIXmjtAqjiL+XiiBaxkOoJpVu9m7rqAtZi8gu4PmbFeKAgkSwdjHS9QtYCm+FKHprF
4OWaMhtsQ5GXZ8O5tupOvFzar5t9ALcdI2PyCnyvkUrbm6jk49YfQExaTSNWWSqioXD3DbR8l3Ds
eN7F4yK1PaWKHwjEWNV3WQhdy/mPf+kNUsStTp8caMGI+mHH43s63JHaLjCQ/YOKElcBjK4P6hhb
2BWuPxmyfcK7M7Xqp34IxWhF/Kxg9JkjLIoA1WYF31CjrKhrHTvJHdX7pMNlPZxKM1Ok/urupSYe
lfXULRiNZamK50x+2xOo99pHtKZAzIJ/74VDeQhWWiIbYCyncEhZatpL1G34FieSRvDpdJMyOoNk
ubqiBe52cHfGTMsl62jFku3197oBJXG0TxYE75zTHuX/3RW3M2i+t1JapkZWR5wt2GMflLJlQTkF
QM6Y9wOv4UxZBaojcgLK/geb9H3eKloND55W/RM73/cXNXU99UMVMsr9I/ANp81NqL9R/YO0gMZ9
q9mTEZyPB1FZFllPqdRkons89X6V7NlmVz3ihdPhDsvzI9uLDsC1v0sH+NkkyRvqjb0C0iYbrqN3
rnLGorFpe5gaVmvJTiRg0qs9PdjdI6hdBbhXqG+69ZI4O8wAg7AwlzD/aOjLlcQ4j4h5DwRxdvPE
40HRJ/1vsUubVmuZb74BlITxNB1rkkiQh15ZI2OeeafzdypKnru9iA/fDc7VZOFpvD5PwB8xGW+N
be5kDzVDIgDRFH7xG4xRwGEfHxEKtZsEVUikhJv1J92F582aO38btXYJRTBpDg2HafZ4shCto7ti
tF/+mdF5NBOiktBpiwcoX3WDzO+zb5M4Ktms1LwUL1Wms8pLr2TO345I/XUGgociTkq6rEewUMpd
IDO4stj1rFeOfitfomwEZqu/dS7eRMXgR1eyhhf2uJypgUd0gZdaW5EJD9oDZWa68GYOIELVhqqH
rlKodTfwYXA45OyQ2W8jUyPm8OvAfUv4jfpRnGBvvxlcV7YRLKdoGx3oyJdLhosWCDUmF2Pu11Ow
yxfT6Ri1ZMgz01jNZid4drw21yI8s1oUBAvreX1YOKMokDHN9bu15QfNEK6KxGq1CNqzDQOeYaVm
cxNesSkuuk48eqOSxkxxBIbO75G5BCKAUFGMr2VKZ0M6DmLhKHTjItYe05qP1WWtth2G2PH1AcUh
Q3c+OBlwwR7KYcBTyze1Og8JY+1uYscBIAljRlDTxsYGa5e8b6XpDYiDdpY8LM1+k9OeS1jhKMTV
FXRIaW4cVC+K4KGZTKrHI8C7a/LHayanZ+pO/Cz6GpyJS8U/eBsmRK9aMQ2CLaaGiX5Ikc4yYKvt
FSDO3IYT7gJzE3g9VYag3uR1ODITL5PXF0TWBIsS/0/MYiO9Dk31SwrK9wTvNZhs2bLJgfiidJxx
TQ8/mlt9pA7uATG6773RntBwWknBz8CLnsY8DnuuAiNk2l6/zmZcRkRcY++LoELgIqJONd6Mw9Cb
AZb6lqbbcXuRe+A0Nz28bXUDzwkpf+FAxe/qvoVGlTImuoqoKC1oW40dWb4LFK+El6dIsdMlbAe2
19j1ILlASY3Qjx92PbZd0o7DDm1UXInFwx6s7KTDYxcJsyn6jWq1Z4St1ze4avWpUN/I2t2IsBvs
0b3W6O/9GtNGMg8fjULKB17oBbBugkBOjLFQuZsQKUxqRQZZK6EYe5kW4a+WkIn0h1dViTbRn9rs
GU5hOzE3ZaNZjr4D4xGi41Atlex5tlh3nBthTnssbOH7ZFA50k2US9K7eeeMmNH1DI3pt81CnbA9
avjbyN1urs1vUfgBgClM0hEaC747E522WfpqWLZZLNj+mbk/TAClG4Re88gTtb/Hr+BxG9KBd6iZ
KUTgm2PqJ/uiti8r7Q1HRWB2LDRg15zo+on5ikRhum3Gk/bpILb1A7w1XGuSKgq2TovGTiM2zyCx
Iijp3Xu3+Ol1FOMfks9vlGUdBsPf80BaYeiJ5/frzT/ZtK14DKct7tNXVybYzji7bmE11UbfY69P
nOy27QPGjhbzwVtEmmTa+6iajESKIUTW8CwA/7262qtvfQ6LmG3J5M0XqDEEkVWU4PMmo1sPD59/
I5jejtiPs778BscuMRrRmVK0vIO+/A9fh82VWBFEFF9sEJvkAwvdw/aegfDDfpCPDOgXlr9FbGLq
fsB6kg8+69kzUmQLUBWfc3KkgJvDoQjhOJU1kO8e1HIl4xOnEtXopyoJUWcqEydQ6iwVMZlzIM10
MQZxp+5gNOJ10Xyxul0x7f6AS2CyiS8sbEkGfLpnb3aYSD6UD6NeUNSZgIFulzKXWVM4Gj8e/G/5
OpSTVKctdGF2XxiAxlY+21ja0S8TlAZico4xYJgE6F3eAtyps/24luW9sCI4+xbosF8CtIyRIzvm
qyADr2T9lnhfc9cAJqB8xLGzRILFtP4me/OgGvhzhl84hGQR9VX+OLUha3qB9NCmVCXDHuxoEsVt
/Dh7+UWMP+53JozheMvGQ2owUjL2ZDFdyF343ODzU05U7pn1gvNd9FWnSEtulZWBa+EMk463rYq7
Dlgfc72aLPRMxeZGyyLrpVF2UwSMspoLdE2/9W11luDsY6ou/fP0qq5yO+IyJuUlPtz0iDBS8mSh
73cQKrvG2l8OQjsGfZ5nD+JvU8//yp9Agk9DF8Kxbh0VJqMpSE7jktMEbSjq8aKPBBTy0wIhYriU
AG3AlbF+KhcIbjV8+LYqKFzvamLHKkuwjH7bsbFkh9QmoNtfQ/WhdSfNA1+S1IXJWxSXJZtQ9E04
aVwRPiufpVikzYNhs07YGsli2I1UufoAaHzlWJ7B4871oxp9LIqP+S3I+e1ufC8aqsFoPHqMGARh
eYKH9qiuqAQf3AjSlPUqSFCD6FDvofAbJiiWneK0XapETvY1E2GG+HRbzSOgijfwD1r0e1KgCodV
TPC2AheESV9PHCZ1Wc46ze16wr+3nRZxUHyf+zxW8OUlGZHaiVPD6mqSoSqzCf+PEoTM29Q8pOzo
jZsU4OuJZGRAKTAXPiN1FW4mDvOWEmvA3XLsouFBD3gMDzy5QCPsz5uPWaNgVxui+qeTwBgQh61j
HfOJRlcxRZqFA92zVAMShsgAc4Y+GgD94wMiCUyDRb0NsIZqlZjy728eWfyB+FwT2d240htw+BkT
LJZx+gZZH4BXMOLR926YuzyWTOQkBKhwUfbri0bMhT14HHuDU1vMwTla27yQUxRl0DvrR5S/fFGd
ex1o5d2ndXdRxZZaqAdix46MMCzjFfNKTXshLWE7FsqDqyatZvag0XQ+egFmsmRWSiIZ4nLSdf2m
AdryQqe46UAGTQwTG3vlaT0eKSzwzwkfjIyC6JjsDCQDqHwSA6ZSnycQJz5bwAtld8pneu8as3N0
CR1cGbX+F3AXKKxVDmGO5066q4Fp78+VTVmWSdhDcZpumbeIPI3CgqGn+e/r8gETb8ySwlyLDgBs
8EWEzTvSmNAD10iagqR21heXWnmf5Qvru7oX5UR7i6o41/UzgP/7VmDN8oHnd5G8x4LrkSvVvdd0
TgjZoUvdUjz6w15NnwSO9Unu6WglP2MBo0Ws7Iom20eUXc9WFkRRZdioMaYu7B8asjtpvDaQ8b0t
s+qx7vJ25GQPWP6l0+1BYn4MwGQE86ZlvXpTojcIaKlaY3YGl6QHtoBR8AGTyKaGVXwQSfrunZxv
qiT/zCPHvNdBkU5xX4llWdrni+yb4vLOZtVT81SrsWUiRGYN0GIKadmuh97oii88363surmgZEkB
pk1j6JyCGR20V2aksrhCzbqbami3tzmyTbGCtUZp38moO0T9Q2AHkgUbDJvndJXJpRr5lRaf898S
Lx1LFR0m5sQarrzXiJS6Xwj1zWptX/66hoXaABsxx1LxaipjTpCgfX4c2RL/17M7hjAhLcE5aJFZ
wTfiv8Gd82l1/oHcMhsfTmpGVfBGDtEJFWmq3pew5nPnvm9bcesO33e/iDoS2jNZAR77fybkpm8Q
LjStu4kF6dJ/ez8QPa1gs64whNgU2YMqR2fpc3qGabrLiMHkNn0x5u51fNcHdBNCP5rL/H6m75da
6VxmN50IyohC8JpiFM8kp2Do3EvvDEJGXXSadIrQCFUeUuq/Z0QTEa5A/2weWbV2QQdWH9ty7y3L
zt71BefNWoUtitv/ZLbm3NF30jmYF3tJ+ulSI3QL+sW0dYX66gNMcDvqM4rXCrQ6CSKefU7rx+su
/ANYh4ROGjVhCCd/z7yZBcee+mvMFgdsuyeeX3c/3DWPj4bFLdDULq6O3bm3dNh4Q13KrvPEq4m8
gHN4PB9hxYD3n9iksoJhN9FDOXHnFPXrrpi3VTTJzXuk13P5GsOZvM4hb+cQ/HQkWAuqoe5hV4wb
mAyH9KVPTkAbmZvZTB6bRNo7DVQWxWvRFzGo5G6Lo3KGX9FpHqqo14+IxS0zKbG5l2bJGXJTgTpy
y76CZTYm1ZKN37VFWoLmu8uRfnuDxUp2VER5AlOw95lYH6/eihbY4tvUq7qdz7HPQiOIuCCLh8CQ
kI2ZufMW/C3JpoGibfbNIhP2pIAAnFbzq2nCm6ibeqU8BjDYfRnnejB2S4dQfXxMXk2Ke/7w6Kfw
kv+DV5sSfNgmhjRg6iEIsv52bSG6VNgrk57up6F6om1ZoTHNikZqrsUdpq53Deu5oAJOhqFIYuSo
ZhQ80UESMolGtnhEVECDAmvP5WGpaQLM7RiRjjsLQ75cUcG3/efxLs9lCk1LEd7TSXZmFx7KxOuB
wJk2QHnFIoiCa+Npz22b6O3/YLMkU85M5aewxZNGj5JD8sm+PMeY9JSq+NBPiK77t+UHTInVZLvy
U2RTdzdPeyC2EyZKUPrHTCG0g8iw58Gp/ko3OEF3zzElJJYTvSWxFLPxuRX+FIM+nzKFFDy3+/CN
m4DKfoa5z3uAQNgXtiMgLrvceTsyoyKkV3CG77CYCfwFwSqIWrF0dLpL6QQ9LbReu/1ssoN3H0jX
FAEOw0sKiBX809krSil41kSCLa9ylx+R98cb5oaBeubu7a4pbndMKc9kiF3mXwxOyerBNUrubWnx
acXx8BX0z9wORpCl8h9TdkqEzUWiOVbtlYy7XBqBIlRPXfZdGChjuw6IKbINVY3TvP+Ij+VIkshl
KUqyWJbcFNMwBSUKD3cRbgxUy7WNWK08cMv4ZUsL4UKi3MoVo7cQxRbwDihUWLTV8uaMGfb5dETq
0xj4UP9lPNjK/GmsOUMwlGpz5qBpK2l6Cw3gH2lLpX0H4VcKswrFWLSlOXIVU2qLx7mVwjl5Dee7
07rtbJmqzRCGcAA1sUOkr51XdR+6Mivu/EX/WQYXjturrf4HzB5SvvD11BdDhDhNDk5QTTfnmL/K
izM9rEpcnsO+EfmgWZbhCLUeUPcauviWqHT9MQJmF5NwXn7++SB0vtrg/RdP6UbYynUz9RcrcoHg
gIq8//dw+Ry8VoI1r40hMUajNO93Fiau+Tfh+j6+Ec/V3bVL9BL8jcY5J/LqfuPSAHijHpHq8Nri
1aaLoHBQ+ZaSMoYmWIcOm85OT/minSNwms8znByPY21HZqFlJFhzc9jwYAFTE9k51rbwnj8Zykt7
4gr6e3GFJj22dDr9MiyXuawD9HtPcy/EDg0J+jD+bo6v/5MSuXcwQjkVCNacZZrxufRkCOd61vC3
ZtSJszW3pZYPJ5NVAE5v0I/gLiBuIige9RtQ5LqbenKnAJQkz1NPYhUtPQfVhadMH9qvBlg40YE9
wxGiUSsFB1IJfdkRE7HGTYtmxlvdfd2iUWn7C/Xsr/0itm+oK83k4+NGfP3qFTjTY+nnBOjOgfbT
vYpKGNUUVkzlHq5UdSO0kDJ6zt0uvm0RMuEZO4OA6abSgZNZ3txN45aNK0h9jhhojsMPIjO06IG3
Ymaed9Tt3LfTXR3GaITKolpoOxZZznGs1Z67TeBe8MQQFtnoDtHQxFUFTR+05iPNbpYYIkBYOdq2
7EzZHhiTc3orouAwuA54934EyBt0sMRgNJHngjdrCRn/RS3ug9/XS5zJEph0hD5D6FGrD0N5zDN9
CLpo4EdP0AaossVMd3yB1ycilpSP/ealE2p7USw7I/i//6cGHCTRID77AJ8PgbAJPYZvv+HQ9vhb
eGNxCWBut0mJu+kHz7m/orhW5ysDfRMOuRIKX5AF/faV8mat8MrA64Qo9hvP2S+2QKMMH/vIBsV9
wW0qWlff+OrdUh9KPdN8qIrDt6L5f1txbWnZFG9+lgwCLF8QNxMSNQma1c6z8Q2BDZp+32p9UEN3
oiKkOpqJzT8WEQN+sJBriUVJkgjD8sEwTcEFgG4SIdegWPhncZQS2w91Kk2Koh5FZBs4V7MAnSc4
s6bZHk3Eo8804OBr1bKnIK1swtRZ4GTOzmBpiTET7ILagIryfZhE+OAyWS2nlaBdjhTGx1/3ZsvQ
e+M5L2iGqgz8Tb00jcNsFuZD9bg4JLzFzv6elY/B0yspTQClxc58mpPoQ6EIluC8OeTgSUVF3LxK
kp1IM00llJlHKveRplX28BhXIy5Ac7AwF0+Mv0994+AhqFDn+H9H/VIppEfouuG4Tg2Vgc0GxLgw
TEQYO0og0HmaiQC86d1WBW8e+7d5Lf2PorcY+9x78FeYZYmcOuic9uDdedg5Frf03vsVVZsLb+Ry
FE3MFkWgdaFbnsoQWSc1gNjURt5CzFFpPzxRLzwOjWNplsSZXX7oqHT4b6b8cBXFaU/BKItBPPEg
jLSA4gx8M6rWVzkQS8q8+dmwLy8ZUCUp7d3FSEBAH3jMrMQH/vGEz4S3TSeQZUh22VLzYTbiQkOf
i6SAceB/RzC9xUx0XRP1qMYh/5dzwoOji2ibv761Mc8U8WMSqtLYDD3WLC3qbOwPymTCSfy5pWAB
SK0MrUrDouP8orFHPuQXLYlaocInh6RXigXRQ9IBC3xbiGWE7W9AtItL9SGhsPPc7PU7Whe0gWuS
fwBJP13reuu0EBZwbfxThna2db8VzAndljOAOSuBHx4nyBc3sJXJzaEDg/lQKRo2nanAH/QF7Zcp
n3AOKj3+bmNxak86Jw9EyKTAFJ5Lpt0fzrd8cI+Fikl/KB111oZSxAVSHFZfa0J6een4WoO59W7e
OKrEUgc2IjeWq3I/WZugDcjS5Qt4XTX0qIAjMC+dhixmu1qdJc/C722Zma0gtiKaVubcDa2RWufz
UtM2B6dbKE/B/LRqfXggHIb9cgGX6+fHqmGUbiN9+Jc0jCVa6UcoaEVVuRHJH6QLf13RPHZQ7MkJ
QZ6Z+SQLuWP0JpfWF2nTvcjd0qgYTJyXpFrqsU/uYJv7EI+4pRKhrm7vI0iJQFkiPCKgechwvZ3M
fYUj/RXaSIgpHYF17BVRAetdvPdC24UGUKNZRek5uIXvZfk9YLPYOsI/nlu1iL+ujfyjKDcmCFYx
wbufc+L0NIbQMXazzcrK0bkMF3G4ZBsHelZC+l+MtanZqZMUZYsojuQtKstM+QuGz/Ex+4OFDeqI
iegAZLsRCjbd7a0Y0xriIeHKqoLgfjAWLnzQ8Ctg/cb1LtmOP/6on0nsYBpj2ckDOkxGHwXFtI8d
WSK8stNTYt8zbqwutcrUjGnLtfH2IAYz2zVBUROwlhfDOY4HLs6jH0RIpSAG0TBw5A6gH1J65lUu
JhCVl8ECPKetNpJCudwTp43Bm6sEMRHazC7XXc3iv/Y61H9MBhkodktrWqBr9sNIkPqA979W75f0
09Xem0SqkY7DscVssse5+M2EqaKDAoTRpBKdEpj/7FRifFazICtv3vZ/Aatdp8kLeQDb7Vr5gYWI
baXaVgmCQCWX/dtvay4G2wfS4QlqtPKwTKNoWtlOSmXOpiD0JNPnIY418dnWM5e49cI7E/g7NQbo
IE2bKBkG++wLS5S2qLFPE+RQUbxK5NO/VztP1q9uwbd9D0Jqj35O11GFefCHX22Md22NUo5S5pjA
H6ZVCS+B3zp8qbFcGR8HecCLh2GpdvALPtGDXNGdz0hsMn5mE3hdlpK2VgPVFxCbdO8W8iD26BCa
B0toOxxuyMPv+skbk2W4bqtKG507G5dEyVCXRzxKq+Y0vSznOsm0XwpUuoQ/J8SYmeBYMv/MD3Se
ldzrKtsfC/Yp34SNOe/V/YEw6fuPHnQT5KwlJ/GiAV4unA/dIWN9o+RWztAFioJKjN4SJYnJeNp/
6WSkAF/Iqeth0NbugjFBdY3HfV2LBvc6KOOhNGPmi18DoGNOuH3i/i5GkLvzv+Q2NdIu54nK4Ds7
5hbRppwX5meWymswShZJrIEd0TS8gn6zwZc0kVdnOro5Heo9SsgcwOvSLZljLaMm2S8iktoM58oG
DRjL/6Utz4c6KCQye7QQym0dlyVCtOjWNmMFxbrzMJF8DC1FjLz1QpjzH3Wa7KlVCf591v5wGdYn
BGs5GjGZp42ogZTUt7Nrsi/TwCt1QxGlATL3AacQkyWVsMKidzFU+nTdZeL8P3LTW8JAz3YGRCJe
6dAsj3vT8/BINrqyEFj6NxsP35QLRZ+og/FDCUzFVYndfEzlZTGJyfrqAWaVtRDP7mHO6tSSmILl
nrNTTrbUHWuXn4ZmJVedgOYekGq10ZSX4Pwzd3SViA+srnSZqpnWciM7xjePse5E1C06Um5Sf/gL
zN5Vsgw6vrFxP/RG81q8aJSTqhMpoQ/NcL+AIGYkj7lhqlFk5U+SeLOB0HErJ2fiYImlzbX2qT6E
6DPupV6/wdrcvf7uDsCkru3iUOTzHeTLHAHBzJB3APJ9s4oQhCxDqKbYIn5BP1rZIDbgjHz/3EZP
YBFm5KtsVf2kplsUMaRgNIR/0V4NmL9hULh+suNn1upI1B7KrYcRgULjdrYdq94/FnBYMX6e94+S
epFwNw2SIPH4WNFWVXaB/bp4kQt6OSWafXc/kfO8rJWAL1As+8+pu9CsCeZa48ih2XnJQmg7Yl0X
42jXR02kdcntk+2urAm28Bm1oNf8FOkZ+FpxG4Ck/HBR0IAwIn6YGD26ot5l6jo3Y00SLl4dOqa7
ffm7vkFkZPRgChSN5OVVhA/UsegJChbqRavvPKdAUa0hjtHIuxuGi8rV2C3Yf7P8Vt2VhayfB0Dt
HOEUCNXampe7maxyOxLRUwhwycFVmqBysCIHNbvpxH2uMveHahm8DzT4pbhQvih0HFKRIanh75Bd
otvmlQOA2D84hKdeeVy5z1tw/6rtobcxFPGvs2DelWQS3LzJNsfThkfbMAPqJhb5DytnkCZl8a3H
IziNoZMz51oX2jbGkbByuftG1q3O9uEQkV5GTpEeAIt+iEF9cB+cn5KultBEMs8YKvUiiiUuJ1WI
D86zdFf/TXP7wjZV7jnm6VFAcg1eKJuGZvu4EZtFo/Pl14hHvfJIYV8fjXU5KeOb2M7ZWN+Gu5iJ
fdTNp+yPW0Y3vNTbogLDDTf5GZNTbJdwav3UHM8dKSCJCS31FWXOcCGrKa615+Hs35q6GuRE1JdD
erYKN9j+W68yVJ9RhxLQeAxc3fRVg10eayVRTD5GD4+MCb7z4lyCSwX7B7gH+WCPTaGb9n5/3C4h
4o8PGX/4jd3M6CUYLLekORCiJ1ShLS/Py1NuwTY5+LRJu+da8+ev7vuZk2/6BnfbLciwsoUBO1H5
AKIEk3jj2JqyqD0jvTpqfJRJP3gbdOw2NZA99T7YCpER7hXzmsePagixsNv+FjebPD48VoYuQe3i
8dlV/T/mo0M+RUTOnfzz5QldCMppoXAV7SI7yQ297SjqtBRACziJZW0aYbpXmWSVxqbSf9CVGODZ
A+Ct1uKgiN/bD0AKxQ/2PQ7GlHYqkCuMQiO84zNh6hrGUSYAiw7lz98Tm/Sc2sFjnm/K8j3zYOJE
8N2V00Fk7KH8EIl2AWXif7NIWreD0URS9IHax8iJSC6cc2nB09Hn5jHYSFHoS4vsRpBd1pHoWv9k
nZhOJ4jOVMMD7/BA9GKyshrcEQZUfzJafMoeaSQtJj5X3ffE4Tm2ayRld6/UpaWc7yRLoTXrm1aF
vxIczt6Cf+ODFsm2qHGRB8Ipq0+8XPTYXeuP//Rn/Dg3nfyjIKj44ygixzwnO5Cz7JtEqAnEAQ96
9eYL/hzbhuJxWKZu+7PGnLeFzMEuZ9+s5OPZ0/76wilcmsKoUl4igU8jaSDeV6vMvE2Rynnw70Cg
w3NJiOJsxIJWAIK0Tbfu5pLx0RCVahUN+ZJ1o5yfh+h+ktwGHQrY4jEHgTPfxpvaO9YkHoO1m6fR
0KeplJ7UxZukY4RDpVcT5J0vYaQwmi9fkPAGJ5ahmGBHq8wLySslEH+lNIwLEoK68/kNJoo0kEGn
uV3PuYN7F0BuneV2ScRHoRAEAtV3PxDJ/jnvK54G1a6mc5EuvWTEfVbtaVjd2B68DH/PuyBT3s/w
q7j1t9gLhDV8kd543U6b5NJ4KQWWuv4Udh9XPk3F8yc6QMvheUKL4KnxxVbH7Ai4sbkwD0S+frfa
/WzIxFJxd3RF8g9GyIDHLGaUsE4okCX0/0Ye8DR2L42U0GhHtPI254QLlJJSiHo3GVL77MnBHNDW
UE8p3VFWP6WHA5Vta/PbrOoHcMuZUpcSN/oMOoqnb+jSXQ4Iz0usrEf3vCRi6IrFFmR2UUm1oyg0
nRK6p5zmoDDgrwKLl5TMsL2LQfS/HgpXysxyo9jC2MRMTM71vlXibslIw8HrYGYy0AJvL1Q0z0TE
Fc6azD8gdWzfmZmgBUP4rCskNCLwLYdr6Qh5r7v/CabPFkdk1U9fMZ+lgdq71QR2fWnCqEKH2322
3x/sacZ3A0L/FDp3ccQ82+1CZ8OkVDrImOsvKot3hxcNbwnjgyXHa7cUi/oZZlNMMxToi4Bg9hYj
a1ILhULLjkCo+j49XT7yPnI1O5Ng54NtZBitI+FunN0EZz3Sion2Mdl9z4Ql+Az0C9cHN71RkbBt
52YzIzsvXMunrB8tf4QFA3KACA08fUVEkm+3IqGdZXi9YxchIhPOPplSGAfMGmKJeORgE8u2cKPE
gbXJA4FzwHVyYcg/rxltvwxUNpcKp9oUf3KfxLPt0xhCDGUFR1DGkOTOIsd5+lhHZGusZBu6hIMs
KPHA0nBhlopuWBIByXxho61WFm5mIyk+VgbqFt7ZmIv/qNPD4a7ay0hBEWXhuCHold4Dc/MDzIuk
lQNKxRWImh0FMrr4cHroU9m5U4tRJP8b30dVzWYm4ydhgtfQCRY8QhNXSbPUbECbGyphkUSA9dV4
N66JK4ytlVdjNHagjpawl59R1FTj0lKwax0iO2pKhXZvZir0sbCCyBhWlT+lJfrndWQUMArBdpTT
stwZRIFFUZo+8ZM6Bd6CGTw+5rBt7lBKVqqNJkTeiagl4jVvT8s8wEXvh5SbYeKQjSqy+e4PUvi2
6U24iUVsXMn2EgGlk+9oe5hYk0WyhZr3CL5fTSiEfi4EZEHXiaKGZnCjY7/LWQz11GWdCiG9qWD9
GDI9H+vLsvCYaqkAopi8qJFnOMWbLpF1GaNIqz9XvDpa1pAUI05L3/O6in6+/8K6Nbp/Tfhd7wHs
gO2rLICM7pfQW6JRQrLXRP6x7H8xByNJldPMjZMGohtec7WZBYDQtbeOzv5ExlB8GSZYsZX2zxfn
b1SmBX6tz6NnpiYzFGLEe2rUY322wabbff64tvRy3Iw8g/M64p4kCAM/VzJnjE4n0yfWWRPBmbkU
VK6ldCubXGo9eCrRP6VIPvuzpNV3RZ9be2qNm46hJHxNIoH7pv1qrBTRU6ehD17+RucCUzrLJo7P
7luSL9OySTyNYWbMqzRF9XrxIB+5W3px+Wk3AgTRNMblciuhUTGpYxN1tQVmlbVTdwDH/TPhejug
f4qH6wOvmIoRz/+pfN/5lJrMnFA1ZaSHBvtnyIz/SJdcmyDPgyF60+Yfh2BbGSd3oE134iFCLoU5
Lb0c/6415lTfyok/bzOu7KIK637C0n/aIlc/C0Cu42xs8Zov+0ZtywA0pJt9MW9O32zhwibuXSQW
iCsSBajhBg50t4Al61YNEm5OM8lq2cRCU2qQE4V/B6hnlvkB0rvnAmIK+nRWgqGH0aD3sUZh3SXy
rC34wZyCGi1XQUtkdkGi5dHUzUt5FarNCAgpCpsHCYm3+2Bl4ziZ40aI8QKiAuAOGn1I6f0mGqJh
DEMoxQaYVk71RCffX7HZ7F4w/1+zQqi507o3L8A68CXtFa8oCdjv3CM84moyB3I4jL3+J5S5y7zH
dU+ZFf/QFzRLwzWoFNHB2fyti3RVMht4qcy4pTrgd+3HCIqjnpz6WaTEI0A9i7y4gbljbE4Ilhgk
/6Ti2Pv12aPSuopr1ptiqtFinTESlTV18G74ioDaPcQ6v+lUZswNpnOd2Q25q+T9A5792M0XZD3A
N1qdyjiMve3nC4aVSX9AD2tzirayOGNO433vKX8LwFWLY9RA3XmxxCP22pHz0m2prMYBcuNSlB6B
Z1poJuJo2UPjIDAR3p2tncXIGWqGmFECVIKv/Y5krST1QIvuYFJDkd+mQxbgC7XVY3rdni6x+fTC
xtQ16NLNHkdbYeei6vu1qm8nBTGfHyTWwxXa5bs5wwUIVIgWIZdjMIew59KFKZq+04OMPjSPRseo
Ltsjrc5KP100unTHjC1QT9LQSrk/T0Rleus8wQLLnxN9GHM4nLMNJnJWPOiZFuryef9R5r4gPFMr
nr72SPjyzTZzOqM1qzXIneIRhi7+7fvgOqij2LwdirnKkaiQqGBPIX9EZBv2hG8k/xR23pn2QzGP
ZG9elD5e1ZVA1CRD2WPC14D5kZ4evimmJtZ5/9hdWaaJDPmasc3gdMmrFkgZIJlTwWWSnzitxXvl
wPvIJsE739bQ7f6jmDGrQpDnUj0b+6dfoQLxxGtJDiyQL8Gjqg00R23swQvp9+bI72XgPGY2W5QQ
PvXu3SXayenzeE9q2iXYSZTCToc51wGtWRgp7QtQ9XbkQDSvDN9tht9JydBZjO9qKTn49e3raCFf
7YcXpNtcUys2qJpozEtdLwoAKm67NJZEFoGq8DlFt4eB5unUi8iKSVyt68VLtaK/HYZ2HR6YbfO6
TjmKdud/ZnXu5L8cBvkT/MP/gLpPocyosexoyqt1JPAZc6+GO2fJskVxE5Wi91r0HGrmHbDUvCpK
JBMOGgKzrOulVvuimSdjixJlNTG4nLn9v4oyIdYxCMHFe2+ayF4mzAmn26CQgOiQDtcrw2JT1XMT
fwuJ/aY+Zzj9jLiW2o36/UOcbCBsd7Mycosm3q/okkaZ/NNPAU/AcEFO44UBzVkJ45n/1/EDXpQj
Usz1ZNCJdasNFT6Ex/j6okLUQlkeEXhOTlrYez3D6EshEdXPPbV7CzwNLBYfeTCiJZ+ihHLd/e02
Ls/4djX0Cpz0wKcI6tS9FtsZ52og7zprN/XN4qS+RDHqp2dr1rwBGJ2MGioPqISuBc6dzftr0t2V
b7oUl/ct1NQUwgixwC38+zfFmEV6AOz4i57xV3O8U+RYV7KjssynGYg5qndYxTa/604RnTpZjpdw
o1lgK/y06eYSB7KTZS9SzOZnGhz1dWo3HmxVHfwjgNsmRZBqSQLIr5UugWIZf3xHsELrB3aBvX0M
WNAJG0+GA9VHePZlM8U/ykkhtCsDNh6tkkImjhhno5mdda7buPSUc09WRldVJJ85GYSSMvETxFj1
nmbf03AcMAhVZrAY0izEUsYredS58eLcSeKw1t5bTAjJQALKfJltSpWpveES7lnV9PxDHArQoiGt
KU/NVLCg2xYr/f3wFiTMurN243/7nvQlnMFy20SlbrazfOclqYH/C2BXEMU2My77YLfRiMkzH+Wv
pHT23n3B/KVWyCuvYVvbDxrebKaveYSH4oYH4LrqclUbGfWzUxQZLmdJwCtoArFlIHdFSk8Xpu6P
XnAiO8+dTnX4OVnpC+675eOA2j4DS6kzYtxRtVnaM1t/jUND1HhtzBQSBR7S/JaSacoVRoTS8g5O
mQLU+1tkwryrrbIZ8pCra8i3aQqunnQKLOo2INA9Rsy4s+bqjFvdVCzq/8fN9yO2d/zcZLiQ+/Kj
IDjE4kH+4BFL/b7/hBwmegxkqWzvgawdHSUl705ans+V0SmUq4GXJI+EqDDeBVEwVm9R/7MQWYQU
EVwh/hKJWjg2gOaTW68DdBVADnItzT87M6BZv/NdLNRfYZ8MipKMsNkNXg6nUXmbMDfQeJv2qiAm
AfHHkeh2NN5I2zCa2z1WyP0gJ0zaSU4SwxIPtpE2MqWJVYx9D8rPZkntPj04pGlVXoA3Ybnvc77i
gUxzM/g8NUrtOHdqLV9QxxwtY8KanPTbuxzVve0YdpiA/A87udSpNthGPAdBoyirmuvtLnD2mHlj
o3gRE9aJllt9Fz7zD9g4gAIsMrXjvSBzO9vmvR+M3vSjwXmZ1/WablC43/OOZr6ooSjG8TACAcY4
ZAhX+TBNThpaOTH9c55TQ+UKgNF0l2p6ndaLlUPe6oTbZ8gK8da7CD8B/4/OrC5EWsSSzTPlt71F
6s5gPLhkcBbNev8a5oEIYHtI5zqlrAd9l2cZX5q2TjaL2laayEXQX8tJ7POxim3pSw1tftbM/cG+
I/18GnHfAUgJhTWt+m/J9s41FjVoeoWdTyq5qNA9Sb8I1BdPYr2lbskUBQP9oqHN/qKExc6eq+1H
UAIwvMM7ETt8oSiHAfxhIvNwZdDN4yLaO7UMPlkF+ceKZGxcBkfKR7t2V+UjVsd1VI4VYK6kGC4m
QDE3MenvDMk8biGwiqmOsWXyo8j0Zaql/NaPr6jMfBjoReKVUg6T3zK8dvDUfTBVTRfijth9FwKM
OIStdRuP85HbqTARDmVIj81iG8FJgI11cWAR7PElAamxx31klfRNYJA2043vL9GX7OjAk1+JZcSB
eUJfKdosLkKEnJIH/i8lrk/10vwqFPiyqfV6qFw1lKkOJGrGpU/m5PCrm0On2ykkSN89GSBLgkH6
QY6o7dOXLo70LYwWTSbDt8byA3PibeAxJdEQxHubRtXQUFRWZFTDcPZd+nCx1N9l61PY5wT92qZz
ll2Mp4zrBFXwinseUpTn17mh/R2wGpEfO2ltzm9s1Be0LrbapB5ySK+mTZaZv/RrWYI3Cx07BxKU
bon2ufPWyLvTS7hca+vv2PAraWJFQYyKafGbmw5xECHjWdnKAjmjIIlab+tE/cA8DbnZ3f2OY8iO
1U9thUkJK3YZyTaGGcy8JVOrbxAKqkGjMehU8KopAeaXfxo0S990M2K//LiCoS3w+q/TZ4DxgvZI
zLj0zTd/T2XxoIrrXYkRcWUPLiwdj331tzylJoNCM78YC6p11hATfsL9r0c3wUHndKCk6Vz7AFeV
4it840EQFU13A7mjJtOKTj4Aoe17aqJYBcp6qMggErO2MpT1Ja4zIKerIErySTiFHY+QIn66UAZE
g5gdtX9oj1MIvzMHIeac+FL18ARmCMbdhoqs+FhRlhWrv5ksqIqQWgcQTbfyuy3bTciSto0+h9Ge
oxtkFKNhEhn6PKJz3QP3EtWgTT4kHxLjsoFZ/02bHncez06fY0EcnZg1fZqp9aUh+SZLD/P69QVw
RHQmi82dciOIWsrlTwBdjbWmOBISeX3o0qqhMJ8lpyV4jX2pLU8Xbzy/jldc1yAJ/tZihRHrgO/w
XDaiU7OoGPtxLQQNvW8S8S5FBe3Zp+THaiyHgwk5sdLSmYi8S+ROksl9kPJP/nK7T/7xwFTDEB+J
Lj68SJlWYN/m7BLzpqIqYtm2/ncINW/JQwce2RAKTZSFJkUpn0Ii7TJorPuAgeTMdyiUMKtv9TWA
TB87umc3C8bl8ZubcKs+L3Ef50lBtfxZwuTKTnBLa6BIa8QYzHR5LxzcD396BOmFVNiSsd1AiBCB
jcQ36UdXWH/LUz7CIO7+PE8fhJUO3m0eIaxed6wslmWUJrt36+dSV8IGNErriIZIOaUB74ussFpR
z75riCf+qVlm1t0jL934NNZw6f7g4L8FXKxXNnyOXlc2GSFYpVcm6gZ4xq1RRaZWHmk0QP/KNHlf
K+bum9fFPzgOZK97ATJ83dxRNmshobjDpoOFYtk0qz3X0l/1raR1qNr9GJLRF6488/U0tAONteJk
FGTDmQ8vlOY+vp3Q7d89g52AcxI+veTHbYYARQmxngXn5ExMuenB4h5ia4qH9P8JMN/Poy8PgFB+
WW8G56zHsUalxNgkgRsv1x3IQrmh8IQo3AWwsj7da/81S3ep9kgCtyDhLv7LQg/2HsA/rZgF7FBd
Z2JEo24IYaMB4LPB9YI5MhcF75gD2eYp6SuZmZ7yRquqC2utpe4TWTv07stb2htVidvTqGXqyZMj
FYOygVjfnfX12UavbVBuPEkECTnuIkDLP7ws7CYCcIGGHft3iactALpSF4n9oiA/AIDQfnpazQ3L
Dk7NWdT3NQqNetkKUFHuyEAEzVxSn8l+iQaLt36bb9uP8876FPFsLYbtt3h+ZPLtTGtePqYOa6qV
Elu84pMnowezLqhHaAvN0MpeAke+Zn7RgDx52N8FpZTiWYaThWJAXxs/9zXjK9Nv8rkWEyRQJb5h
i0i7efkNT636uqZ+aUt/cigdWzrkleo1D+CIyu87+dT78QKSiVU2S5yuTsMt1rGKwwZkEjEZPZgr
Unooa00A/RxZnbI+UDl16x7yKlnpU7c1TUK7ZQ7p+yUnVq6MuM4M3yqsrwlX0k8GSk5Z01Ud9NvZ
4QSqpUpU06NLDsjXxMAvelzF85KGTLda0logKyA8iBF8J94VicP6CKWUbOSxPNeKMn6Ih+qcagOV
BGJpqqm61pYzQA/ZBkJYdpUpidNBnPTmStz7zIlYccwb+dNliazdhQvYdlibEyKrw6zlexWuHMas
S6z0ogzbd0K/aUSzxNxz70m3xVX6ChK+NPw0f3PtiRLUlSOFBWm8UptrBd1X6erDG6uMd7XSIEsS
xnekWCiXXXxWuBpJSfa0UrN54YIJvkN6998mMLwBcM7LESh0ZIOYEVz0K5mE02NA1QijR9+LlXDq
GTLtylENn506Xr9bfjWQbnHk9SEjEFDUP69JPiO347c/lp/RUz99ZlFXpNtluDfBKWHIzUsBn/lt
MfB9cH32JfqbbfNWGRfLv+44YAEZ034PmhK4cVOi00KufzmlmR6QNv9rUap4YBV0dj96W6jDWuGF
seTfuCU14VwCiWvRB9uF4dsdXEHhBC8otDMxUVrMuK1nVe9eQYcbJS0o23QsrsV9MIHWWf3FH2BR
KCgUDnnp8bOujcaR1z8bxpJ5TKgiLIOeBouWuDJ8uMcuCCasXw9wtm+EUdHCaKk0OjA+wNLQiz0I
TSPLju2putPNHejdvT3AgmEpSXDFYHnMBFTbCBSfXbzX6CIaGUILxeko2F7v/D8okBt1elLpXZ9u
TBUePRBivTe9tEqZsWBhIBgO44W7B5VVZRu+F7fQQHNCaVR/xSqdswXb4tME15pd9rCH/YWPFFJ0
pe8UhDTorJoHbuB0Ca+yQ+GfP7ljTrqwc2nee9++ltCa8m1SE/qn/VP9rayQ5DpNvo6FZuq5wT6z
bK3Uf43gGBBDX/GMhOtM37bkGro2mwYlQ883DL2tbqLXTMEouC7mAIf1QATRhd7cYglbcCi5p0Af
FTsb6Ch/g8sc1AfGjATtnY34Rs4NDdaFFC9o2dz76owecTbB+Z0B7ucTXe9f4afrnNM1ziqbBuHY
9Of7Ru3MnqiINC6zkkJoJ4LYsM0DZfZmPwXu2Sa7uAnVMzQtL0nkwQ07ZtRml0VfAwIZxY6Cw1lr
LN3+LVa+vOLsunDk5J5VDw6jQx5GAIFnmS8ZXGSeJExfiuQjSBeD/OWD7ctxVzPeqEJvwCYPZRj6
CC2AEmUD2gtTJF1RgToGVJRnI07cg8mQfaVQouO8I2/3UMqBcs+sAOm5sW4ERjt4JFp6DymiXQXl
aYjqS6tZPa22lRGu3mXo+7Rh7iCygvK/miqwsNuQHgdkdsvT3Amq1Al0oqlbT7BMO72gzHsVJBiP
SWVB/5xElEI7ZoeXFFr6z25eUr8sn58XyifFJb0hCoziWV/6PZgPyqE7diXOOSRaaJNWLVframLN
Yyy18ZtxQr3MpmBh9sae/ClKtZ2gYBV48VyGDnkfW+Fyyu/TxK064YUQGxY6OF1yBR6EyfYJBQS8
+PA7R64IDExzv9cQLz9aDNhOVDPQ+dbpSfyMiGQXHtTjjtpCERJ7ayjGOwvRiB8kVAI+47uHFdC1
rGD3xIMrymE4D04ruWrcUP1BIiJCKrOcfMD+AP2TpGhHLQ+3Yakv5Bwp01N2/1KdyL52Nd1QT2OR
RfhLEtYv9BmJ8P24eKd7Fk24AScTeH9PP99jEdM5ZBNJpOk2Wgji9rdXu+tGEfMn4bluiJIVBE8H
73PcS4FKjJpphhHlAY1VaIQkvk7kRFUyGqtch5ZkPPHh+xbIAqiesMGpTKbFugu5m66IcbS3ioO8
ewi5JrbCTlWgZVMhW/lprN2XoAXnf+Y+jv1ateXWoa3mkPk5d6w+ONfJRzfA+G9Q+rskqfpe7e/5
5ED8z2ywe8bFQW9sUZxS+HlsqI6F8/xWxxV/+c5i2qMjZLEffGTtBmpylX5w51wZUBUoNLqrqu+J
VK439OhEf7prZjpZ21DcegKy/R13b6g9PAdIlJgr5gGu1Hf0PzfQNnM6oPBUW0aiDviCc/YBTN7t
+qfhLP9wstFWqtrj3mdgAsT1fYfwimq8jwFFH0mMjfl6p9cFMVPzxgUPlfKj12dkTwpfR54DfBsF
ERTjubT783sYpMoPf03EKC6wTxqCl0HiWRfxJYaqRCCoYUJ5FaqKlJ2eUcIH++2shbt/yRaHiXYY
FbgLDhXUoesd0E/dWaMKoI3dm0q1Lt7CWsljT8/BwKESn+7y+miuG3duX3kqDlSq+YrPRf0J8b38
3UziGe82Glzw3cFSAxUlQQB8eGfP0QjEd+CkClHn22XWBSUtNA93me0h/JWXp50veRLrjak0bq9l
e6O7kr9MnnYKg7BBQR95h/4ge2kX40NmChqUW4ULDVDgcnnUvBikkpZg47u9PtP+pSgP+nBz8Qr9
kf6iDAbFH2bpN2g77f2hTc0pNrU1rNir3DvInH7C3WRplwxMvlDVbM+7E16Eds33Qme3k2mtFagp
vbBZQTclY88OXkD8IBzqmymIeUV3eOcuXPbGJ+Mt4PZcDB4uSv0hJ0E3/iS07UJ8ygbUgKeruhhv
TrhXrqF0J3TmQDuyzfD+f1i3cEslP/709tj7bsy7XddoL9KUWu7+SYitQ335HDIYFVt1X8OsEbjk
zicbehP82Z79xlQXYWGmOjuWqYP3aWT60wtYkMh3U0eAPXUn8e5/p8FQuB0TQqe+1eUFwZdXKFdr
Czfc/z4puevz/H6WAJw1LAkUW1NdcuKvbcdeywGw/XU4ctw2dTWXA0dN8VXQxfWGsy0Eh/sKYCEj
YCjAwYA0u1ly1c2JCBPJYcD0eN0dFs7uVyefg+xANxLjog1nus74TEG2+AXUU0390e/SafG2hiow
/RqZsllhPg5074BB3QgoYfIRmwoVEsKc/XvI9yIRRCa5PLL5ZY1ALBwWWirLcD9MDEGw4RK6jbYH
h6gL9iQniyNuPhdgvfgAWqpw7EH2ziXgEBWbvGfacqTZbv3MdooY1wlIuRmgm+LGLV9mH7lYyvEh
ty+fHRp6EZp+FWv4X1JfKWlOZIZ7/qbT/m845AY21ch05auyOiR/2/nO+AHZFmMp+q8BZtxE+Zmr
T1faYZVVd/TNVRAqPRpHoqEisSipCbwe1HvQ3Ffu6xzmwG0rUpuOEc1X5O7bNM7r+V5jkPM3gIxN
t5tkjYgfb+v0XacR7rgD6sP4m36yLb+WFnc9YWnnKoZUbekWmHHpHOr08Ca8yr3ieMreH8FyKu6o
h9vpNOQCN5i9ttKKmHoxmLTF5lobkbn+v6NWvL17J93/26yZCZQcYByhgigh4cnAy6YQkVYbQRHE
3C8z78QJmLsmyoCNexJnMW101OeHJntRfgR/FpgWLejd72kfXBf3tEB2Z+sqxjG9YO1SDiHjquC8
Ls+Vjr//atIOUXxLhNZ72soUFFzPyEEvaOTe67ZQ30EG3ORb1ztIfB15R9lZny1PIHSkkfNkWInA
qWMgNgzRO/9/GNKS+szKQai0peuflwq09m5ryy6JJrsrSLnnfWWc++MZBOeJq3oCEonhos52kDmK
bZAAm0h9Dsx1mzPfw53FxnB6nqcN2vESpcs9nvA4oVnthKzchp3XjTOk+ZzQZR62zz+pQl541OJI
S+eKXu47UWng4NKcn7xinpoNmDyd+0VG1rLCOw/Y5XzaXACEQAJ5+o0oKMs2mhvUOFaHfoZfCLXh
FTAzomQOisxzkG340ZQtH+FqCp8Y37UB3kmDFMW03tMBZE0BqJ+7fi7W8b+vBeNbhkcZdJfRmeas
mxoymMGu4cSY/u395gfMTcLi9Z9nCRm34adn0o6vE/Z/r4Eh4zBe48bz3zZ9za1is3t45jbeQnc4
alyMKCJqdT9n9bcuEzp/5DjjknYwgZbIaK3DkjdcphnbRXXuVMQ3d5hiNlFm2D5opz3ROC8bnut5
eSrwavBup3WnKiwHo/1oS4n1VNP7ovTHod42CTj1DMbNfSL+GU1NVy1cTUJD7E5WMxc/5zkv6cOg
GUyOasM5IDVlnxX+sNno8ZawmJnaZ2OrMC753FMafaHsJ8h0hIvbbgsiUCUUAJI6zrtLeTvymogM
k/z/8BAXsxO7xm5ba/SusSMMeXyCUt9SXuuBZah3wugVZXW1DBHSWkrOrRXKdD8NkiTHI+O/sf1o
Nb20RCA9Yq0h8fBRpyLLWXmKDUUKSVm+TEPNoi9MXQtuW+fvS/HACLe9jDHZoSbu1ykgXXUPiUUl
/igEziaIzywhUv66rW2oqscIpoRtfbauUIpa9vY+2eS23bjtTPz2OZQC8mkgXiMl6+V5aJw1PY2f
UXn5v9mumIYptb2La2tinexBHD37FZaL3t6c3Wk1mtqDHAC60GjhuEofDfaCJSCEF70PT1Qkkdt9
p8ZvXx2P8ptJE010olUATfFzQ6CG/kev0BpMQf49s8NWVTdxa4EugLhuhsOlqIjPyhd5XYNCdrrk
D2kwoNjuXZPeuZnfjX0cEXyrqnFePd+xkPd5DizjJhuFuvdmObuhsrVURYQ4vHjyAp7cjEbp0+GM
AaQne6AkLa6fvMmNiZTbvMcNLdv+aZNcKURIsSg+A134oMUOysiFfHF4kJIctCietVKug+GLZP38
srnqpvMVFALNxTzf6bxFYrRkhpK1CJBF3ViX24uBkUrD+BptOfNItqLNmj24JkKxaD8uRc/urlpe
kyaap5pOP3te5nAeDDg/pHvmytKU36AY3krpt8ud/STVHVEH/pMHrFzyFmP7YNucVDs9a/TY5HPg
SnZsGbzNHEOzxefpmkIWXsHaMscSTQvhIIDNtMppbAGpX6AUMBEMnAljXufySWXvmovd0HCV23SS
D0pWoHXGviNs7ZU0kBEpggnMCvTmEOKHYOel8qxn+dwiDiY0Xif0TE6I4GAkpEpZ0BPOuF6NS7Ek
YNgVPUTdtmFcsUmdbzcN7QM2bBuOFwealZW3YhjHGmjM9sKFrlKGT2Fyorj0JhMrJxf8bYfPwYAs
O9OH2gRZwyC54JEzzKIcBS+06XwaiP3M8DswmPST7WgDfexRrnzcGgUlKrzDAkW1v2V2sqTB5Etc
7ShUihtX7lMCUqH0xkRR/NK6m68nPYGZNijU9G9DqkLEGp2X3gsLI0NWzRCafYH7VTO7LnyFCfZ7
v/l0PlUjBckNmQl32Y2t9aCPaEcg/CSNMAX+k03VToTIC4EgBF7HdDY8TFqcNE7cnr6W5hpnDcEn
iQTFw9J5iAxrC+0Ki2lkJVj0Rw8h9/bSpjnJXdLnMNugVyIcRTuVTsxCDWQaVVM8H+DpdAG2MooH
Ei8Mug1j02N1xZjHYk+pxxRc3aiSKeUOIqmYW7H6l8Bn6gkjZqdx4m6gOte4pi63lfgK8C2eneAZ
kH1gSd6UzOsxVTNjwe6hjfOIv2+okpq9Yv1MXJDSUa36SUh5VoZmuhvF8tfNioRewAGyunDFOAf0
6pJCIWX6SPwK8rL+LTImS4fXHj62TPsUipJWmEElYnjdX6947BBHSanDkrsYQqTy+C64zlItzm0I
KrfZmVlY4lBavbWkl3+WEy0a+WxrWswIVSUQpZSPjfg9cOXCJcWQH4ikqxIPEFa7pC9fmB/3cw1g
PXGiHunEW5OXr/uc+MzMefQjlEUApSvwAfn1J2ANcu/nEz6q4tzm72TlUmzY5f0BC7vgGzvotj79
Kv7G4ViYXHKi2zAo1jj218jegmy5t3j3ywWgzgac1id1xwhHCotLEgq9MTiiCR856ZK0JZPZFCJV
eSzb/pOFkezh/r5OF8iyI0Hj9ElgGhhyPBQwzQ9mWExaYQ4FB4VD9L2eOfcjXua4sBak60TZUkrD
C9G2UH2odU2HCwPuPMqYAJ+I+jrx9ytjQRr/iz5/JfMDFrNofsAP/bsBD7bfZzg1ME0oLY/6E2qc
TbttkrN5Lwt0xs2rHlOJF1FlnyWZc0l4JZFqKuEuBBNhzXouM+TWXdgHi8pRAgCeErAsQOTNgdZ9
QeGtQ1nwRU8YlenUlWVqMsgfmtLeWrq8WkCArbXA4WuRnEUj5KtypECNuVZvs6+H4weUiRmkg/ax
fDn7PUoGQRvh4LBG+l5k6H1VaykUDajl+dvxIi5U0zt1fU9fhSfBB2nFi16fKkwEri+pQpZH9Lwj
FmhgPBmUwYY7AwloCWDk+xZGh1/5O150wXXa+s9vyIzKHPVyhtnhNe0MHKD4hnrAZaPTWHjzZD6u
vC4GuZ9I60b1KAoHyVBXFVUVHbeYl3gMjg3CMQr38cM+aMpmrsnFtVm6aV1f5in+zjZKoKcaaUu2
aq5QbJaiaFGh0PJ506rZlpNF93eP7QnynCp0fm7KyWqGYCaW2lJSuXUuxODyU6Fr4p8Ix6Z9+xpZ
8xpd+aK9jGaCZGXu1bYOsPpIP8JsS7bLLN68WqwVYhnXVVhG/r/JmMOdDOHty/Qh/qiW+qaB4tbB
gl11Sq6rFlVzOGVETKAS3FdY+wFiI3/tAvU+NNbU5ZwXc11HRkBX5TpNSWqMsjRIC6kCuDJtWa+3
uW2DwiZhUbGItbhoZVISmd0gYvqA/x879EZzBHCILzNt/Z+vVLKxNehr2+of0HDKWUksNzl/qdom
ilJWfM7aPNNr3joIc1j/Hifsb8wVviYbfW0ls+0NG+JrL0Rd6p/cFz+pGovpaSxEOtVVAC1kOsnJ
l6Yo1ZW4NWGQYjmXF3f92/KsjvFIzFm1XDmOXragvdCqZ4jsB3XlRomNweRlzKbQfqOLD1qm8bjX
OSHmtBwgz3fX+N/6rHf42KMAWqcTO4ZyRY13oU6ngW/AFj8J4+ePPTXvSRf9NyTTBQHnExR0bdYN
Q/vH5WaVkk/3x2mwqyd/UnGdKWBzP/nEdRQFPH9dq9e6gOGc4weA0Pkty8PJebU/BK3qxrVq/aA7
7aIo61ph+uuXE+VYbvLaFEhxT9bkac79LIJUalF2kBwkKa2ZrtCJH1lSOa1LRrQbLMvwMTMZvEB1
exjq1wUHBV0D6KYTdnSJt9g6UzMk3YDOVbiZnKLuQBwCTQnycs7AwMrABmloRfnZlsVopv/yCkvr
VZ3hxpcdv8/t3xEd7kdmNu+dRAWUqiL+OWwXO0YuMSFxXo8JoeTHwGKdVKopLlOXAFf3Y58U77qu
/Z2Si4PtM7GLedz0xs+27+ehyOxcnUrj6gsQYnreGZEC9kCPY9SpkOIYHJVrQmaxdFW3/C3JGEU+
NSOjk4CcKLHC3CcwW6LFS5LbR+D51bo/5XpP2gKLjk6lj24lhB46E0sSdO0w6iFsWhdtNiOkUmea
srt4FbZtP++8r1Rm1mU0Uo4CB7bSxmh2xob7Ejg9u7kKd2I/nYX8Vb2tBFQUYWyDG1b6nRnDU41o
UNgRMOiGcM5VvLPwbI64CbjBSPTU4d7OJvAHvh6cMswqF7rH7+wXM4LNylLcc66880ADHnVPKCLX
5QW3PUEGUcQfbtKS5LuX+lNXAJvDGIdHzqb4iwYXaMv41Hy1Ypxc/9Yo6ugB32dgg07/ZGKPrNIp
V8qkvMv7V+ohnv/YVFkCJioUXBY8429Os1aPBQ9BXySPv8Vz+l80aZz7PsfizP2rbcXbkTu7rKma
hc2Tn9/vTGrbQC4JDCQvgktsumBEWRQCg2F/QOaVU5PQYng9ZaiTCjA96pIqCXS6yHer+GqPzZxv
SgQ+5KDhCUApcfrm/XVr+Hqnx0pYySba7G7Vt9Qw5tWJ4MWAIB24KJL6J2FoGTvA0rspQII3i1Os
fhM0OIU0mulX9FTrRR5QIQeBdyxjS9fJ5THX5t4SE0Fknr/ZFMbUeLsj3pBHZqeZQDRWcvkQYhpt
c4HZZ+0yTIO5c+TYfhQ87UKurVjlrLjY/Os/bymHgMIM2ScCP2XcO+sr1hTdcxn/qOnHf8qdPNQt
5qlB7wbNLXEOFPzz4hHrEhfeEPvvuoBScr55BLpmqQVIPOqMRbmbQ8VxjLLUyiUsrNiZGIWXAaCZ
kxGVFyNPpg725uOoN1vGHnmuc58/MjuE/1lGqgJPTAW8Sv3ClPkvU7cQv080SAg0IZaw9gVYwxUs
IBbVrQ0FC8DSYxRljeCxIOoH6Ih7HR01t+HbRbtfRbMNWy2jeztmB3Mg6+nOO5C6mI2hGKiaaC2A
8/TiVkRDRgJkJM54GjsKbWVSPfcl34qqgqKhPj/g6TFMTIx3CNhWcDvMWG2mZUdbN8Wx35/RUqSK
95466oK8Myacq2oa1NQ91v7fkePTni1XwGRKfjrVROGkebfGdvIY/nQxBObCDqmlknyV2EVFIVGS
Y8dqhovpfYN2QFKl2SYSd5hk8ZIUJHj7aoB+lOJIa1bsPGzfVJ5xczxtNCnpdcJYkQ/eGjRFICal
iG2H9bMYzwSTPTG9cdUyBst0w0XC4EKPtAJLDGx4XW5sHpE9xpX1XzZJLSpzjCWKaUOZMHsdyI26
L9bssY8k8v/sbeFxtrmGMjHPB8uEcFquOD8mq1O3xi0G3c63HgYt7gG0CABVwYUS2o2u9HSw1Qor
BlkS8JaDHtLBekvTCDq1Af5v87HDNJvVEByXDDO7E5eGijXOsHnC6goeo+dnVVNL9nvmZNogM5bB
El9wOmvcLLnMHJPFdfTUCejwIQ8HDghgcKwJ0zZZu7P6f++g3SeMNMClC/DsPboCAbJOIMnKK+ur
Lg143pZb/bt/MtHbOVJ0bIJW6OJOvFfaHORP+oFxfveC8Rqgg+w7mNz0Eo7v+mGSQFV+2lnLUl9g
b/sslzOwfO+NQv290IVFNU9+DNa5umrDMjkMeS6Z67uVnWCTeOEhiWbo20sLc75HgVZDf50O3B2D
+7dFSO5rD3YVK4lrADcXNKTQAFqsPiXBq+3EIi5kcdoKa1/AQW+EdBtjog9SBwa38+TGrhOmfsZ+
KRjb5pIDKfZJ4g496sXPRxK4utiiQ86XoGfVqrdE249l96dKbjGU9ISLdd0ojk6i02OXPvXS6AcG
r2ITMfori27HdM+s574g6bqOpNQGL6N9fWXcfNCwOvuvVYcWMKnamn00nbr3vSB1qm4zgvh3xse9
4umzyJRiRlPsMMbTEkn/kH6o5fBlTJncKZOV5o3dr4pZM5QN5UoaU6QAYQY+mgXubV0P3a7BXWvO
6o5G0Ix7BV6U1J86TDpOkNwyRX4y6rULhX2WEAgfq7uTYR7RU/l93PUdE51fkDmBvMEsCJqioNnJ
tAP21k4Lob9gl0eYQYHSRFcIbitayZrCIUcYOvGYbkugfEzeUJnLK5PUppgspITZsUuhIdgQxlD3
T5vZeOLZoTJfYjoYv0edyEB0IRwsseM10Feb5rAJnz5pPXB8fKN3vNUSBUjgwQGE62gbOwAZbqCL
4igcJtzYVv53mAQtcCNZzPOAVRW90OT3FPbbr/JBau5aCJN45dVDSSBykoe+cUuXzAI5aXBlecUp
LurZrfLd0fsxdPAV1BvG7fwZ5+x9dNHPlc++mZE47+DcK3/ncaMyMa1GrZAdCX4C3NU8IMCppdUL
At7fjyanR3z2jpbVykGChvXumS0HwwrLVQz0uBIGVRMR8yO0OWxxkVpYogr8jPjdA378ARfBedfu
sGykAiCo6aI2BjwNjC4MDI2MiwpLwBbtlqPqKQzzPL7A+0XzhzLRNWKSNXXTTa5fjqRCmj2eEGfd
JJyJ7C4WSqNsGVGpcWwXPvyRxhknFNIkD/l+yJ52UVLwat0idwAPRSnwVJVZVMYKst11uIgI91uJ
M27CRD+3iJU6ON3E6FLKRDspcbJSMGGGiLGOclkc2R5aBp5QsmkV+la6V8u8I7qKGIfmjG7rZehv
u0Jrr8R0/B+USzCLC8bIvb/M75xuemkyK0r/0fykafVmm9CSuF6/C9wQSkE+taXDaJsStguB0xMb
fPbbmddhnTjjQ0VfLImqwlxF6CdlTPxAClCfdWvgvYh/ymEBhPDXs39QdUBPIUrftvrbN3jwot1P
PJYPYbtnmv04M5A3rMgltzP5Pswt3oJE2owOa1R3Gc2jTRps5ohlss6lv3sGDpBN66eY8GyzKR0i
qDI2/fEovgsI5TmQyWZn35R0YHeMeiabzJSTILnUy493ll0rVRH7s6B1mKVBi21eXkk6qHz/a98n
ENbq6fAFhM7pYr/F6YRx4+2HTAzKJ4T/flctSlmkqhaCaTCZzx/WbbJyaSM1xBMMpD076RvxgYdQ
jQxXNCMNRZ6QJ54wIuBI9mA3dQ8g6v4cxi1raJq/todPxfLUkfu0CSKBjoKzQEFAzWTlXx/PhIz+
2GcvDxwjTwd1DpyRjuLN0mipD/qdmqKVjU1D1rFpJDFzI8hV90jWssU0J6RLzCcE2vzu3+Co9Urp
+iBT/KYy9ylzCO8YEqD7elHmP9ZDHreRFwE0EXVgLrbmmj1qkMbO65rfJBTq3gKpNGpPnOLz6aqR
ELtfSld2ZI4Nlhutl77wdLkRd0sYnWEavz5BnjRErJcOkFhKyweMJ98/0xSKcVtd9d+jAtNaMknD
/6GLUwtNYerSdJZHEHGbYrcNYqzrL0X9ZEMas0mSQzyGbmmhEIiolP/fZrQa7KNFlSx+Qy5JRlt+
9I832nBz7ILk2rh4MukIRn8urUzlo/Kas2Hg/cUPGTPL9JuCp37aTQtnLB2TA14ikRMxtuo7amKr
FS9rua+uf6LsHlFPz+mogh+BCsaXoNhP4MEaUHJ4I7R1H9omWEIYvspTxiPFisYGWucdUR3EqoYq
hxYmjwQxGsDQGHxMcVWkTpk5Jm9hfj/hSmoyeEnWvlIPaSY32PW8wnQ9TwB12+IEmxLaDoXEKqWU
8z4r2Sk20nZ5o20JAwUtjKKAi+na8MESIz+rCT2nfhOYmw2XFaRm1AjWizg3mZBxLIXjAlljt+fg
lTtGX3kDi/pwsosdnHBmfA4+6AJ3E3k9w3uQ2wB0ICo6N7ZZHz1Z9x8x7TaWvxR7r6LcPxSirNcY
qCxRZZePETtXSFIwTx8kib1V32PVa60etMZFOH6QKJXJqjjNvAsErWqTRMFA9+0c+7KwA5yhPJUX
3XKmsACvhAqIW/s0iQDWL+3S+/+Qo7edYJJ0Xlv7P2NsBJVKasmDJb/KWGd61KHWrGzP3obCpMVX
T+4PELnsZJxzjojuj2/DM39uGgh7OkV765vnmZC4Ily92MamBUAVFQ9aP049k6zkHG8xAFDJusSA
vjDSu1Sg47Y5KkURugmW+CyrQhrqlR++ncgDxmWlHYt1Qb1Si5+ZQrAhg7E8JuhGbp6BAIfPykUJ
3TWipUfO8AdEpwOehFnjGbG/ElXoLLF7mW02nLp5AktEFG8Q+jeGAGzuUnTayA8vwywCv0vrEzKI
vP+pgAKOFb8RENHIrCs/weIg8MKNFi0JWCwbEb4YCg5mOWAHaZkdvL7laLE5KUE1cAfUvZA4BfV1
/1szXct3LKdhtd+Dt/f8C1k5xkYj+VJHHdTWXBFVGR65gsyxb/DmREAowHDIEtBWvfVRylw1p6BG
cTklD/pzMNBh3EtfAB0aEfpJAwp/6C5YBzFQAlZNVsVDOiqGdRUS9bLcZ427DILzG9UEGSZjF2o9
+ervJ6WDGhsrIl9Jl/ZExDOA4gYK7ekefslPu6gajU0Eq8KHBMXBDMGrU6dWMpGKFPesAGcQ+HQ4
56O3IoCLgQDFLloKSc9nqTzPD4g4MsB7Y34jOYYaTUcHR2IxmDFDguOXu02YbRHd/EHzbQ7JTBb2
BTOY30B4FKptBiGt/PTVVl6ndbAZFHR6XEIFCJlRQjC66Ohu848Iin2thHJRPIXSRDsLljs2pDQW
meFP8mOS0IuQsKFiV4j13UF7jIzC+E36lXW02baNWCfuCnK6N2r0paj41KAXjoaLinmm7Fl5R4dv
saodAhdkmYsnlpR6XmcXGNymbJBquq7VLV+OO6qUJw/npvWl1LBO9bbqCck91OoXEkT5X92CCZOW
yNUO7YAKpkps9xGONxFmksgqVjLryba8IfTbEF/0bLFuglEHO1NgHZBEeHJSZrz7z2ghCZ0s16Dh
B3k3709DxvmWsfDsS4VXP5h94fsFuuvtZnZW40Lecx/YiMg2RgyuuyyrN6BZOw13xBD4XT/mS5el
qimc301zROlkXFN5PqTaKOpMCHlT3+VchCsQJ682hs2R/DA2Nb89iW5c7LkCZCq6b2B9mo33ZVRM
ZSilUNKcamKX1iGiZ4/WCk/vlGJIXaLq0AP4/Eyw8RXu5RQZtxTnGxL2C3hDjPF+0OVL+BMXNn2U
opSgJI0QFFfyir1JA01VDSBE7l4B8g0CQABuO7rSR8hX7dSgt2qxTYTdphgvkpOIzZUOFfFgs4UX
tTUV1g6U/7KTomjRCjbWHqQLSWZXiVYSd/TxoarnHRu4eouYJI4iJfsJZYgZBuh4OdRie/0YmNjn
ux003AANsGdqFMe0hCZbkjJmIKc6vEK6UJCdMDRBwad8ZErKJX/TTOeSaPw78GnZSZ3QLDtqaPRa
oNSa6n8ogh7DAPkK/zza7T/dkBcVuw5TEZChYryCQ/8rxspzVdi/x2KG1lifWqp/Kt5O3qOxshMA
4zeXJRcX6KxkCdFOal6QkgMpLQfnJRZ3TKSp+7vJDoXnHRY7EnzwfOA/8cWcAGJPcxu0i/BLS5iP
OAd7FkOTsJybnX6Zt/Z27ueUxssXkeMdAPcwhHcZsNJGN4TzXtWxGIJZrI8LsJ8j9MqK1CVmOLPp
sGtSyuWLy4ChCrY2o2XuzTz4Ifgu5POkrGe2knt6vHOH5G9ZXZCk6GEVEmmYN8NmuzjaeRe/l6mu
v8CXxkHYgy5GKzJ/NyBn/xtbmfWVDO8SENHJ6KKZv6K/+rIsqW5vSwXZtbXUWWXgYzw0iMFGY5I8
aNoHplopXqiGcWv3YVWvuN++aLqVz17ZhGQkOXlbf/6gSf1SoUS4R8J88nmX0kNRTjlk84kknlbJ
88GNPhfpr87M9kva3L/lTTcQftwwsPoXBDL5vqAj9DC35fiFlsrVajWi+6c1O1WOi8mSK129cJKf
fxDNnrCmolbngKMWaleBvOQ7rqbncbr1gAi7/tz1RWo491MTrXt7a+3sfd60yIvNxDNlPMvLeKtE
pXtEwuagbiBeEI/3u9lsJpFjPPPPTF9Frhjdq0N87kLgsLcSRU7wimGgdMLJ4ty4hcxLfkG4J3gR
i1V9QvS2eiy/IDa4N+ZnSrFJmKkhDpXit7Lyg9JalVwFIF6YPWygfjIsqgQ+nFaDPn9q2VuI+eSU
jSGZIdoUv7Q5rSHUbmXGEO3VLkTpjFEf1Iqnv6oxUcJnQUO7zXJksBIyrHVj291+qeHIdwZCuVKA
aW3sd+lepnSS3bb6kXNv03OpObC+JicN0IX+ny85mThxc4vagJUbM0Gg21JM/uOArN8Q1wY/QJg7
UxsjzBfY+pwaq7tBCcv27rbpXCrMjxORxOdY9x0+AmSFeABn/i6/WeKmqsIrHnD4bKo/Bcon3hqr
w1zugyexdvbgrV2ls9It79mQ6qywyy8DtV6o+0lZh8onrQsQIwueBDmeK1j8+tuDlnVJMWDuNGBa
2vgik4ZwkCK1IMj/+kxQlabJ/7An6/j1UbzgHPlN2Zsa/FLohzZXCf3MilF+VWjb+Lgh/ga9nVcL
yLl0SCOOHehixPTC8FgzegiM68BTZiYWBriOoeCk7deCDxqTpEvsYthnctnfe/JxlYAoRPkzTRP0
b/38Wb3ZJMG7+U1ehjmw1EciThNgFMBSdmF+NIfktyei73FfXp2MXdNzckvbt9Mf/1/fH2+iqMra
R5meRqo/i1RTRYfJ+Yrvw0NU6pZni7Yzg4s1QnLJU2JeiqKPMTd4iDeahulo/r5GYuDYqi4GR0L1
KyEz2JXq0njn3vpO5PejVKVyfbkGoNc0kRKDj/zbQ6e1YDEROhO+xBn+eSqAfWNUyy6UZjbu40DY
xftBf0j/AmJXclhvn/339yqVGOaxm6nPOk1v/0q3KjXPcO44QybioRmKV4mcjk+qU63T+HqQwi53
AX7ocl5M0y+rhajQ7FEm7ntilJWdbN/01v2ar+VbQPvNpeaoMBBZ5cbOAdCt1R6ntEVSRF0v6dcW
RO1qRNv8TVFv0qPNStp+ZoF2P6F+DrhhqiQ0cjWBNLE43ot5D08qECCtiQOSQ3qq3cIlOUkQZYhq
8pq3wwdTx43Mi2KtQlDtuIc1vRzHibr2NGdd42nOOKAfF6c3p4fgrvdO62QnjOnnJ0vcR+IGMbT3
ZDKBplv1DAjyNov+EHBr3xhxCRqPuu4y1AFgU+OeHALxONgMsQnJMxp5aWkW+7zYm1gToF3FEYIH
My9G6gZZe7orNqOEUSXxXl7yib9U34OrGhbtlLBB6M2bqAT51fr9BZu6apjndgJrYPRecn0prwP7
adw31DJPaNc1qGD9TxPIPvH2F01QvjVedBwhUX06aDH0BJK5w6+ZFoPHl19AWwq4S6vuPjuZ3Sq/
IUzBgNFzrqKR0xeLQBRPcL2RBtXYZSkGoS9v4+mU0G2g5oufNHbwfldKm6cfBLUDnL5rS8F/7Ypp
SUcSV+EtSNi4avBsl5mtoIkJ7wdrK0uPIYInKgkYG2CYLBoAOuRmMlAmcxNmMWSgSKhQkjSqtzXR
Yb9Od9QwL+N1Gzab4qsVsUGxVKmPLLH4sPZ85qGSdZnE+Df4/BQO+BGSYpzzI61AV/g+iG8Cq+D9
aPniRgy8Y5KW/56yZPgdYLB8lNRAYA2IqADp/FVIwlrJPcF0m/43met67oYnSKERgXcpvLpIgC1R
UdimL+Swsr3LpTBpateeSclE2JvCWtyukAlaQKAkPNWOfMEFqAMeqgj4ihaKPKXTFeAnXQ7qvgCy
5f3HBKZMgst0WCVot+1eNs4XdVqpDOgFIbSFjhb4/klnlv5Dd2UpDO/JhXMjlgBBUsuVlpqTAYNY
ONw/7UisXAnuWBtDqY4qhSeRJXRVUzQIciS+4ZnVm0f2s9bu2zZc0DU33cFTD7j3j6z1R9X0FX45
P+ZWhbccPvNFwQXhUeBfJg1Z9JNySif348/raeytgi1tMIZn3St86ib4oX1C7grEKS7QjdsJcrub
l4Z9Jp9oHu9yjOzjddPOOzaygELDX7XA7dngAm6D23yUL7U7WzkfCh0rJsxaRb3a+0dMyQqFdMN3
kxLE2fstI/S2y7b3R98ix+qYxw1gzR6W7c/qZLFPS1WtkjFMork9zdL041UouDm95+dBG+4ocQMb
AwAB6ZH1A4v/9ODDl7JAuQkHOHuT5VCM0b3s+9C0+zDWmeZ9HY71W425xpHio2BU2xvJi130viqR
EvRs1GFnR4MvYqu0mLwskzaRgeTdZqE8k0iaTObjBKkpGL3XNw1LcnyMn5A/yYd1neMp0JkCYyqf
yvcSvHk+li0xkTPpG/ESnkbChgZysRfW5NAXo71NT87KESe/FZHH6FFBlvR9v2luP2yt22tSVQat
ay2VswJa/VqvDyCLK5oIkuKA992w8godhWm5n6k6Ow6UmosOkikWamKRxjaBeN8i14cfanmWP4R3
dF021codMkBZZCAz7/cM2kA2qfAPpCk6VdumCSXsM3IEhQnfMzk34NGeurCmB1JULw/8vssdmFqW
FFXWO0yEjdeBx3W5v/ISBzrQ8Im/f3VnGZR7bNimPUnphqAhg6ii08rcZGJ8Wj3ffbUe9B22Ib+A
8T6YNBcYKT5U0kl+q2YQcTfp2y1gYzl5p1WbO+HJlV/LM/TJZgn11LXwMrglPC3bC6ZyJATq1Y2H
zG/M4bA+UxsKG7lkX/0WHKaL8MxQulQH0Xod0ka55SdrBhRN7ZaZQICo8TEUEQb4D1mTg/+PhpHs
UiBs0ZlB6rp32LeG3pR0hlci4lSYVE8YYXr0kwfQ5G/wvRpbMey4juEVvXqkxk4GYSBdi3E01Dn0
B481vMSxxXN64ktmZfjm1qo+WxeSHXBClADZ6Nkj+VJWMUzk9NRuytjJ0Yw3kCX5E5cewhvYAnUq
qnYzu3qLIzKVSuDqXyNNHubJmHSSvklB0cD/IS06uBBAwbuA1RQsSfURIcDHT1u/h1kFlp4mhO41
9QtK11WGzfDJAKAM5RgSIJZu5xyfCJ1dtjQy/gytMDM6GJs5BCd2ha1jOwUXWHBJOJyRLbnjGuLi
zx5rYTk7O8OsNjHoPE0XqJNxQXKZqlWksbTbpPr1y+j7JFQaoXrpCCuGZYwFk6terhANY+Jc48BN
2UzDrUX19dMb6Fr4ulwfxpOUAsM7hti7HwJDLdKBlQeL9R2T4vx7qHT0eI2l9QwpZlw49Ovlu2nP
G2BOY04QZSvkFE4g+5bHDLWztaYKWXX7JSdo7mv9wLwCgcHEMX/DxRV8Ux/3kQOVenBGVQl0cxP6
nC0EOSj96rY6gIyqSxyxT53iiYb3ddLdTpn8qMQ2/HY32g9Uli6jbBz/CBfa6NAV2J+vyKERAeX8
YP7mW2YWqh6SYAWz383aE/i8vg49uMYa/C6Jo7lfOi3lOgdbxauigg22hpjg02jWzcNCq4SDQaHT
B8leaW8WtFW1OCW+QsfhQa292rRAnE95Gf5vlvehWzJ/Cz33HTA4JO0z6i3WyE00ABdcHgybQKk0
e8VgnLuahA+csclLU9/PwDrf2E0DIDSOYlAiFqWixhmERM+SoDUFJc4U1BSvJArPw/8Y8zca1BWU
YF2BwajS8hAmgIbhAVpqweJRLGiPMcmNKcU/L54ogRYYc1KPQA8HViWeM3nyFfYWs2RkptfhfZNx
1jKWWlEUneY6TGu5TCQl0oThAyMS1uncu69eiaG5bcoaJMzrMAGoVjSvyxrDb5lkmdz62st0ktP0
77r7IyoXUrkk8SVhkVYbxKeuJCFB3NzKJu7kL+LgRakMYgyK9gnX8WLg4NMIQ/T13oOgW6yyxePJ
cUeVJC8hMgqY6oC4LvdzkR0OOFQNq49qsRy7p3NBQUlWbhtIPg5E7q43zkk1Ofx/K0VIKM2aZ5VY
RJhtPr5MTulBibnWxjlbVv1KD5CcI6Vnqmq5bYC3oqp4BcxDzLF331CmcszKMoM2vGVk+f2l4Q0z
N2EaSVsp8hr1G7rqPtOJVoJfvcT0pAAJ2tkoGP5+m/Yj1aJGFOqA9XO1CRVtfFAGPTNwvlhjEGKn
R5NZd2IRmg7+tYbqhXuC87SJnal4t6bZOEiFwVsaL2KhZ+MfHnDe80zJZPbNgH3G++OPN5ZYFnNt
tl7oZTLU7fx7owIS07qx1ZaAW6whqxhGHKEyqejY/TMtQ7lpMmEEQ0v1jr/wCD8yuP2SjtAtqu8U
8/+yPbDa2iF3T+QB36odHUm7k+fd07gPZNbqnFifKdnk0n9YybceJosyjTcWtuQr6Uae0YCoZaWK
23Dlcv6CG4UDN7/EqM92jMuPfzrEffzsn9Jz7sm/fTb7OAoc3B/CzEyFVEPVaFWyP/wG6lrzelhc
p+vTSoMWbHrDzHjSSEyEaQgNL0mzZ/cT9scaACet4DYtqcJPD7v1no8b0KnkcoKzPNRT2sZvj2xl
hHsdifq5DJ01Vc4cQ1yGXs8wkQxQCbIU8Khin5enggE7+amfURYdQXf7efpAkN7qwYt51NI156WF
PgLkkNOGvMgfauoPI8MvVT7wjD8iCK0FAqIR9m+92wCSM2HuOfOWMbzhmCgge5oYmyYZoLh9xOK+
X0nfw++4JZrZgrg1l/8ArSSCJvzRYIV5f4fqSZX3AKVSvMNd385E2FbBaHXwgPSXxc27fkkuReQb
zVDktB6PCOun2MfKdhUP8K9CC7s8umk2ebmVLalnhM+fdoHNYfw05J+D+4ynI2Mz6CCqBlS8QH0x
y3OYyJ0f9y+NTjpcHTl4+MmP4kwZ8Wzu+qZebMqjck0dP1vNqDZ2uSGID6PxRdr84zHzRXDg/+lL
OjniYbTmhJJBvofNXyHDvYOvjuilORazK89UzsbD0C2XGMx912adrLUPqfmo8gMOUnF/E6bHTIL2
CCLn63Xg99A8CPNcYIRUzHoap87Qix4Ag/FFR1luLrJU9WrTYQFl96z34FWgsgnlChHBK5sDgX6Y
JUKjLi7iBpU7hTo9sEgGRpyKDYi45ksipQecMMClAWkbGtW1h4Kj+bGMWhdx2NX8wjzPIiVafgRC
IHdMavcfhQhDuMFBOzQmvm6X1wjpTx/dkehHtOphrd9eeNYhUq7kcEPdJQKPslZxXTv9kbDCA6ZB
4gYGKOqx+WR0H7/NKPB12fGK7bMJJIl5gV8aSUhnl0wrAlaNc/Qdd/3Xgf+ZXDYqrepVKdfMAUfz
syhkRtIBPC6xcfAFnFz1jUuvmrJ+1Q6iQDFp91H9Y19B6qvwdNHnbZdT84pcl+xb4JsdnsesY/dw
3jcMNZcXUuP94d0evzWDh9JmdIDlnpRiF0Ck6J+fMCGmi/cL+pnDbSMDckSTa6ASEvVbyPssosJy
vrBYQcFIPu6LpCpZR0YxG17jMC3GY1ZeBtjBmTIdoSKTAYyhq+TmjJi5jOJsMymUyTU6LNv0f2lB
YAR/wf5M/4dTNkNSRuQVRy1x7aaH5RbSS+kxtJB0h5KLRXzYkZIQ8nFbAG5KHe5KnO7Y2kWppGh8
raUG+GOgdxPB2iiN3RUXoeCo32SiQ4mazjgRFrsYRTfRWCRTWfiNk8j23kzdPjIlzwtTGsKLpbVm
qkkuBXguQ6Qo6oFDcKNsrDHpP0Q8z4lCJvj/vDgR8onNh6IgQN3BNODnytcm4qp5Dc6oWE64yD82
VeMY94edvWLt8cBgL3b+/pNqf/XXAS4ILPdy2Xc99upHWA2DKDF+lNU0BiPoBoRjhXyakTTp/i/m
cSz08UQQ6rfrMfzW/ZiH2YFCnOnEYPIQoosKIc89SGWqXAgy5Kle0dKaeNg7tMmM4pUGFxRWtgr4
GaHAQaInoEhmCuWWgHy+xjFZa45jT1/wZ5qzZeQcfDqdI87tYH/XgLGH0GzqMe6OAMIX8E1z3+8z
nRXsU/QOXbOkQPSeWe1g038q3sQygYWNdL2wwe5qTS7eOC5axD2t2bzQFXJVYDV56JSOtIbqqN5z
M1fG/RZC/Gp1yrLwocJqzQSIGBmLGLh0Z6OkkgtcoyQ7XumL2OXsmN6k+UuvoVSJKSZnB2kEBGcg
PP3weKMZ6MTS16qShWbdnp1oKCW4cq9nxsl/902VGmhQpUAHZ+mGMbVI6tcrwy0o+gDx6C8bhi0j
cb407LJDIMLz+Jm7O4jMmVTyNrvcs9aSTsUOzlUPMcMlzpE0uwAWEoLDQheANMobfO27Qr79daXz
OJLVQm1e9EZUvDzNg7w8UAfbKRE2MlQXDsU1kyp5oKuYrqqEtecfASjaMXxkyBKXE3DXONYgz+Lt
UDuPyJ9s/T5pZrsBCVB8xArK/dmkreuDpQT+fG/3WwQcCTlyGhP7LFHvXzV1qTeyQJYKRFJX8z3q
0+fCs8mnRLHZposiOxoV23jcyMN2r3LGS16h5b0+aaGK9yIyX2KBBd8oDL3iVhEBZ3Z/c9bvvvTj
j67vpzJbxqJHNLDmOVdmZH0V2oNjCwJZIE1w4v/6lGI7OEbx76RNn3R/QtgMq0R7TrIIHdQRHcwn
S5waXjHKzXCl3pjbu2WrPBBOGTL3AsVXWdTd9PKnrHlDew+YE+1tc1yRoSPbTYwDrNwTbbGMnNzs
XQwiwUd8VCxMknr0bG+uspeKaPTmbpNlZQYiVW2HncRfNqVEu/davtv1ndJgy+zuiBnODqWSbsPg
ZBc/SnDCqx7CnA13rP6tcCU+hJdHE0ipLICJGkO8PnwPO624WC2Orx4CPJbCdfd+6u9lK91IOvAk
5nh/N4GccZQvrX29h7ZIsplJSb9g0jLtQz1NFtrZCNiQzYL5uD3NPtsYeQvzlAfuKiCy0fff1Htd
gUmmaG+XcV8w0zGJuJOVp3OCSX8Z/DR1npJRWz7UJLJ3FvlV3mCpConTMn7qinGDp9ZyGzR6KLkP
7G8nShegmj1sSZFT6kbt2YWHhrVTqH9tiHW5BVBre1m1f05f8F3URjsEwc2nbQ8QePqDgRhR+0RP
HH3/Ei40UtlAf/IDaXe3dURmVcjKrudj6Uy4vKTj768c3zgxxOBF9her+TO0uMwBBSFJW0nRJ0Jn
cLHX5DLPSBEcop7pqrL42TJPoUC/RGno5rDT6L912DaVOJwAT2c+NHQwMjcnGgl0rw8vKpbU+OIX
j7lyXwDnd+Eq8T5CqStaqmQM0CCVt7sTZ04mC1YgmH98YAUTdsNnBQp3wNlYkI3qo+w0BA/pmL0T
WgWbKsDknZR7O0uXzBWNhluAScF2ObOPWyi4vWcOMQ6OGbNEx4m9MnobGrK+tuEGcmoQqDYnbTFP
UFK/BwKslGrbG3ly8C6szWtxbcXQ9l/xcM9W4kG6LO0JwwgrueHzLpTctmD2X1rTIHnJYaleHmnM
axxb91RxF+1LgT/faK9rqDwGlYLJmChwB4AlLAaH2l8F3JmBV7OdCGpFrCjY6uhDdqbtEGkzW8qL
pAjIQFNBclsYV3ktjNNa0zKT8lflbSnr5y4/3HmdCqd2cN81Ridvgagiw1Waj0YpuQ3RpwEsAE6t
6r5PdD97zJYepJ49+YBMgDYqyOqg2eza6o8bBrmoaXLPlpSGuTVK1vrC/dmO5q7jrKnI0tw7aApV
eK4HtskmaWZhayGAxNrg0je8IUhFd3NldiRL5VajDds0V/XkM8njSFFZ+lbbtzEoG177et6Kxlzk
yuPYSLX0bgeYSFLEhkQJNhso1W9O+08imUTRQfm2ahgIQsvo7HgdjbMax3/jWzvoPPRoF25peO1j
icVZoreScRsLylz4tqMCK+Mx76IwNtM4nkGC57mExO1JRNgmYYrtR40oVw/eItgPtqIVDPolkLxr
iX5DrsJtc+y4jOO152PI62MKVm2XLgpXhOQy24u/5ZBO5ve4kbmrZxUiwAcCm7Fs0EDyi8ZlFwzW
Mbh/roemYWtOK13wYop9fVunhlxy3TtPz2C5cjY0KAVMnsGRE0Q6lkZ9EkQkcM3NcH38G19bm+UP
G5TFc/AODU5RupX2+lI3pKdYvTTYdxabVVkqaMsbZ1+7qJEu3037K371MlaXlSU3ES3ni+ORe9eS
Jqvw0c6+svSUtpk/uBxTJTaSvoCXyHWmftqzgczjYuRWCxZYXGM9wx61EjqBiHUxlj4cwuOJOhNB
DVHLPFvQ+d/RUHmj9XNLBeHhihJAwrz4fw7ecKz7U/ios+Jv916Avg5Wc1tpTjWaX5f91hS0mevi
SfhdkF6MoV7YPH1S0V2+fnZ1zNvjg1DWw0kC1ECFSeXw1oYI+iQP8frxRoVJ+g6Pl4ZrDGfNRcyP
Fzt7R94lX6uT05ow4Hjp89tcVxWunUrWrPA5RxODLtus3icOzu4n5boAZ8h61RIjgSIxzKNkcOv/
zgepFct8IhNKiDHjg2b6n2N+7QZB2QEWnBs3fd5E12O4C/za8R/S1ncmpO6f3U7owsYd74Je7/dC
y48AtOQhA5RAHto1HKr3P1EwZ67LFXV6U8RC2c/8AzeQWWkyIgHCIfPaP0aPwBcXd5ZWgwAmx86i
yc6dWFNJu2YpVEnb5slQILRuyjZXm20heg+hmDxGbYGOGy8C+A5GVlIb7hphh4/y6l7rNynrnAHy
3WmMRI6Mchuth0KSsVFM8iijhnuUoIJKJCqfBIyak7c4xCW32mzD8Y/yomqXDgMzDgGDLAykOQNc
LMp0RZARNt2+vfZKzf9EDBOc+55bc09oRKj1LNhXaMUj8EisDj4WcikON04nUFyCXpDOV+QamymP
BmBUFtfhnOFqp2WqOXQ3Xpwu1sGVC23mkB8GXNctyPfwZQi/ASOvMZSv+wneWkR9S1rW9Zxt7Q+R
3unUegiRY0I4OoOld8vD+SJL7DVqaWK2POkjL49Ho8zVBxF6gxNLwekPRr7oDjbbjfrwOwSdtMwj
IpsrowSKLjZWeu6vkrgwMB2c28a9vtlmxFf1QwY0zOa4AdQR1n9YKT3il1FO7gouii2SyeeWwUxE
VlHF4xzuTSCV3gKOvNstALzo/LBqQAQ0L2Jb4ehVlPoFIy3ry89DJxUcF06wWOIviZOnvOx3yTQ5
w5XxNCcFxmKcyZflv8u+s1+gJ1GgqFzHx9KoJBxA0OcMknASfXeIixQzYEYDorfqowZ2abJ/KJEG
4hcEm5DEUJX7TtImOgpkqYSRwmJyUY4ZuNCpFVqEjpZ7EsFpp1/OIzypN27VKTR1LnlMEmppyfMN
sP+xBCIfFtb0L0XxLtTTc4MSKgEFadqZ7TCVb3F2ia8FfI+bbl6OWvbGLSczqacM1BpzFTwtbAwV
qngTvoVL5xcYuXeo6xDxT2Tls7Jl4zEN3Tat5+Jxr70t8tGTiIGym7LYS21rZsLZWQrcO5+wSVU2
cxWuZV7TPhUtPLbzIkcDRQ9JsWPjnTJ/+gl2sNJBahK5K1vRJMhuECXVJKyu6RjOgjw6VfCb1aQ0
67BcioTIHF1DruuAms6bGvXE/gPbrLzieM7rJrRJc3XVuqA1wO1so+kqTwVIS6HuY86Pqo5FDL6T
t4k+EnoLC6LvJja17gFtVheVOux4xi/Dk0b4icErOh/PxuFNPfX+fb1WdKWPDCxVXGjlJrSlOGhz
ke+h0oPsXmXU+Q3TqEFtfLKCwOdFlVJ7yp6tHTlDePdz0y0Deg+tZ9ieW2+tknGoMOC4Hlv7nllK
yF46xxcCtSU3DRC6WaNpK/ckXy0Z58QDlqFMM+dhWLuyyYWzDw2COwuRwtEQ8CWCAQJGG5mGiQuf
otTdZHtNsFVPJj6VoU+7dEE8ptYlRQ0oPrnEV8C6JVfQl1x4qpeDb7E2bRPqv/owaAeUIAPHEF+Z
j1XXe2HN/dwuT1ui+DQDO/Vksa0nguOe1jjEOyW50fsowE3dNqacbUcfHD7pDWRvKqghFCaT37c+
0XTlLN1N5W3T4o6+GDMYPxurxiLulzaZqwcwsbnYKcvX5Gs52Pc6grm3TkS0qXNOYhs6pdq2T0Va
yTWWOl6U4kApX0CJ7BTt7XRqkpDMJD6vSKg7yBkZ5jjGC0yRsFijheso/fSqiSPeZPBAkBERIhzz
vny3G+bw4AQDV0lVIkPiMiqc2hw/OujSLFtZmGt6uRDWGcC4GDQe2QerRMRXO7sgG8xpLAVw3U4a
S8CGiavOOfC7jpHjY5Vs6kBD82yxAEnaWO9GicYqYFTcRE56OwEizBtsYYhU6ToK37EObqpzKgx7
UHfHA512yAIUic89IwAT/q07pdTs8Hk6sk6+DbjBbh8/i8GUmWLluSKgyDT4Kv1IZ4Rath6DxWa2
QTOFE7Iyhh3RWmEH2Ja1WZpMGI+e1QVZUlapPNzjKIvIxTgDcRWUdr0LXOPFWA4hPdaazD51i/4T
be8iu4iOtx6GNbzulVs+UmlveXMI0xjcUUl+Wt+nI2g2dzuzrBrkJ/tGzAk28WUHCkmuoFQxip3U
mY4TabumXIzb66r1pBCD2fvsN+GKZE2VmFn3nPvOI1amoLaR16y1P85e4+3+B6vZgBCuue6AP89d
MWs5o0c9w8x2YfuYBK0lNeB3KkkH/O7E4SaspPO4mgkdyK/aTdVdHFxNKtIXY1axJTPIxiBxZ+N0
INETA22vqKowzz7+n2Ej7sgw2tyMWjKCqJklpQbygncEbzROjxWMuHrr1TQScG4xQ3AiTX+YoWf6
zphqCzU/RECHOAnb0tytGn8Ya/ArK7WuVoNA4v8Yu0u5mpfr/9eQAsUjQlpRiyJmgctVS8idRWQy
VZsIzPEXXsFCAv/Pxim8OtI58XhX0YyQntKikmk2dW60PZv7Cb2MMmD+U0/+LwZWoWZ5gEgyUKKy
7CM66HvKiY8iA2JhVcpNr1YdCJSSbh89ABtKtWoWilzQHYH/V+jKFN2N1VVx3I2o4kg3E+KrDqVB
0ZqBfuISitYkmEcOyhvDxIpjIPZj+TmN4o24btZJHnk8TKxEmQDuCtLTj9FmiNz9kbxcM6/4IR/X
B/A6MFVJcFdqk2AqCz7McsGvEqHOMSQfUQFyLorYtX/TvU46QUnuY3/jpKid61PH2/I/xK2DX+fJ
MYu/u1gP05DOf+N+W5Tti4sLVG/b4uFUnkL+/p2YSsS1mz9s5RaAlTrTX3UKdC2U/u6L4sgGCDQ7
PBegoDxETDVbEWk4ASHbn581w0jsI3YApyJr3XdiDpkjEicFYI9upP9JaTs/73JXuoBmii/vDLdy
5zbtwLZPqTZxJ1+o1bNJRho9FzFeaKMjR5MIqll6GET4FR6WKkAqfwdBUb4+AJsfmSxC6+DuPKKY
K75VJSmvlZncOBHE/NBFQrsFBuMitn9Up8n60dpeqe0BY+ToTQqRukdBpG1LWswM9ce7w2Cema+5
YH7S/0VgvMjneRq2ZtTHqoq7iTzpOQxxw7OhbLgbIR7ETbkZHAnG+cj7xsbjckr2X0HariHSwOgQ
kai1rrsm2fVpF76ex3iib9CqQ2ROEhvCWy7dEDlFrex/RdkD6BKCTF6x9qZfntYuR+lt9XIkCVnK
48o+R/1Zxma2N75Bl21h4LUxOVHc+FfXGD5OuFMmhHfJothjOIcHv3rrQexyBtS4+QlIGiqY5LZT
wsTZNAH/N137vOmDnGtuD/4xxlwZmo4UUpa5WYRy6+w7qFzIiIxxlNJKx+7f9bUcMzbT67YZcC/h
xDnfuRomx3HjqrizZ2q/3tleGzu9fxXFUK82O5msxx8vRNOz5xYq1VSuG74pea4hJMxd/umQix+s
SwKlwEMoJ/GIhLnBKQmQg+Gf6P0LJ4R1EW53rvzAqbAHBI7xKZFIwL9hW1zsgNWpzt0AsOm0jPTk
3APFYTknykBvXM4IGu+gxP3G+29CzB2SJ8UsNW3pfjqdiqD11lCGR8rCtqAPdHrYMiK1Fo6XwyA6
hTDJ6Drx9yFFQ+F5/atw5BafrkFT9GNI7Ax7PoTnIFNT87orxkKfzfEzRT0wTtKW9gD5q+K1/yT3
MRz6f3J0+V8+l62wTSBNEEugyxTh92Mtt7lmwV24yzG4DwNRff4MDbd6kC6FWfcbXevuImPZYWaO
1F2wWzZ5inIjhygpfZXlOGJMKmcNPcFufB9eHojNjWlSWcXnNyt/cv5qT/D+oU/sdQf7/EVr78qY
VnWjWLWDGf24rRg69f3K78rIGOb8NuFD9KHzpQMmDGxX2ZeT8FZXF39ogdQQ+6nF79AEhw9XI73q
MO2lu1dpiMexNYENzXi9uRqOiiaiGguhFbHlDkVqh847IUt0YwyzSXDd+NzUih7kPcfnx8B3U/+C
AJlSUWI4588QpFQ5Chbc2lmapJiJTvnXGlBfOXomrS0/wr7+U82Ad2fbsZXiXC3bqh8WV1m5FMmH
KrwDZunCl4UIfu5Y4yOX0MPfFTNoL5YEWTTXNHaXtm2J5wYqQRB46dOGFARFSStdzk1R3knP5Qvc
s+fdcQZ/V/xrNTwcz02QIo1eSKiTcz7f6VqJrjBYtMoNQYlc+uy5c2Ax8mygNYtyNJsYvsifDSYw
Yi9jJtbZ2yeZZ63Dr6jZWV0TC6l1SvF+gOYMolcffsVBrVVJJ5ea7rZPQxS1KOGuB49QImAvJEXq
MiMllWMJPkCjVzVpitcFwUkNJKKc8GJDdsH0REXZOCSdnphtxk7gFf5PuL5aloG2B06ed82UWeJJ
/quLtQsD2+PMh3qAgueYDRJKIIm4ruJGhrrdE9axi+pdunk9Iu8l2D1RIpQiJAA3C2VAtJojwed9
fhlhAKk7zZGzIewv1aCUbEjkTHLVOD6cKEZQw9KExtjnRPhz7IrZBoeWfsU5yU0BadEnxh0TBfzy
MWvjNBV2/hz2eQHXrm4Ek3JF0MExG0dK7ivGbyr9a5cZyHE3tYf1DFrAeCy+69BRl1muehDnEeo1
uEilhhLxVP9F/cy5DVZyvUdQAldzA+9gV3veuQ9edfvVgedGap/rIpxWEfHQJGFzRGmTuel+zVfC
mfi0C/2XsiclCmCAJKFMwti5k32X2HjOo8EWxr8fAP0+qWBzCaERRMrsMcPE5X+NXzcyfNdvC+s4
PsZZKBz3nUdQ/kVh6NSDudTfeha2wPtvMN3V9qiNykaSAvOL9nVg9/kj+P+A3oaDy7e6KxQGkmJm
OZ9US3vVPiRIL97TjAN82gmcEqU/lJ3eTFWsbFtJUke/sd5caLFZofKitfVBmpiFEbybbQjO34Kt
5y/Pi/+k1W4BZox6+sSE98Esi3LkauytUJpo0Oowda5NbtEO9HCsgElbOF8QFyrI3jLPKQabtWTf
l1nJO0A0T/atsZ4zUm+eF2p6rUFf0mx52VR4D3eCkyUlm5ug9REbxins7AAdzjPZXnbylIvUETvw
nUUgX/4jzYacWzS6ICzvlnSQtkuWuSBorLtNmARD8eCeOauv0yIRlsufD1RLZvAvHWZPXVDB6bDS
sQspcR0jLvoFgEPbV2oamOmAHzlnW62yrN59MfI5oTdU+sji9HD9IqPSVff/9A7RT7/5i4Dqoa++
cR98EDsqgcffesbd/R6yfU/I50w55PX21fqQg0YgnLyUkUhqEjByPEmJfG5mLcDI8bqpoJjYf19P
dIFANd4guEzUvqUnSDjX4wlCI/ygwN3wq9S79J9sA33P3tkRnvKpJ1Ts7hW8n0Ar6IAQTr3Xw5no
Sy0AeXGo6Vxt1RQopl8jniZKJqL6ORMwmAh7tjUjeoynl84YZL4RG3jzwyVQsGuK9u9bCt/5mOMw
CBSaZlo/PWigUCLInygl7Zev9+8XqiaD1IKRH53pq1UmACraLQiHeZKG+hIJ5TqZdnVivtxWyTGo
3KHSFmVqOzZUzD2NV4BqDYCTXCyxIdcnKLpOmt/OwYrwuTxB0o8JlhOuhjqsOjq16yA8f+Uj9112
77KX1K91AvIFRK9rkSG6ATGJ/P+pnJ/nBzK8bLjz8vv2qQ/qOyRr4AOtcBzFlyPHN2Z3KGUj3Ucv
VRhcUQu1UWNzUqyXkTrg8YEN6/mQfB2Pv8kLLtqwM8lPiPZ+igQAgAZGGSplp/S6cCBlcWXInDqb
lRKxmpBvgvAQeOgQVGHzkkoARPNse4zxBC2iVGVL/sVtj+1m4eV8oQwT2aOYEbwb9/IJCC7zAi/Y
GmjtdO8Tn8mW1yrdud4IiqmyjM7FBZiSJYd4AGpstvry3N3HF7IMJk01BhMrFWL0ZZ8WMojeC0te
pvi+71w5C7mq5Iov0fXRKKAcZnSN6tVM25W/MYisV2W+0M0IvWAIqGzdlTBYbdu5DqWvmmB09PXQ
ESNUbkXIQ30ocVXrh/juHljPh5nG5ET9G13HClCWlMaewoDXeWvEdQtvzXddm5Gf/+LgY0OSkB4o
49y4mVS8y9g1RdTvi4sfLlS2OLiDgqooZiPSZaDVM63vOcWXPhtGCB8uTcIcJJzPLBGXO5/gr3sa
T8VnS6Zmh4EQuzOPYUn3ZzoyDZ6Dxm4BHiNBbZxHaIE6QPUM6/dUmac1gAjwrtkrJtfRL7DwqAV4
8IJRoQ5bMv+5cwuxPsXksjKphCHMwjE5+1hUf06o0PmlFT+sJyyFG/jSMLe8XSTcXZKf5RMc7v7X
dZBefgOCCwEDsrMGkkvex1/wFGjiWUOLXJJObbDrk0F5+H6OjclC8b3AhgK4aNLfzs4PAVlsNp1V
ziUMsqGA8HEIk/boPXc3SX2pFTmsBtECMefY1Z5q3eui4GgD5tyR7qcN2QgMdLfkEG4GY4UZcViA
rDQnfYDc3ZDK3bc3pKfht1lcyDYeCUw60+swqaPHjbeiIxlek0Ob0C+8VOSr3oKPykcDx148MdXa
NcqWppOwXli0YnadIVtu85zI0zuLP0zpguPMN5I3rsDRrA0o1MIMUv1Kdac+ctnXHkxUGu7lL5sb
SLfO+t/GeKcCZgAy2uXY9jdaoBoHygpmA8n0PhB69/rqtZQxU7fBqF9R++VHPA/DVSKirN2+TDpY
+cEkCmLQ3Uv/Zj8lHD0wTqWQ0kp/6WJDkhPYch9HC21v6QIeBBdRURlSdmUyXGYwQ3p36iBVaOHM
26ICFNQcv1w6CVqpVL49vAvucgl/7q3E0uiyNqyKfBWugi0vNYnSzsBQ0S/TQx0BiqgdFkIMaPg6
vKLALzrTgGzX50goik7v/+peZDhmVepMxohktWKwPEbyBpa22RahWkwULi7NOtdZG/Q6JnKDp5DE
Vx+/QEKXg0dJBLw47QWoCMz95EaCK6UZdmPLm/ZLxYD1umWG/fp1j9x5/efl0JeZD2MT9Fdn50EL
OlC46MLm19WlfBPAgCrSN9FZDyArbFG29AdVCA7wpMt5F3a7sVdsELsRGJDjnQnqXA4LUHeysRGz
vSa0pSd25yCWGhMRsOV418gxTAn9sN99gz+8LFIPTFojNpnvvOOig/lRvGw2QCUhaFZoyxPXiDLf
WjE85e2KIomXQWeqslRIc4Dqk6u73cLCaajyLXTvmHIfm8Kt/gnpy8rXQdGDipQXFFSPahg2Wv2U
MMQEBrxTwBF+zvNUmtmCUpIadiBRkhX/4cmyXPng0QoP9eeVPLe5NEv83teHTJjY/4e/hgZNhwYY
IyR1WBxy7DlWhrPFlvV5r1ihhtAPTF/0lHXpH/OjvT/wCy0Z1eBTgKo/P0yXe46S/++uttNJM/NB
iJkxbxKejOSvIXDCW+GA8z8VlMDqTANKL6dY3QV98oDgT10qXSnlK7GCVvwOcVu9xwfpeIaInB7i
qzgglbtDeRYiVMK2PbQZeMvZim3rMco4GYC5piKYZzPFRt0mEE+umc2vO8WE2XwOJ8GKYvl4Ia7a
wHLIlcat01QWEarsLRJ368omTnxmrP5LrBmB2ROD/hZzInKFl/qN8Z3FV8xtykK4l+vKmYnfWGEj
jG0t5pvLGbbswATEjJjkApegBLtXxcnyroOmmVGGZDgmj/T3FDfsp2MoHNRH9Hb1NabzId78mHWZ
nc2YBqG1KpQCeoafu7WoQJZeZ96Vro3B7ooE5zdIP5Krfs9mpS7uxG3LbpN5YmSuKJOW1N+W/DUK
5tWhSWtE11hEjvchdxzQGuuIJ0U0YUNWPW3uRfydgNJpGg540/Fl96Ty0Bz5Zlzh6pqS+e6yJPDH
JnjboB7gB3Rj41Ve4lJJIOemkkNhZjOc+uDBMFHc0Iq/a2+ANu3whWQDWHVk5Tm4Auw/x3WgnOVY
KyU0O1hSuk1htgVe3Owag/FCVY0zy9Bh5hIsOL75ydYV95yo71mtycki37VYjkiTf+gIGNetqGyO
tLimot/jcXCiwcO5u5l4DxG8pIZ1Nei9DI2/PxpxRHU/N/HcXsXDMySx8f/RaiSJsLuJ74Q+7k5I
+r3hDnST1Ik2ZzyplZjBmhot/29VhkZUgO5GVkn7p2Nk0GJA+CVG2f8xJmaNvS2/iwhxLPLyJ0Ve
oCGdFATPggobsevsALchuHLN1f+MPiysIpZd0EkvZa8b/ltvI7sDjXx3CXWlPd90Ldhc1Ms1kpi8
dcAJjrqytV8YO61kXnGpOkObYG0HUF1NhumBg9SFXQLyr1o5sIZnq8sH4lTOwVuDgpwdHiKZYPgS
524AliLuRpIJ4c4MbSiRJkqR5pm/Ka6O2WaHpZ75DzERNCbQMjdMBabVHgohZywxSrRWkFiDfw9Q
wctG9lMm1BdScd6cNM73XIcGHn1LJLudqJK4kcIz4lod2E4z+Qd2Ln3o7HwAYWXnj01U9lx6At9g
kPcQkeC4bBmvsEt8JEnekOZGT/eyP2e6xSsPDzzAwrmTweCdN6N+UVTyTFp3Ey75Ct+56hCqUmn8
hodQKyx99GqmXAhTN0n5Prqavb0SO5VBMTYBJHNN6OqSWLVhy3/GOo03tFGJi0mdGW6B0EXscgPc
fSaTQBFIUd3BJpt4pyTgSdg8UPrXA5Oh+PdgfMYS8tqoZfHTRzI8xCJs2tCvhAVagavJbk5S82um
Uq4ntZ4CBZwrxxOMl8njI/BinYh1Egla+en+sR9QQFUCiwnSQxTznQVad7xcXictNcHKdsB3Acrb
u7syZqRQbSAefxHy+MJInW2YEOc9AtC9a53N9ZAIzHraosmf16mxu+pIbiZWde26PP8vz0C8GXHs
/17SsVfksUK/PcWR6n02AbAQG2RUd/o4yHJkEkL1kbQIg/XGQTjcK+bxWZwrLJUkjBXJpao5QRmE
ECy63RcBeOOHfuc+JzM3jKjytxJ+BCNPjSsVwYwVLpEICases3qsmkaI52trnax9+Vc3BpYmkIf4
9c343+YaBIf9RBCE3ipB6uUMZptOuo1LoywXdpTKA14T2SKLzHKu1lTc3v1I9Dr1nTAARirr1fnm
ktLEUtM+Qsn/+A46aY9EI13OXRY4LkUeE3pQ15HaWm5K5MSBfUwCueBLpOJrQHdhZllFailyp+sd
5sVl+yooYfg83CEdJ3oVvRMlTHNa7QrMxQAljOYaivq6lrepqBazPQxg4CnxhivgD0orcyquUEpl
xmYe73gskNeyqlMG/JvZw6uDKOvQL/aGKeI9EK/ShXZOMCCAhRTm41fYykTS5GnyMhh4nPj0hBeZ
i4JuQOARNMl5K0dxQ3S9NaUe3OcEJm6MRNS3XwLSmRNyxHkxaWcJFjtQpZAfED0d6wFk+7/FVY+u
UA8PAvQELmbN0UY13StQDxkLuyAVWmdpAxQqYT7yN37jMoLeQwZewGw/M1oJ9kcFmQjwjcN4ZDrB
p37sKplDX66wfiMqlX6Ak4knXTh4xQmx08nbNzk+9i66z749TlJB97m29wAmar7wA2f6fAnMvZn3
3bJJnzug0ykKB/6N1KCXWTu/gKRd1WNqiY2VeKPKNY3LfI3GFJCxhfDVvFX0dur+i1eCA4YPbaBb
4sWpe/TOzXqjSBAsKAtxLe4DkfNlrVP+9Se4xc7pVgzwFopJkwBpjsUludjzfnszUlu5N/Idm4Uw
RYpwf2N5KK+/FBqgn54ttlPnObuWjvv8SpXGyBjf1olijuewniNFzvlrZCEkYv90dqdRnGFufyPo
RMJVln+sdh9wzdXUN2/BVt8Dx1GNfebImhMb4M9m1LNXciABwlCxF9IO1x4c723k2BbLurAQSgeU
Yd8BIoetKtaPSRN9CcDtBomctv4/r36gX6lUs4Ani27OeLbUzhz9yGB5GDR4EAIyz2ecNiitF6EQ
ckCBFnmBwt8mjRnJ7qL8iWKY4L8jnUEIZUJSiZsTBVCafQTNTOpt4+0jUIGRbk6CvS07hHjxGeX+
phLRmaYKgJv6v8Ju4NGWye++I+zHzCO65K5QkP/pmbB2G9lMmujtIQ95sIFSjl2KJf2T3wOIdHVT
W+HZ7+bxDH9tz8q7nEF25NA9vdvdFDMGXjOJfAnXkder9oADSEQrJbA3PQPruSE6yO73zKGUPLZT
UMf0OmTpaRwWrMG07/SIru1fPX7DD68sIbjU5xAkazmkQwYBI+GWFL1I/9HxbScwrOsri7O3i9Zl
CA/e3NQM8zRXr1H5GjEpG6w0NCgDR9eDQ3xJa8cl1+7xDIk+xn4bkUf9Y4Aa93j6hGLBWyXRnk1+
3hW0+LZvYwyjYA8461X0/INKdM2XGCZSMdBF4JWMdTsIda0DsKYhx5avs3Cd4tkOmtXDdp+vJ6UB
bn7EqpTSBEFbtkL7oWX4U5mlN4GUqbIHnXVIKRt6T7pSiespBqxWCi+hCl4RHRHPJPrHYhAcYaR4
Ldhm9QJfhuIPtLfwwJ638FkDZHc6x9PpHVO4oUMWzI+N7DC8xjRAiWgarTe96YAir2o+Qe//mkhC
iwx1VE5mtOJWWwzn+iVyd+HTNV9P0TMVOlGII4PZpyN44tiQXp9WyjitZG57a3V+zFyu4rgpnQmi
xoLskKOuN5jysgV6gEbAoYbqmw6ifOvJ6nuKHkDsQCuR435FYNd4nCbjiIlFdMZr423lslxDeBbn
KwCq02Vs5Vl0+CgcfiOMho7Zbqnp7Xi0F0rZIeZJ3HCZ5p6uMPjwjf+vK3xEFzpCz6pvcGm/ARTT
hpANmnsfpMQvnUf8wrWD7lcl2bN+Btf4ziKzHej0x8Tvw/fTGRf/EKl5DayO1FW336EgsbSiIjHd
0HEwjyzfNaj9EsLbH6090+/WwQLvZhSfCEaDIqdwhZA+V+BYJ1t3Pn7PUO7jSr3qGA0lk6eH4G1d
Y3c4kX2v0eqYdCTcHK8yF0fx5J/8VRXxQK1Mc6N7oiuGxV84IxjrWA05/pMh8iHL2Ytqvl6JCGax
uR7z1QY3PnVuLh1bPTiugq6x8ZGxw92Xlcgc2hwUAw0aqoy2N0i2aYoJcZfvtaUIFoXu78+BjKSN
dWK2rvUROcFGkqZzR3H+8JBtAkjnJAn+ZDLmAlcE4VIeQ4n6pFOuVaLanG5akeYjZOl5TzOoDwiS
NJP9+uRfVv4nzipvKf7vfuuJk/14g52lizmPO+9D/Sd8AB9JZRaJRfkSy7MHOJf7pToEncHCEuKF
KAHa+ptvUfwstC+205MsnH1LU3bBgd13KCxLYRAoWUjm/Xof8TEAzyHN72CBK4SWSjRMseRjE6N9
0Ohzau0UZWvy+k3nVabcth00TwiQ1kM9IcWZKa1IabcQ7NbKF26tK3nDXzvDidXlN62ES3NJ4BAj
Oaes0ylBCFIMYo2YbtmvIF5okCR4rdagdPKZxs4ijxahcAIRiAbC0BhIZucVB+wpD22cWvyep6DA
maLOdnKrIwUtZ3ka5v7vu2m3TcBOg9a+F6mASqC40RNuPo4NTfI0EqjsW/y2c5Br9uCzAi5A71Ge
OFd2OYBvx7HJpYLsBWpZ8MZYcYFVAo9V3Ae0WT/eL9YgYNfbWIK8gbDHVa1AFuj+gwcj/t83uF2h
zptuOjweYUIr6vDFsAhEtgzg3mmVyHbx9IVe8cqh40KrI54D28HR26Q5aC7wjumcyVNgN17k8F73
8vNJk3Aem1b42Kq5df8nhcY2uUlhZGr1tzWVeV27DQrrXKAXO/oLnG9M3vq46j1vBK3LFJSOsgzE
IgcIUHwPoxprR09Oi3PEvxq6gydBYWKpl9UyPqYorixQ+E+z43ghOdunGrAlwYCtJXsg/sP0i6hK
ihU2JWv0/Vo5q4YnR4ASV7m57pRibfjpJ4LC2KbW/hDkrlaHpLRjn9K14z2DlEUIZrFYJptUfVrG
kXEoEz74W7qPDbYBTQQBSdGEsCStQW7Z6p0cNW66KfR3P1N4WPQraxKQsa8qNWVcCXirpoIL1r1c
Hz9f0DhGCqEeQzmQniJQyrzli9zXjDIqIKYfEw3qUmlL71lF6LL0g+LUUEJseBxiej1u9xk5E3cX
i026pRnh0hf8tjlZsYLmBOeDczDAKqhfzXvEF0GtawRGsZ6OcJrXJixHCa0f8D5WUwhhMqPm+MdY
qIVNr1aZ8QmRS+U6+W8LkQ3rsV8gQ521O2wTToGIz13aJPVPO8FUQMBFrcr8R+NJd1pBtUHreB++
pTKSB175DE/Nrd7DLitn3eX7P1FfIhDjpyu6zkp4eKD3ipjg27mloj+hYCAI2Ykj8/xVshMjl/HG
+Ms5znODmf8D44qvYfZ/oJ+Xm2Vymkhtc6pr4xNXSaJrOGv1wiPaWjZH7ttVj3Iz2QlDIEbhkDbt
q8LSdvspXlL5v7hO1hAW2ov32Uy6wJ18hp9xEeEepqQUltV0h8O5e9CsRl20R+j7TYk3eH39lfcI
aZLnGexZ+Rh8P9sNtZ3qZ44RzQiD5idXuuIIVx98CJiImp0tqgkZlZ2KW5dXM8Rbtfg3MciK5Khu
UmcimtCVeqEezmiyG+ehu0PASTdieH54zHcTbQEUNxo//x5U9yDQSn1AOICnGKNXUXCKaygshEwI
JqCSC88duPySNLXXoIpijYWL+SiWzzjmKX+pOFnJDdZQFUjc5PjSVTG3NdLeEeQBN4vtnQE0kJSX
uvItFZiCu97R8L2ukALp6Aqo7eULN/KXo/zgRjAerd4ERMw0MYYAoJRKclM4bU0Qjc0G1VvUaTAW
Hys3exZ+ulA4N/MouXP/VqQJJTzizFxYh69zgX+SuvnVAJ6kcHYmKqyj5PUSkdLO4mIIRVV83wGg
ge2er+xTBt/MnqO3GDXfVOr5m5RK0hxkYd6iALQdL18j3ab9yS5iC58UEmFdCOMEFCyNw0iHfTHh
0VGZGubslSkL9UUA6BEICgF/vYfvXhYfTYSh9s4bT+zBAuR92AIVwJbBMLQSZ+2BZaPV0qC9oeB8
CIQCQ3fJkrAYY6AgraSrqfAZ84nYfRUJwwOy3cDlS8D2EOH1fK/ptB2mt/xxDqsNky9NIOoE4+c/
RUK0k0ruMS6ihz+vJOuhpc92TiyDPlEQijAXBFJWZoXwZV8ah9LXDsSBRfcN0rgEjA2yEXXYaSOw
ZKMCQw5gFL0NLOnk5aCuh9Svm0ufiFvQEf10oLqNBXXPtMudpa2oKuaMeL627xioJy/J9qXWt0xX
EDF53cBBW3dTLwnicpnOJPTYrzx1xmM9/kvC3sbeRaHp9B9V/Zg+lrvy8p9kpirZCgweybKnwRYB
Exgm4lbHIUAm9EIMvosOJ1F9KFBBcYQQsvUDFaD94TbGpvRlX/oRhDAo/4gONPeXe5QpdMWWJLk/
k25DZcrcNw+YMEeKKTAiR5C1YST3byMmn/SR9h6XSYsqJrKBVXIGLUva7vbnqTt+cgXWPYISrhnH
CxfwW2Z5yg1BLnDVY70rpG24OADJ6UXLIQvLB9ZewZT6Dh4NRgTc74qA5WilgjGMJgHZLY2ndD4F
lfEXoBUYSMTAW7RLfsLhz1qFGmrHeJ2n0LNkn8nHt3ZAmxZRGs6cLGu6u5LGe3RTRrnY2CTKGoEP
opcuaU/X7ZWMqmC27nvOQYAV9IyDnczI7/UlqUVkAntZgeod+76C2Z0GY17nIuf2Jc8eiNv2tJBX
XQ1dxrKlfEPoASHTwe8IO+JXJercI5g6l1ffEQ8GFvmRN2FsJgNLkYfYIcthOKde6dD5HY/i65sl
WVRglgc44zTpUATB/XVaxULxC6NYDV3IevC/YKT9RfuiMwnljJSr37D4WSZLHO2WkXzIsPwB6AU6
27I+jE9J6zyc7UjwrTtu9wCququT/0ESSb9sryI0punDW1kzb0HIVnKxpw+OPUTx7bCWEf4ZcDC0
7vAod+Ah5v9vD7M6aE3oswHo/aORABbtZW2wh5hn6me04msy4zu2ulB9vhBsfQwpp6hJbSJ4aiwS
MXA1xem07diiOGmHFMgrVNPu5pH7kNY4yDHZGrR/7KVHPeMgsjUwIsQPka3i7o9M6XwMD+5F6Fp3
3EiPuJfMbuXOo7ICXTNbYASo5NK+DEHJ4WK5yqv0kYuMbS4nOWWOWjsHaVymCmZ/CAsCTu9eyttl
oaGUdIKgf+QVZnH5oUabee9T7LwUapqeBCB8FkYX5/cxeUJHlfupCFkUy1gWBmWOcmNT41BS8eqs
u0zYlQGWbG5NvR4DnJYWbE/wMwjWlIrb5Ax3wdEFgBs8JqONqSQhWMRJBdByVw6V5NIyUk4kssmw
2iIY6ogxn/jqgpmLNuCqXHJIq7vy7EkkREQ9XZVO6pSAhDbQ1sLjCHMxb3MlTMdTFZQ3x64/LcNd
0JpnTHL+8b1x6NtpPQ819vjL1QtsFBfh8kebizPI5GhYzSf5pqwTFLCnuWBN4sZk67q29IK1I+xS
ORMylGQifj/8eMtsbRK/vXuat5hAQ6XpHwPjDqIP5yXAj7Wpiafyd/neHQAT4p3oqK5HE5tw2To0
kd4H8qTkcLVRCSwgst5+xLak5Mok4E/+3axRJxx25NrtankrP2i1YDI0YKTcJqjls1Dk0sEievW8
t+flrPbXn5JCd6gNpdvtjmE/6vjEiMx/EmABw9xKtNLRKdmj/JBGdB5my2P3EDrxeTTODw4y2P8/
B1NxEtiYoemR97x9/m7ahr4AeaZhSPIgNuayvMVukLX657e0aJjxHua2IlrX1AWnGG0Jr2pgo/35
+xoC0xA+Wj82h7LtlMvzmhQzrgMIef7naH67sZNvFPYElNqsjrBWJ5xMMpAXZQXp94Yf50SHRrAr
0K71eNvKURNuonSNj56W62kLhLM6+diJkIGKiwpHhYwuZXf0OqVquRkIZ3lliN/FLaGodPnjSogw
i69xjs68pYg63aLvTQalzbXC5jRdOySw/B9ewgiN1PxizQzicsIGSJKJTdZH0w10//ZTRPOGEtUd
2o1eyfioREd16x4VbepFyI8ygdAOc+HQ0CpBiUO+iIEin0OIMar0PikD7YqyFOUbMLdp/eCSAqKN
ebjYmnKA00eHgJ7G7pUDEIj+1NIO6Ma5XmgqbyTi7iughrIN+EszEzoR0d3Z2guEIWXhV1Dxn3rD
ons4lSzcH8lCfG+MjBLrUe5vS8IMmbwRjOXKhad1jb7CAD9UBlts9DURGzlI+XVxF+034UGl8yCk
TCsaHzLpYfH6A2CrjdciwBv1eevZGpo2SVheXxGzm6b6hlJrI1BFQO+nsdcdL2ryYxHN7iqV/Ms9
suXiMKqD79XmO/LPGgE9OqiE/wLuhYUYYrT+2lCnVRH2sZtxQwUKYpsAU8O3UEBbzb89WeifDNDb
GXzu+WvfZvfAXOvZUPx29LW+piHCdrfrZhS7znAm9rTVKxPLBli2SMDDOd/aCtPVz8gWX6C8Wv3o
cbg3R59b9KXQ6A/fHtjNu/zOnirVSdS/HQ6DsDk+pMHm4luYaI/f1JiVLv9ziYpm+4JMeXTJCApA
LBzMf6SwczJM+3xU29VIxxxi8pPYSlOVCCk6fZxMbTohKRULCr90BAU1WEXsz0d9A7MD5yhj+Koo
1jkAQ+mqHeEzFFbQbfMx/KHJKIbguHynu7+rUzDKLoEQp4KB9RrdpY6ZXWa3fliNll0wW7A2yc2G
rTD2eIi5MTakK9xR2C6kxEiSE/I8pPLzXW6duNO64iFBLgP5BPtgH/FB2D62JDLbGnBc+7lCY67u
0at9WOQFrMr7eBsMRMsc3M6lYyf9jv+9N+TA+aNn8+DfsTDD4tjXEHttbWfUciR6fUh9mF4wBmWO
oBy5Fzh4yN6z4NcLy9nzCqfk8enJUtucTL5NXr0OWRc0WoiKbVU0kEBj34tMNiBPJ1JElfmy8QPr
6GwaKWq6+BQd08sekw4pbb++gFisZdDQ/6pVn9qupy+8BhAk8iC4tATY0mVDYVNP2YC3hDwdnq8S
g8UKa7OdaE0HgsKRr8vSY74lZXcwRRlsNBXDwzmYUG2P8fHiTPQf3tV+NkC4YEL3jnNhaG1/BDNs
aoVG7/d9FxWjIm42An1fLaUSeV4k81vWJIPw0b9TqKMXYRU25TCV7wFuz5P7toP5a4oaVJ1aIQlG
BVONfV/v8Ur6Fq0C/dC/vf7ulsCB+8E/e+Cgo4yYX9FrQe+53JScFtrTEZtMbzKK0mSFXcktHnyD
omUYcGplANwZvcXSAtlQDYWp9PjLZFY8IkksuOmsvmq12vErPkq5/Amc/Jg04EuW52Uld+FeORI/
8bm1/sToKEebntAO2TKb3Yj5RtrxN+bfpAZ8q6ITLQfodleIx0BBgQdLvujqrKQxBdLbF3G1mnmB
dQVUIEltvG0B5sasAqD+TeYj7r8V4N7dzXYNTMCFTeFB2q5FZrbvBz91Ny2omMBfSFTuWoDHjG3a
UCUgPsjeR1VmzKgE+i7g9mk4eXuqGZEBeWZQtSbUcT0xTOVNeKmY8YUukyNc6QYEAKz4jhvWr1yV
cqtdWjCmNh5ZYyJuEbx8a/FuLwJ8trf96O70FAE69+ADM8qUSWcM1YbXy0tzJlVmdpBhzRPwLL6J
lcwgNZbUcq2uAO0xPcNvPZNe8Yo9SJHU+dBirgdGkxnc1D2tVnwgnAHxYamCKb2k/BEKCRq4lqet
EVTp9EKmbDTbbreEzcRv17SyIywT1u/z7P5Xxx9pSMqhdowv0z5iMHu9ZxOYsBW2oVmKcEpSz8YI
Xxz5WbgqQmz0tGVasg2cs041Qmx7PJlAOBYxgGNJzFpYzb8zhu/7OPy6wFlpzC8sXkY/i8MluMfj
nqymkrMxeRYzT4KMm6ltvu0AYgwsymDTiicTn3OC7EgCaPBIVNS9YCzbsTW34jz3VlJbxLgILlhL
8PCla0hzOXy2enJCxU6BaIjK4OxMeaEgSxYLSeTHO/v1Rezb7bV2hoTk44oarqiKMmUldFoXK9Sn
kxDyQPSZqSFwcqffyY5+YcV1poWz/oiSQ1T1gwy+kil4Tn56Ilei1IYicFJZGsFuCDGb7q76VPG7
2Y3vIltljjU+MiyTrGFvFdrVrRRmhjImTLZxFD/xkP4DNDgURKrodzAe2lw79JJLqrqOKzozukFL
2YmMlE74AX3onBuvryVKVN5BG9ivqGXvLU8lJEt66t87zZPqRzhxeqsxAyjkeJI1fjP70ecg/Pk/
JgSRRQ3c8Q+TSghlxiuQ9VpdPv+aIkMa+5QcVArPxtzm0ttwnxzwhPrfFY8MTstpNAsvyNBIL57S
F4yJ69yXNOqYy5hv4fdMpT9Uwj4u769CjCVdbCLjrL/ZOpWb0zWsAyZg/iZAGi3266j6ZWgFBd+e
Jjg/sIz9SM8FPNyrkZhFrl/Qa7QDczLuYHwQPNM3vNUq35qE+L4mMMhnEzCceeQwpWCW++6ZBXVs
imwrC+MKGhTVhIQR8FL9ykEhjnf+yr+fA6dQNx9NSSocet8ecQAMORd9mst2nah3sxT0FppPk8p0
syyRkHguP/megoQMYElCj8ERNCcYc0rfx5yq1+tNlnAbaHRt8y5U58Lnxw2SfL04t3GbWA6YZtdj
6kST3IW7onWEcprQTlH+HtzgIGIvImd5wsdVx3FiQDoOyY9LEzySERZLJGPXo8vyoPD0ZgZrl6Jj
F9rmr7ZMN4hxBwFRxU5QZMExe05KcbEiaDrYHyN6Vf4oXp6bBhQIiy+c9AsKocosp2mmYEbTkcIv
N4S+Km2CArvPJoWoFRC/HGgW9mwxITlPrgFDnBlig/o3eOZCpIOMQOvHg24hMcz4lNrhs88U6Aas
TFaP3kCc/pK/jRiopjZnwRFw7zm06nytSaAwjdkHhV+kEdmB60ajjtyOh2aX0wXgFI9bDzJZBevK
+ZUlCTmC6McxybSdaJ8ChjP6STaw00v3oM+sOl8wpU0kQ5ASXKeiEE6OX7O9qlIA778vJjwBfPjB
IIo3itTG3VRzqFk/GGzMhcKbrJ/ul/nARU/Ix9ftSCsB2/HfiXxJ6LzJgNS/nyvz/iwQgxkE7roJ
pdk6eDQO0nwvHDJsMyYFdb0aWMEcxV5BSeq6eM4R8NjBw6WFmNVQ38UHCPYfMrxGiyBaS+H5A82T
+QvZ1Qzv98NMcdFydE4GbmMu0/rzb+eAPXg429M8mX2bL6zqRnsVBn23mKUUChOco72jX3s8c2E2
pqkqam5lV9cgk+JVVBqB4sbHatA04qLe7+xOcGMH3zrfVe0adS01uzqx/s+K06so9s4q4QVI2q/K
3nIbbO4iZ2onKAsh5wD/Vu3XqQalJGS4hD8Mxetx34F0WsNF97xkgfYCqglid8SiFg3Ng9+L9UBp
M44cfy/FQYIRPulpiaqFjl65XbnPy7yuTnKtbnUOGlcSOpPg5cgBfXyxg/L3wRNrSllXL4iTpwPu
LLkqcvSpPV+4eEYbG6i5+BudvZnCKqtKRyccBzPUu32+SpYFJnXzpQowaQFcVjUjQuoKxogU/P1T
LYuHfZ/0Bj8JKs/reTR5Zhi//EOw8eD6tqnabpPTeSyM27p9Wh7AQmm4eWyHGNBb8nwdnjL3puAW
BzJr+WCF/VViLu8eRasDwgWoU+M82WEKk8be9NF/NkkF4zo1bRu8Wjef7bKmNWi90jJzefCrv4HV
rmDGy6RYM43WAUwUq88KUsQguH1+UjGLR2VnqbiO6ZfufW+MSFlXEPj9tP9FCJyhoQAFO5yL3HGh
B8jW2crzHGDs4DAyPB0kOiijJ1vHpNEC3WL7dWAfQSMW760LlvJdtiRrn/8geLRtDeynH1QNJ8Ok
TcySxXx8/kFzDKlYwo5hOoigFC6exBGqzSfNa7vDF3NjSXXwotbtDbj2nHPYN/h2sESkKR95xynJ
xoQSzstryPX/PbgX6RpvlPpyhguS+P14vKP2Xpd6E4ZcSo/v2B2MPCGws9hKSs6PLMc/gg+igs/c
9nea1pJd5HnRcYT7mRXBoc0wx0VsWpVTDrj2GLejkQ4vssr8ER44fsNYfwM05KdZfRgFr+v+Nihl
polKVbzCPXbAkSj1LCcxEy92OFTD0w54Lykn370KP3r6LT6rGcfjjPiMhOjDA+5cjtlgFOIsdGgT
6TqCQLF4ugH5U+BHjMW2gg9HIxutXJ11EVnFBVrFkIAZzL8VcbFYiViPELao8THW3f3Go7Xxf/Vo
h1qr8hLSW+WFn94aaIFkEPANyjFsxSjNwC/P2soarx1o9yH9XxWc77Ka+4MLDs7A2+yJL4aXXcgu
+j7mJng35jmcXyLS8jL7810oXlJwjf19WcwlA94cadtpSjrmbsk/iukpE6Hb7tGC0tm5F1mBXxjj
lInUs40tmLGrO1781Towk3C7G3dQHOHx1KGtQIyzhSuRmr+TCNsZTE/R0OmWIjBVl5oxdp3Jff7K
t3RvkQ0YAGTf/7G1yzqjfqjnfXhYgFlzgMyhWzBYBnr2dUHgT88BxAIMIi+EOxpbN2eRp+SlhqqI
KE/ZFfBjxeY0gc9LfcK5/wKkr/ZcmG2rSHVEmpOzgVB0WKjSMPw+6DF3GcSD/oNssKjC7+2bUc58
WuLF/G1YFTy7xle1bk4O2yUmnuCZl3bvVhEeebFDHaBfWQ1vpDXm4eAin6lXhlSKaB9tASCVZp+7
EP5VQgRUSNoxdKM3oo5REUTpqxFj1OGhjpfd8aIFaUQ6UxJ6Oc9MlThLx4WhxgeOv37rYOtIsIVB
/IogP/oIOJEXgGMiQrNzkf/htmKaSkKdmcOXKilgRsHAqnvOdWRylxCHDxyPNAkGS62xx/3pkzUH
Vmrh+3+FLX86WXxppnOeEtYCYbHKxqdwQeD6pQkpudb8f18yUYzesaXfxBt+4W00cePHtar1jJaA
3H9vHvTn24X5vOtabCyPDmDrb2rnuJyBYA6vS1wRdgexrHLELWuQGz5ur7pAfsp4Ga8WmQ2KLBXk
w1hRK6C394FsuL9TZuRra95Z8RogGPxNJpBW4F0rinQ9fWbbTYxb/4RcQgguLD8233NXr8LmFY+A
o5vKu7cvCWU5o0hEdrExVmeE2zxcUKu6eRZPZyM/mZgPglBOf5MBeNn1oRofkNrChTZo7pe3R09o
oiwzJ4Bl4QRlCfszxKs8DT5SijsDsYCKFm09GVzLvmHJpbImMJafGZi7D0bNQcxEI1dLZXHCYmWO
dgdiSChvlYUJGvMPEICiBg9ESKx2u9NGjcp76SFTOFrqqCgh06EsnDFbeZUTlg6wHhCnOGd1mhSt
yl2/IRoHS7/s8d9Wo1gNeoXMFQtujdfMavOiol7yHtrTPeTqcK/oCnUVEXjGD+J8SAuwTtVCBe5g
dr3rnr/P581Y14SiC+40+Q62UkVGImhq1fAaft9DG3ueTesl7er0gOihTsseIAI34+F/1MpSQg90
t3wPhxxD6Q8rdXv823n5j63G7AdqGj+l1b0T0CVWMGbTiuB75XEViFNKZlQYwdTa47A07VZTugDs
NuS6adW3QFbL1orlt/Ok3mGrMxJvx1Z+c6IJQ58IvHpusJizAUaIvCSz0ED0Hxn/6B8CIw07/CuV
FAZ0GT7+WbG5yH8uOB/w49WQpIOt2EKPfz7kASGvcXz1Im1Bprv/9twCndyHE9bQaejxLecH9XeC
1d2zGfUai4b8iaesAhQx/xC4ZczZI6i0e6qbnAvZwgCdbXNfpB+jhoorXepImdtRRLiRgfNVrcIB
z4b+83E/WJPxNgd89zML8BtKPogjwkuaJYlan4XQfZ2H6sZE5SMQDz6ViKdXHzB3V4oY/S50Cyvh
yBtaPRvhgPA1yXMJzugfK5EfXfClNI4HHNHRukiLV/2HlMY2HgXlAabRnI8YUCbdyDdRxRH9pX/b
Cp66RKqQLPTJK+nxRC5QQLGAd6AgvBvmQNULPAxlPh2GIr3wFFt16L5kv1wGwtfvzwZinfPsd4dM
ieocA+52N5gCJJm2h9GFHmFcpFiDqcXj2YGxG9efT8/9/P1a+wOvIokVFppoi8skZM1yJ0NEVgXG
QOtAtlzByOWRZTWOCuIUvMwl+xblfk9WntKM147ZLIQLKn7DySwtHOt/diLbpe7BxaJ5fIFT/V1z
hJxTOGdn5P6gUsJiz4UuNZZ/IocoEJbkpbuH5/i95NQmxaQCIodQOuP3Qu4l4jfN7yjovshD1565
mULmV5PF/GEIBQIUIIcAW1CE8stQXrDxP1KOURxzRWahiy1bLehGe5M1jW3qVMLb/jFWIe/Qexd3
579Lt6m4saVmRLmOjzSEQ/zM5Zq42NiAflvbDgbfFxUzR4YAvAPRJhYcrBeP7ZT8eRm/J3K9J4KE
DZiPomjVxWYhCG8ZfoUhN8ikVYc7b6JOZL3aCy9dm4/OlfdzPZRAJBEyQvP8YUfzZvuawx4WAcwh
NF+TYudwJ9eNzRFKXyEb2FoXNZxspoRfh2WHocv6y8hr9lW3GkbY/5h49xs9SlGqL2bkHs+L3mRd
j6WgjgKb1EmQTtXdU26E4uomXZNr0QuYcvUGq3Hs87PjjW6dtWJAP0Vh1309ken1YhnLsqZXhHNs
3hGdRUzziU4vb+fu5dg+6JLprYLHVqCQZy/jT9GeZ3btu+BjOzlRGJ1KiHdAH2ZSv4wejKN8cG7E
HWwg3BXoEku2sALcSxf4xn2xFvMFp9pCspujNPrsG0dU+lUVKYjvqthFMsYw7gvVrlmtAeOTtcdw
rEuJM4x1M2jh3e6C3iadlNHFwn244TRueucVY2uAC3VArakiYefp9F3SBurn3XWD63IRfhcnk77k
wEh8xpt4na0cqmfGypqQRxAcigU+cCX1murk+7TsW33QwBaofHXHgBFpbljFCG7ykxqSdErrijcp
Sz15NajGX80moo3EC/ySGEk4NKURia8eI9RSu3K9Od59sSvpE3Xv27JVqdiN6xgeMGVUMmeRS7nI
FfH78Dk8/tsKSn9CuXCsYO75tAcieaTAJVQW11I3s3K2MgzT83hFAZ3FIdXftrYXNj0Jzhsjtlld
0hUUxFH6DxmvL9udX3+pPZJlHoGT025F44Nr9nDB1uokp4a27mkNwY864H7LqBMMQchbBU2oXEae
nJQqyQ7c9VHmPEX5hzkWrFJAcDnDfo7ZEEkfrvRbQlsS7s/99dWZXE0oJLgq/YWZf9Qmpjaw+Jd0
zC+i6D/6vAEPbae0gO8clM2Ealt7NCDRM+Rvc7V847FQggPvOtf7t+V13nRsy60tBtHuAaCYqdFQ
MoK9vLsMrGpi1C/naGEpATxjLtcqdsU26eNNoKY8Jax9HkgjPOERDM7kXEinFuBFnpyKgAGk6mWN
Cvsq61eyuV1X0HSUmUqo/bWtEmas6lXFZUzMcu/9y8NBjZ+FMAxhi6ygY2djglP8BszBS9hPbVHN
SJVd579zsVluDj0sYZk5awF8XjHB92OIidu6+bEhthJ8rRZh1bovqOtTSmq4u4/zsAHJcluq+e9H
P/DZhyoWKk2sJmncK2yI8lz7sXpecpLJ+lKMqnsJXTkpRCbojd5LBg7BEUwN2nLpPtQ1u83Igw44
4xyfHcVAMz0AOfA3EHD067Mme8wsMAtZRwS8ldDFA2eVZis9kXU2txmEpnt4qZp1gGsCyQXk/Vsc
65Bc2D0zO3pkJUenpZfkVzRmjPg60c+/Wtf5qBJj7rhJC3dHboarwy/OZgTNT4JRr/i8MNq7kR0y
QzYC0oh0kx3K2uDep2cBk6kFE8uwZRCLLtjibu+i9N/j/r7a+acB80TLG6ztROMGpcpweQc5ECvs
OGUDSwa9UfZqDMhNLZzd5OeJgO2Be08ydi7+4adaOiO+u0FtxT0kz7gAJm4StsWkWk77otEpiEAM
fy46azFqXqF1elQI4Pdm1/FyQIs5NdS4k9gYSGkcT91KLin9XhSpffX5F+CeHQEal7zJnGCvD9Pg
2tyNOfbC36TlkVgfJt9VoVuhPC86yX7aoeHT5N59vo5EFktKP6Jcyh+6O43XLRfMWH9KiE2NniJ8
dcnEP36RxR0ujlKWJGnX4fKwLcmndK5M5G1+p4Kp/NWageNAMEq7KJZRvCq3j2F0bSZKrS90/hqZ
RcJbky3z2LazpsrN1/ZuL2UcoYCSI84p9qtqNTNW7DhvjlGV4hPJtt3I/Lhsn05UokvDupDJkhdF
GopFjpcaWyA4qlWJNnA2eqGEmIT23O842GpvQ+WFV1LuOSB09aKpd7lKBqWFOSC6FgLAH1+0fEpj
gGimV/5draHjA5VnlJVB6RYbTXc6gkjiQ5nLflvxaGZfk++VImFlKDV00aHu4fqLVyVVwmCCXLAL
RZ6rowNZulukXUlwG/+v78Juazc226UIDf0ybDdEfo3EtcP5tmE+OLQkmfkK6iDSR7ImEkzAZnA7
+30HT+V7qFH8+KGzsHP1rDE/ZMnM/FpETlhYxQ8OdvwYwdXbDI3bpjWFIGOvpY+oUPBmyzsJfmTA
BktZHrzSGS147k8AAzwP0UqhTfC2j8aUBd3y/NHm85wpIlo19y/37xtVoZjgZNPxdIXJ7Z6EviLl
aGCnkMpsSZzmFD1Gyeg6H8BV0vHvRpn1XnuWZRL+PPPBVGb1XJ+JGBYC+RAkrZHYriXXOPgBFr4F
yJFHN+gwLYVcuTGcAPt2+6ievqoPqltWPQH1i0/nN/CP3FJ5luKQupiFvxoDo6z0ZP4yBG1j8m6/
KBdd8mPzf5JDCG/Cis+1gYfoa6XxAURJsJBYRZbg82Tzer25xTjVQR8PigldHL0okDnC5Vi1OJvV
CeRU0ErojuL3NPPrLb8OM+Ke1cv2jqOTsNzPXtmlixcrYgkQ7j3aXvAo1IV/Z/7Do2oLrRopcg/s
dzLxp2jstAZeQmM2aaZRHAS8ent1Vwdn73T4qPAIEZZb3t3gcdaB0unuk7u5UFSkFZAeTKLQzcna
bwsZb47rcIyF3oX0N/xIGFTLB0K63SByHeTXk5aIPqZOGHzrTVm7PzvHMLB0+of2zkEWjmXktCvP
+oNgVPnXZUbvYf5ANP3+4tKzZ4My5iUjNwFo2F/67Hnmhy4xv+UDCrPSZJIaJ1VVjykj/KvhZAhJ
M0OdfJg3MmdhkgLJvEBZwXkUMWnvWWc6BkcBOATlnfaETmeps7KDbgAx7iW+xfijpZpic7HgLteg
3Xr+oDuB4nqIRlgBTcqGV556ol05F8M5mIFI8UqfG3SJnrM/GBCZ/9CQqtxhMhpCUwF+wy+6Zqp/
vCwf8xmPK7TuDX+fRC+yVzDUZ7pq10leZNqDl8lYrNznDyl0P/TtJYg9Y1y/3ISMoFkG13eVSM/7
Mt7cjf+pWNkpr1GVGlWAujgwC/XCITfq8SrH2zTfPRv8uM6fFfRFMU0y4qO5BtV/1Vt78rlYRSub
VzUIlO3Ml+0hTHXuaZkJQwRoITBegrYYipDztRELM6q5hwkhJtaDIz+ALKDTdKPYYFht7XV2uK2r
clvutC3c6tUOXYFl3L6qWtSHl8XDITyrSbVe+g2FcXAQd9eOrPuyX1Y1FuWsZd+p1CrNL8+ifcb8
W+BNXzRNnUTfc8xvQw0UpxA9/0Sz3S6+Ukwit4mQP0OPnM8VhNDCvaf8VruNo0wgqL4MsIm/4iJf
u3JTUp62Jw+jOHjPJVynIQRC9dxhscnSzAKqSVjxQFLxvGFeYN1C0964gvtmqZvmM8VC9dQtclmw
uaoSZcg912YTZw53hvOweLJDpFPmogGJ/VFcb6LGNjR3JtpqZeW4hl0M2p4ORmUb6aRe7YQcY0V/
xYLPZKpnDmKWZCzk806gRSHSWKtH0Kdm+x3Th9xsknKl384ak392CJp0ydaFMj2iMb5rtewnqREt
9qDsrCFbVYVjEb8cSzxM5kxbeOMfIbsfG+v0l+EAuBBQnz7t1PnlKnJQn6MQQgJY6ggCZT/c+b3Z
JG2zuAjY5nFMy5959Ng0YFpb0Q5ilMK/xt/j3AqTN4zNSaiSXK0twSO+4o4yWtf0CQ+c5iXpXf2m
iyYJ25t4N0YzmzuHSYzrcSy0KxiyRVwWE7rK8bFxaa0RxPCwqHKGvUWyxjKMlBwL9ZomGget2Z17
u+FWRrvuTznLTfkk7GlljvrdI87y5SPYgCUxWtunc01F1Mk42iS7glw0Xhy9z7KMXj3gT0PiBjvn
8SWcifW0rKpQYVYaLZIfYo0ZyCWAl/qczHIN0U6/4p0tuxsRTijXnkoOcS1ARSnZ60DOlphui5va
HPrMf6sUj1ccmdeVCeG6OuIK7l6OvMT4AQtdmOgN7WtKFYa/LG/3L2AdA7xLt2NZD0G8PMQFO5Rk
/8UixQhQgtAwnTBXxKcp3ksvQ4pMXqTaVYbzTByVkF9X3givK8RCsiQV8nBf7igvqM/Cw3AANMvn
KhaNm5pwn/5xkaOYv2Jgw42DLfI7Mpr6beLDKY9GROoUlzrWDluIelcbDw34MUQf8EwIATWxIo1Z
BGttGgVJLGKQfEd0Dh/OPgQkot2Yh2JYvVdgCLsb15Ek5QuR7MzDjRk6ZDYsQ7oKEw31yfOOpDCi
vjynnlk3awJvMA7BHm63IcumxJZb1w4jfnsdmY7K/GvJU9/Aacq3brHmLVCCGz86Js8ctiQwg+Bt
BjccukYDUUIX/34Wc6GtZIav6Dn/qDtcRZQkUQ8TnNSEQSMmWV97LuPt3ddOPmWgcGMl4VcOrpRD
S2HB6xq0+ccdaUvFWeYf0EZNJBPd9DF+IwD0t5Tz5Fv12bLHC1qKNyUwbv6yZSsTseAkipKuDpwq
vt+8hWiMMqz0o7UVozj7KJp4lz56tgDjGIq+Pl7w7QvrZNJ1zDKHnW8tbtA+mh+5Iqk3rflztQkt
nZyDRqVp4teXI0WdLXx79KoAcF6jC6Z8lBqU8ccMZCPtqF8BrbjzMX4pn3fjb3m5+QnKRRLVrF6Z
qAMz2l66Z/BURavUjgTuNIIE97LmbYbASiZWYzcxUkH+s2nPmZC/LtaN1ngNXnYDJiH+BPFmdDs8
zVb+zA7s4rV4d6OOJq1GpOVW01ck4sccoRALefosts/PR+Z+fVut1s/wPpuEbwufpP6ByQOzyK8B
3X5uLtC7yGLPgYILHgeifbp0ZRfAuepxcpFjxgSTHffxn3hZ0So2ULnPpvG0uc2zO4bpgz8Z0dn3
g1jDS1XJG7i1y+ltoLUlmeqVYJVrqooRTA5xPlUDYw4MxxN43sJA4ROEdzVR0pFzNrkNbNWYn0A1
Ri/2PMJJOTzNcAuokGATqWZC6C8E0N8GS3MmjPDiqMOrzwVtGpyQddAeNb7OdtUo8JlJSg5kCuBC
c5PIOpdDTrYbr682TsnF7NPkFlTcNwWE9xHkDTySCKM21Fn6V2VtoiR9Cfcv3JiR8unl5Cf/1cwy
2mSmAXybqSnF7kQy+6OXCAcVcO9BzXLSE9mczLzVszPXCk7nSGdtPDajxN/EnMAg1Oho/6YYAI/s
qt+e1FkREhRKk65FuCrO4uPJUi9+CKxrFT819CdF2G56HLBwESQzimQFafXum/x8qjGuzYdMgv16
6dVkPRuescNWLRil4H7eHBfeOkGsFQOhbuP7TRLZe/4eZeIE2pOcChusu8tZW91cS/incdUGUEBW
Q4gdaDqTGpWQ/ajme1pCaOR22P86Mi70SCyVIIzM5oo+1hd121TahM/dYOgQZ0b/ayrztL9GrWV/
7JalEJAQ+y5w8ETPP5sPqVuobg/nVJaCpjLLxwx672U6QbmctyvQ4R5E0KCr7h/Ua1pIceJswNRn
rkPTxUn4WwWB4s3ubJ+fWuqWxun1FsuWH8arm40U6jnGMQV7nN919fFoFYB8M3FyGbsb6MyGiIXf
JEK0nlG0spQo2jui/zd+7J18fV0vupzrLh3N8AcoDLkqRgeKYIPMdDUvhLWRCYokXvm2KmzCoPan
MTL4W1zutQ/dApSO13d9Fy/Hq5UctCuS6uk8WerYTrgvaied7glDXy5aND/5uLbxCb61wXXm9Ljr
Tw1eqvupIT4JI1DqsVazJzFuzERoWygerACZddGDM949S3+yBaMxZrP+wazLxtREjkRSzT8v1J/J
3i4d1lyQmgNg15ib1Q2vQDPFYZZhKeDXz16bZurH0EyvFFtf+t1+90FnM4UgxtNNtyaRmgg21U8U
MkQabobWBAuOVrCCHPXXBPlh2I7+V0kRSU+llqnA3FOOGg3Q4OKJZyAXvGEdAoqbcfS5L3UACbQ6
BJGpZUPLVvT6uv1HfJv/ZxnJ5HIb/rv4lWukLehEuwKx2ibVM23SnVNsjn1OiTSOYRkfFtEvphSO
xOXePyw9+22h0LRC0q33dLgwaLBwIZkDP5VgIof9tKV+hhufdO7IDGxeVOTDSi9T8m1T1GFu6uhB
2r3b9XqMhzTvw9CnHmCIF0WNdhae/y3HMql1YzQHUB1y2KMjwtDgIdKIHFLlSY4s7TAMZLSAUdT6
6X/R7QlIRFUK0/lM0EfSN2pKKSRGiwnNE/JX0q2lA+Xc+PJPJN8myf+2T+Fmmq7xDDJZPJ7AsHuO
gO2i7GJlLeAwGJfWP7XUmZlb1epc7ubTimmZIJblKN5GJLvD9f2Vo72mtApWgsFY7jIvxHefgOQz
4L2aP/TUfAm21kvh5A2RK8N3kixm4+hWTc92HQ6e5Y38K7hzNzPnFvCi99vVW7h0TCjQKc+JFExB
7sEtKJ/FeyXEI3XRQF5ZnFDJhLlpHmcI6Pjo5nCz2Qoif7zq9U8/FU7tAa9Yedj296kPk2wb3Fax
yVYKiPzBze5+ALG2gszEo07HFuzTmsyRJGsQ1obrWxshQvqVdrDpKYUcnKy0gWvOnGocrL4/CgdX
AxnmytoshxGBowBv8w7r4doFY1gdehjltzQjp4UZHd2imM/aRPk4+vgiXHxozRi3E5n/I8usJ9nJ
obRlFV1MZj0y8HQY0UVNsSVg8jJMgH+nl6TtdZ+q4zjslCvtvLqmdXxZXAwfofgHD5j411y+hcOh
FnQ3KFcrpLEIou/hkVKHBGQ+fxk0gGD1nCIDmAcg4qu4j+8GW0wJ8dMA6GNsMA8kjar9rlQ8D7ZC
krrbSIsplLhIo4qJI+ne+9RTkTkd4k42jyawggaLUqhqbtwGy+41DpjnvYMgbQJos0Qr5HZzcAOx
Jcuc6Oqo61x6zIXtAy/WtdnP2xGaN1aTAdJMgudiaduL2QdhvrEIEwCZ+9eOC3JStMcMduQ/W/Eg
jO9Yii6RjpREN71q/pdgkEYVBe2KV3fP53VTgAds0jzcGVWRxKngthePZdTIAjq0PZxz/TnVguO1
BQi53t3/Kh0kTstuqhJVD7aVKKcCDA5vYjptlvbHhyCYfVvPFlXwh+Jmnhp+RgJfAWhDnItPT/2A
08euvg/FAEosBmW14e+6fHSNz5m6YrMFxQuMMSBR4XfPLTwFV4ZgX3spM+K0er/cfMATB8XCN1yJ
rgnv39+9Wk6mEjWcSTVvxtNCqP/OpHv2+8T+1dljmq921JDONs2iL0RL0ceZLh7JuV5zkujQf5Pu
Zf0LQXBG8K5qgdUMR6dSQCGVAUbxprKxBleB4/tDO3ppQBg9rFnuQD9KjrFR8/rX1tIaLoI3BBQ2
WArx2M90vRzLsm56pTD9vhgWn9d4/OTXNQyLtnqgWWQPfXEGfIg+JcX7qn0t1Q2IilfUPxxaDLTS
hh+FyFZno4F3KsnE6stFKuz+XN42Kah2zzlHP8AoNPZLld6NQRwsoNKl9ha+fWl9TYhkeQ5rQc3V
m9B4U520zeN4XQAl1ihIop/6Oo16lRnRt8Xb05K+UbOol5h89N7LYvEkziG1R0aWX2e8lDJQZkfn
dRn5mIW5Fd4DVknJ8hxoMVQXU/3xDhmmIcp3kQM5WkDOQPNxFXrvZa44owRPnIQCdXeeFlsGC0zU
jLeCrefYa63WaUbCNszrPQpM+HV/qPQQuU5cGTbWnviUO6zxx/n35Ry3pC5R8nj00rt0/HO3TVbz
IjR6beRsSk7M4tqz2DS7Z7qOjjUzumaBrz2hUGPpnyIE9OAg0by4KDln2bp5LNvfFAZojJUuW6xk
RkPWfXU+39gBYRW0Y9ea7ZD3iMu4V5uhE7gU6YzIpdRCIe++3gV84rzxSfOP0iVn9u4s7p1kfpQo
hqpDntu/oSYNLfUC6k/vVaA2gD8Tw1yeMiO1mGVvUv22WLVtg3wNg6X5WtxFoPdRJybKJt0p7IZ4
PV6g3MhVJHjQf4wPzpJxMMjFrshXpHfKZkcAr+14HLwkS0MwHxISRDgbEpNgoqnHcb1zHSKd79fY
QTVwvi+KtvxBkyPQosrfUPUuRj6SJSAsqYu639TbwFMg4fZP89KOM30xAUbNAw12qnse66ZFfGIO
OqjR0o6c9O/bzEFlsJxo3VFWQujVDmDcKLop8KZWL8wpeEk1DYPBq/fUqS+/IlluIoWysQzH+2oN
tux1SgtfW1nsdxeWEXCC4ctyfpbiAx95zxfmM/yioMLhmkI+ZKd55I1/csL1A9VyvQ2sNT7lzxrx
E9xblK2KV6FT+Wie5aXH0dwhMx59pKALgsr2FcRCokxmF+MWhIBmooDAbkVYCXn4RGxHudylgfI/
OWVkmb6RO2s0aQ3RN7v5BJPFtxroH/D430DhU2e/iCXYAmRdYOYcBYbkTPhzHPzfh3A1OFizepkd
LY2XF2/BKjJkOReVSuxCl2GDgb9MQptRufcENLT/AVH1owhxG4O4cecbRWRUqAcmMhTIXnlhG7d6
23QBd860U/mBTg4QMaSIK2QYmr14l7qpgILzWbP8xM2SdyhztdRAlufXZdWkUu6Dh4gqlhWI3jCf
K6YQpsGpULewqY3RiyxMp2+5IIKIwKDYdr2gW/x5Lz+7QPNB+uTqZxW45WvLs6I8icC/JL7uvWdX
3pmZKZJhd9Dqx4E/oDqdptcDQGAPhZ22fixypBtmWL73OwpEkDAN2mgfaav5Q8QXdr/85mJ0v6wX
+dyZ3STSilTVl59VFsC0kQBfPVr1KY3Sqv9M6CRz5XxwcUUUISa3ek9QY9p2h7uC8AoUVmNaUVzr
LM7TNZ1AjVOfL7nPMrQM2gxTMNHGEy8u1LSxMOvyRG3ybGaKspL0vtJOB77HwVtnuNs2zFPDkIl0
QLJ2CHHZJtRgrxMBa99UVeW4VUbDKetfmCJpoluYSPmM/eRUNx3uQhN4OzpYgcbqbR06LNQYrlem
Z6BopEdrIeuXRNQ8PvSbBJms8WW6viZ4KWtjRPaRGqyHOLMhsYq27B/nD9LaTIdFS7YoORXlyXCo
/5kauZLLn1l7VBbxwtJWmGzW7p+gITtO85mAqIYViTatknq+pBwyBWaa2WLT5wQ73SbIcWTiqe56
cONl6E8GZBCMAk1OmEtBiMeDQvp9V62pUBI/uLHSq4CZgnfM4ULd/DkZuSbV6NwbJmXjlVCn1CLX
xRmadDRNYeiN0Zf+0B0mZdB3geBsXDJ+09hzE40rwRrkCwS9KhZ1CCYLrl3FK3r6xi3X+NdzmqTq
heSy8Y/B1xJHgfoA9O+OqgLeC6W2Vys5HM5XFl8mvVKrglFda81z6yYqbAlKjbAB54cQjREJynrz
bXq5+nonffZaXlwFDb4nvJfPPppzXBbr3NypMAksLBY/RKdlqXZMIs9jnNHBBIvj318z5jhacqcX
xXcNdI8D+gjl/AaxI1VLpjIYBObQkMTg7365K54K5qvRV1t8rPqKwe8/FvqqvFYmv8Bhs5vLb0xl
tKpxArAxf3ZeV5CSNsn01z+LDx1Z85BwOsqzzAgcgSV1HhSQspw2Y1iX/2Eekmavltdplqms/Ej2
O9IGt5P8MT9zxJROrxffRrPPHR0w92oOeENpySTS0CNbl02I/GmfPz9ZikWNCxtd26m9cHhw07Rn
k3ZmgkY6q1lr2v23wlIDuMV+nax0WtOXolPD+wD0UjvbkXqCxK8K/0XXdCyrkfTEyQ7qzDeggLXH
j0dMsU5bCL/hJc/xQQ578IAGNcwy0GZ4MeYqGLJXV1Awhk7AVwQyGa5aLoelBoUQShsBPlpNjiXB
eeSF8mHJfnB7FBMSFW8UCPAP38Ysqp6bg+pW0aMYOEZDHgL/lRA9y/NjZBKlp8iJw7kyIzzfMBcY
nKWuuGX+xFpbSylPKLlyURG/IoLhXk5C4xyQfWpr9/x2gcXWnYurhOLp7JSaNwOOYOXJMtu1xzay
aYkTSiY3aueFn5NO7MhbvjLwsn1+APctsrglViE14vcA1Tmc/LmoKNJw13Z6RmEoaty8NLqQ3s1S
5yvy5rqjkdzDVA8om2y3T+ZVU8JuGjlemvLRiEvlX/G2L8QilECoqH4PuWBU7u+YRPX5yuPO3AMn
KSdOy1Dn/rzjGsaJc2D4Mx7oTZJ54rGSPnZfXsz9RINmspMQC23G9JC/HeCSt7jLn0RRRD6I/UFM
qFNs7UCtef26RWlkDEGlk9aoqR7d/bGP7MCrP3UHi6dqg8LB/n/H593WqY80h7az/JctzVR9N2gj
kc+/0xPnL2VXE7ODRsYuxU2bZUPOdUB9XucLMXjreBiZJwKJ9yWizu1opR1ELcRxZ61wzUYjxAvG
cBfrelUO1Q9PbPxlOeCkd8EsO0cMOq5GMgqQ8xCehHh7QWcWnD7uS0jOZ3g+d0jBA4FFWEDcz5T+
KFFFdqCeRzc/tBnnj22vBWhEkAeoGtx3WUXksH7fa2kRGX0MjFxNFiygvfQS6w0EVLLIc3Tl+wbp
vm5f3YE4bTR/ftY1Cj5z5P2Q86WaxTY0lg4BHVqYcXmdchgQahHbi0u39of28r23TUN74xhZH5yq
bjhkhkbjcNXa+m6csfjEd6DWbCmJN0ea6UjKUypfNqHCs2FCNI6Ch2HeAI8/0ZjY75fqwpslcngB
XGuz4XiSM/8ynWO9b2p2i0fP7QgAWmxlVEjo2WP2cSvHhuEmmaUSwlDSaRSTZzb4cTFzFKCmE49O
Fe8Wq2PL5wz7SzNc0ufv+LvRFZslnl54LQNeumeaG81EB3rH9fizL8DOsLnBSRYwa1VvZvcKLdpY
1ALE1Gwl6VZVAycZ80BBR0ehsnkvrYhEkEJN09RbYDP9bSsUqOme+U8clJp97hsLjkk42q9QXqaY
D6b8tiMgWZrdO7n8nKTTWOVRhtilmL9TW8TW/m7PGKmUQxP4iBTIsepRCGP6f17uEUXFJ/TVrf+J
kDpAlCeSC5W0aIHd7o/3gDRUSPSCpRMh5kF/0WIsT+CW46QMOAZKUID1/ATekHOIGCiniydWCXaC
/Sw0gFnW2ZgAtAcrveTCphloqZ3d/sRnjhKV6QpPFINbLK5oMsoLT5NQNSf2syfv8Gf6XcjeMewC
dgw7N340Y1V8lHKBIr6uJE4Jty2w0SlxNo/SLNGcUtvKFifX2u4fnc4iTPue7oohCUG444qJfgap
DfxNJYAKXJRYZHKiOFKph98AQ7I9Lg6MEw9c75MvFRaeeLy0CwDfxaH6xITnWfucRbzjOK1hPY6q
KK7GPfw+s07GY3cXlFOy//O3j94Mxv9rRuO5eMExn17btjour2TKyTyoat+vD/toGz7WYD+WLrX3
FB7cbN4R9UI+TBJdNVuvKPN0+XkyFz+6MN0DEkWyDa4UtoUdsysgpgCsgsUcNOyhJnYko9EpbH7r
fREQ7Q6vrOX/tQcj666YniN5N5NbooPcB41PfMOkvU22VbqKbNsl+71TKu6Ntd48puW7dussnSUI
pP1Z1DHWddLpi9vKF1eh3OakKU5vAnV0hI95Wykv2RAAMIqUktQ7/8wRB1ST7H/LojG4mDg9AURm
pk8pxESLljQ+CUgKheu/T2bWGWe15R2/WjCIOLEhVKghMpMPehr7/jrF7q0wrf8T/MFEG5WQ4Wpi
3xTJF1ZdmmTM1R9N8DAMuq2HkKw8g/KivEiwgPPbZAhT/p4gAoEF4VGAvj5IMWtf7UAIo/6MKf4d
2YuWt5D2lTlK3jPSxbXjrKzD3w4JfErVseSpLKtAnd9oY+Mx8Jr2pVMSdBl8Q7WSjYtRcp6nQ0NA
JHxI4CsKUeO5PBZ8yRwm0BBEIiltClwckUusa5lfoBegmfDl38DC+GCLBySBPjIXqJHpkW/A3wf5
Obg2IqrXh3RunCvQzh6jUGumiC9XRZOBIVqGuAkHadUXx7v6hM66NdxP7fH0hVoeB5cBsVD7p+jG
MQggJkNI7j+6sE3Fp000PGGT3RP3lVmrXP2BbBm/3Byphov/PWgbnWm4SKQ2A/vLma74QstptpTB
xeQb5SM/jtOMCBGLQFvD8Zz1/f8NlgMuEyg54OJ5ZTb3XFxmeQbl5T7YlZUG+a1FgXj/RDbD/NAx
bu3rMVQicUG7ScHIxsXgow49jcZpQPFS75pEKg6wkMwA1TM/lSB/wd85+wNKu9YSN2zGaejpKfm4
f6ywblXdMnPAV4No7m/jvVp2TKu4SDTcMvT1i0Nix4dZIdtM7JAlli+22/tpW4k5wHH0gq8XkchA
Ez74TmwBrxd6UnmrhtETcSmogndnYxePpdTUhsqXlrhsg+3dFw+5YTXc0tF+CRhx/GoofAGV9aMP
v0kwQpwXLnLkjf+1IB9JFkKVP27p6tWy0aQyjJhciso4YOwopJTup7x1/ew46yiQyGWtCEqc94Qp
yup60WYOhNGnHZJM8IpUbefDwjM72ZgP41r5Vw6/JoG6FpDjKLrq9QHrtO/S9+aQ4QtElaXv9Cty
XRiIUUNLY2CrwA83jv6Yr/KbJ9dTG1CvG9AVg5M019OUAtyTyFq20O2KwujRZyuG3RDtBf1ne1QQ
BxiteGitVislizLh5mbkAuWoqUMUWz6t7kspOV7tKCRWeugl/O+4GbOXm4NCRd212bq+VZTiNTnz
pYBaX4eqii2T/CYzqKV3NrHk5pfq4wBp5nZvgnZg4x+1CLbtJOeSKGyG6vOrLAXaWrKPpe9VlclD
Qugfm1LFpoY/2C5UsYnAGdH1rptw3fIafXx61CwFFUQmOvtObs4f67LqrdEUp6KjACcBMmePXg/N
7zCc0tNge8XTdl+veuY4hqgibakU/2zY5okmNOJ8ZaxwrhfCC62Z2UOVTF9jrXJpeBQ7gnFKO6X9
Ybq+4rNEDHUfTn25HvzM3oeT3GwiUbEd7j2vs3X31Y47nz8F5hldRmAMMc9jFAnmAq/AaSkSkMPY
WBklvKLfg2v/SWNYlJk3qoyoU/8O3r8FjhbQsMW20unZk24PGtF81y0AgjV5ox80IEnVZ9DksvS4
IKUBwVBw+c1yMiJYKu4xfYtnLqRbWqW7G27X8LuXNtO9S15D+PI+jwUIcOkgehiRagEC8vDF+ojB
Uu9tdsJgBWTuFI3PiAc5ch8MuTpiSqVLFZslzgpreE0t1cHHSnBeYw2Mgb7DlK1gmFO0GZ97sae9
Pjg8wnTCBWrXjlUgkXVVCYVkN6xVmtBYqj6hphjCQr+5Ne7pfzrAYwwR2RL6CPPcYNviWXXxXgZg
YrsMWWCZ7r8BqWG13tkVC/+nxuVq3Sakjui/xrxUXDgHAuB6yq29f5Z4tEcQbJX5eNDYElFAXRUg
C5ScRuOv9QR06d3dDD7VIigly5gzWT1DaJvxPfjZabGCkfelPZuZt3BF54HPW6IhFpr4UnkE3l3b
HN9lRPxn9FBfcCgtvTSi8mV1B4AyGnwXz2GmBYR7VUl9jLijjQgfEYrngpuqc4O/Z8kcVAlDsVsF
HrYb5WyZu+2d01WtQt+7Q/ye+vc/wQAIZ3IxFuBe/zI5EnAFszQeVYdEPubVbNHd834Ghvcwxqor
pREp6n3dNuQ1TMGtL7WQGRqZtQZjS6AWc+WFJ3K3WNRBLHESHIF+AU0OGe9evKyWGuuoVk4s3Efg
H9lS3kFNnxzVVst7TrSaDW+UY9JKUNFCkB5/3npW8wvSX2q9trW1hVzS9gxeitx/oKAsAT+cDDMJ
2GIcu4oawwfx4rlhocjZExW8QQbDXmyHBE3xpJblUmP1KIH1Xcn7o1H3ZzmyW7b36enVOZM74iW3
LYB3JeNoKNUSpnRExwAPwh9yLJDUBRCl13aRWOHykkmSOM5IRTePf5iGQUKX/wqKCGNjZAGekQYJ
ptAfujxbmYsmSIjfor5HOZ5rCnwykUy9jtn/FMTbqbJxPji3JRhmn74Mbl37kYGnshI8f+1HXj7L
Kr82bOS/a4NzRAPRnHr2us8b0iEbOc0QJor3hvEeJgJFSkbnqRaunfRFi57Moxho18w6p4DMa9FM
fpik2Sew9OagJELPMFq+CA6vWBNCIpC0wqqrwkg717qhxVhjA4MT7ybpgflc/Qbgs0JB/E+5cXir
K7wJ0DuF41d+jYYT/d3JKw+M7J23MrBOmcZyiXiDvwlhbJ7XIxxH4x3rjHOAQ1y9xgUn5dpaXd2L
8fNckth0Y1ORKaoNKL4E6fYNSrY4awm6Q3dJcYqooDuuDJrN3e3SAQzFocsmgU+KIA9K9sDaXPjo
FVrBGLPfw/OS2CtJXCR3ONoH0hDKQzm13KUyMFqWuRhpsQzBMxic/aiCLsKKBvr4gtyNbd2h+wW6
xSY7SwlqMruD7K9N8DGIIp7HqUwquYXNA2yHQU/QVz+q+M6ArfmnQA0fjEoM9JX1FblLJQJB43zz
r/GDrizlbfeSWqmMu3RDVX54jpAUeny0pNaUts4RiFDu/MEhmqoRnvrphzn88haBENFSW6WfRb2+
1WWZyC1RWgpUvuc4MCZ385PU5HuvQzVbNN3cuEsfFJYzkgBVSEEE7ymIcwOfMNACJcEeRFD9crww
XT7Wc+I0bHqM4H5dT4HfXNmgXJ8w88cgX+p+CyH2Qa12/pfZqNMfXJQsZMITCHS8QZgmxnaEQSl0
Oc6Bh/tFaC+QG+CKMSpL5DkAzXWK5LOD85rq+h3w+MKQQURY2FMkaD+O3XgkCGyMVmqM/MNEQL1I
pXGdE5w7LRp/TDNWol0p9JluZud7xlHD7cISmIGdovRlUFxCQT8ovUOxP2wM/ycjuTqPYed3U+2/
YVXoxAmO1jj2ieCnP3f0QDNQmAQ9GaO5wJAc9JM2k/Kmu1s4xDIMDm25RwQffkBmry26C6gANpDq
K0re6vBRIL23myzcO1K0+gkpWZUnj3nekksgOxJotssmDRJW0YpIW/hxIATczK2UQuRYInI/PjMj
0ylnyXITK0KGtX3lGMR457dZd2cCw2nyo0SM7TqSjdOFTUL0z1Ll/XEkLdrrEXBwnwkB2seGrghz
wJMvVWVmCwOZBBOHTiYOQje2ndSazh2czM4X4FS/XWcLREQ2uP+sBXgxyFn2x9StSYqj1raMFV8a
9ocb89cLdUONHMy6h7MsoIt0LnwM7xiNiiv0g4t/o3En+nDVQteyldTC/yFV3fAH6dBqBXpsHng+
RUYZjGtuu7YBYPo8vM5lAYNQPx3DU5vE+ge5CO3td8fN1vTLV9DNboEeBrzTJ8mlOOr7HTmdVsbi
PuJ4/M9YGzrIGLWkZZD8bSuXj7bUlkh0GttFdQedj2xJtYZQhN49As7rgodeuJwD4FgOaU9p3Q+6
oAbRNjVEXgxkUAsnrO9T/NxMDBxPNHi1hLpChhdI7lC4fEvq7ZBkn1P+m8ioNLHS9le9L7viLDII
OhjmNXQzcKq9+UHRfcsHlJDwLd4U4vrWik63KjQhHdnkN7G99FZbhum3M0O48CEoAZF3GZeNsHAT
Sg/h2CTFCs4G4XJvbnCOCJrxKDdki7w3zZMeOB+ORrT4I8Z4MqEuSZht7diIdDmAJ50f/ax522j4
dBZx0jB7KfuxT/V7PPRO7iMyYFNU+BpSY1vCAdw9ctPzefH/+vjeDEa7QKqo/WwwlZQPcf0tD1Es
s9rML7GQyO7OX0PgW5Ss2bKLkElABEyu/ZAyWHZm9QO0zcv6qTiM83DUwkFHEUqIj5nYhTQN4VGy
AgXQTEdi65r2nFEw1xp80OAFySA1U8XsQfWcAbZdLzt7Jf1PWvHckf0Zgf3xvXRSr0ZNgLcykpFT
ihlIbMhJXL0nPyTlHDJSYt94+BjTmV3X3kAePh+T/y3a1WdEfmVo7nB77uz3A6+GuvuFq84pvEkz
jVbrYIM66REic257SoFiWq4rI087pr/+Y3UNRs9nEsR28H6kP1pXrmHPjH0eXRHGdEeaw0ibUyOm
d1mthejrBfbNCFJ7LgGhup3TIE/wj9B+fE24Lgeyx0YS18vAo373yeKw4TUb1GwqaW0eZJaemPXp
Ki4rvQGF6coz4Q/fR2x08gK5/wdAizRATEFUC9w/nUGq3sP1GiHID6sXQ+aXDuzudlAn9TYYBheY
pVGycTN6URzirQj5nRWY8UBUxKAAW+n6M6rU43UNIJ9itts2KCwo4f8P75A7J8yADF7qzLGfOduD
RxMiiMRyiGqnIQvRs3iTQVKYa8HlSjrVbxaUQdLJ8iC/k5TEwGbYNc7GFuaJRIcLoMFT2Pe3QJu5
dpJ/qARLmD31aVKo6aeMzWZixq7rqTd7JS7qgsjTYZRfq/TZ1TUFBu+QqSi6UaPyNXnppArkYfHX
E89m7Fb8EOSDefosJW7YAR0BNAEoffbXfWj2/IQ3dfGr7lgOT+OX4jhITrqoid+xAe5EbWp6jXQC
sB+B+Tztut2GEPyxlHtBl6Ba/RX9GSP6p/+DJUcJGc9tdcHiLuDRDHij4pqSgPy2Sc5IrRAZdRQS
3Zdhr1eSkCUGH0hT/pBh919ov/qVxQif+4Jk87SLlab0ngqYdVpYk7+vCQmo1rGIhYedx+LFd7dg
PUnYy6RHXFj8JjBMGtNhLRQ2FxFuGE0vA50NAckv+IQtUCNKmbC4EO/2ltXPUI8bRYFBvkCbz1m+
vNHHBsKCZjvnOwvcxYvg1XygchgiMtRfjipnSuODFqNtqeyVAmxIznlsGnuXdZ8LkZmvBBuEVUvG
UUAbteaNc8LFSsmIANV1gJXJ5eApi5e0s9uQTW+JdVAvXgAk4BpvFX8Qg78H/JIlNhkBZz7kLlcX
kgnCkw1mKYRJHcITPvrUE9AKu1GGZwHKeACA8xIP3U3QAQoM7LbacbnNxM/PG4oq3y063uoXJ2Ep
GcICs8pwo8eHwEwtEksNGJpqgP3mwzzxrVVe6gyuTtYaRBDlDTarZp91C63hit4J461AnsYRjUl6
lB2pcVytw2ejcShXl/qAqtl6obAh4JcwNbaNrywGLQ/fzoW4Fru36d5+R6CIPwSkmF/EiJlryGhC
JEPPu2TEYycC/zIjRGZyOQztE9GxrkJxigRrrqHtsMEmTT8+SK+CBVEeDRs65Sg4Uk8BkXAUjEcc
yY1eje4UBAyeHj7IxhGi7Vwt0HwhCN3bBnFsQc1vivQ7YTTsPsN786fifPxF3Ut3YcpbOQxxNWuj
B7YNSXC0QJ99AlHpTGPceF2koDcHZOFrY2ODJcysWLc0UsmXU2bnxbg8CGZBRiPOHMma3VxNv4qN
qJm2BLQ5bOVSGi3fnMKs9OtWVaUejInJvecA4uWMQBFhKJmvK+bo1kSsUecRvnmw5iVXcKQun3Sn
lrSFR+WtUl4o5+Mg9XEKjGCOIXiFccWu/aCFGdh/luAVfcVm1TneZiFw0he9koHJccBXV8SyaSdU
HvSLzUYjcziCxkz3mt2toTEOpW0V+pghMmyBFZVXrKe/w0HnU4CTFtuoJMKxuhBwbwEk88jKqeQm
nol/fn8d51KJh7XXCfmUfIwYT+qf6jXg16zO7wwJUYScytVYsmAtJ6dOLCCsSiTFSEYBpUbyL3K9
/oUARKrWWDsZ9m+0uOMsM3/eaXlalKi8WT1oJoQNvIkaTpp3wwwN4vrHLdG/CQaynLrC2CyqXiEM
Dl+r9t8NKN2sCMVHotTk7drZHRzXgnxuXjvKUhPBTmx9/jpcJDGYDIHrb41GlKpJbyekiVI7cg3p
rfOiWXr78y2mfks+eoX3R3UT7I6scOpKnn+paTxlIiSnwcHmMi6B1ZqbyMUsUPzwruPpgtz2Kzry
Jz94H8y3HfwE5NTs89nP4R/RSq1fTL6TK3mf+jR7hUpjyC3JeHXqmIbFhZ7hgpfjq6Sw9jpfEW9a
5t5RZDbHFHEHf28JbwwyuIcX5SmLH4Qfxlkll4G2Wl+h3ARw8QwyKH+JZEY91I4dGjYTEobj6ybk
+F6xkhTrT7XZpTipFpUWxxgSupLiljCvZx/m7LAHCmtGQDqe3g5Psf+nQLq73T4tbDwTW52UDRLB
J7uiPChJXEy31wdZ6+NbotyB59WpFrYH97WtCY+L6NVMwmN4pdYZgtlzSo/Bfaip7xvO2lewKPr/
kGPrqNdxiNwIX7CU619DB4gPtVlF5Wqqe6VEY5hnPN/lxV9ZFcYtN7+Z2pe4wqhuWiCCMOeo2e25
j/fZdt5Lo5TPKlIcDzzrZYiI1XV4GktTFOATHr+z+SVEBcXeHP5OX0aVYmei3Ar31dQSIzjVTimg
Fbp25IyeawijQZ3raH9abei0LcFTmf+3xF6QUychsh+oHnxYeuep73mnV1fTCJ/G2OnQS2EkhWyL
FCf6XXtahUIW6PCxu2BdhHGUxzdz2G0sSL3lfY9O8d/cuIX7qqsnhSzy93jQTmNGFxB77LiMAzI1
n55Aw6Z573Ftb1C11csJbTX5So/OKd1NNwevcQtrluEoKjP4PdGiVqV60n0sXn128SB2IsWE2L5d
nvG2CjFxZ70AHAP41F/t0fX0xQkEJJniFiCu7W0cDCpUDYdmW8PxlzH31jH2GVkFQUjEyohtmfsi
yQfxQBg9oNQJaujVhjeZs1gXI9cY6FETiU4Ui7g6A6nvgvjJ3ucrXiefaHA3Hk5SnY5wh5T6DQ2T
7GHICDw3EW6ZDS4mgwygU4tHPh8idVJbBZV+qrE8PAscrz95D27zOaeGbDLgkhvXA1susLTtbJyE
LEm4jrJOfWvzF9bZSRYLGySATiX5dJstNl1D4Bh97Ji31IKRsALBI1o9LHOhnZPBqNJ7WwKXcUzo
EQC8cNgU2Ku+yTe0lmoZUXCfd3WZ1nHJlmKEmJzxG2+Zypgy6v0eDXSj/TOb6c9LBJM6uJQWV8oT
4DMgV2g7mk60O3ImDnvNK7UaMclPMQPo1dZn/+O+F9u7iN3s//oFE83oKScPNO+zGVXGAdpH9LxP
kEt6qBIIcT+jnz7yyy+9ccDqeGgduEPbboe2c4XFIYEJJqoBQSO1e+IMo1lYJyAhx1mp1ttC2/5i
DHDwVXvWevjJQ31Cj832K+MVXDrNv9a3zz2oX2QP9XfwqlIMep2YUneIqUfv5akakLqYo9wgY7GQ
iTFMkSpcPu9ygBr0w8VEIAhQB8e3DnU5MnYlkbP4zbfedVkqkqrKRINz/vg1hEi9fHwisxkr/VUx
UTd/+5EEKg8vtL186IMFi+bB2L1dKwlmfk8dkjMVLiQuFcgdVvDd3LqhrHXXQanUp/cf3ij1W6BX
UyFwM5MVX/hZ2wWQ3xVX6sNXaqJ6kWg0VL0cfx0n9xsDFt26zuHkfMCzKa6zfiHlHxuSj7uV5R1f
mMDYgVUDpWZhXcrOD+r9dclynV+9kcW0Nu10vyB2yJu2J0o3I/9XeXIQJ+xI5kwvMFay/dKZz5LW
hSaaNKX9TL/fLb8iIPTrcJG37zNcdtz0zuR35OZqEApH5ytUWpfzNSLPE++PhakSOaeU1k65Rb9i
/0rhpLhAPm6ViRiHFpsHdk6C0Gs9iVAKEx5g/tNJIQbsyNn58PQzz2dYz/C6R55sxmSSr2FDnb8v
gOW/fO0SPIz+sCwnmPF9oVnpGNq3jvfpD9Zdr8mkPPm77/9o7h7ymAufXfXXljKCTzeOZz/QAd8d
ACqylP45nBxsyJfo2R/D3BQjGiK548A5th2MzNSsLVSJ8GmFrm66F8q9OaeyRwKl5bRadz5MuU8G
QkX6WYdmUIqtzxUlVyyVMcq6sid0pzQLX8fsMvxeqFirDkzPO4N4X65ot5/ZmN7Yx+NID1UIk87p
yAamP7NKatZkUDbvf1T2kg3rdYUyElAICGEDhkjALwjGp7hR9TEBeIPOuizKtgAKita31WzU1DuK
4+t0NS08Dd2n0TCiKwDU1lQvO7j6Mfj0UXWUOp8REzhHMWegzpUC2NOBaRoBK34zi2FMUyywh/CK
RN6Eg+VkW8TePICtvGLdQuIJ0TiTVLH9P0ctVFG52QG30u4juYbtYJObNR+zrdEGtw/ZIuTr7VtU
h9IGMEQC6XmWRKjpHfGXto7DpHUjS09ZZpvVD8jvGwtPEuzYKHxglDlbL347rbrN0Yb8I5zNnIzT
eIBO6FcSkLiCA6KYLCcVoF392kXD+U59aBI13HfyFMb3R2RFshMCisKisb3S0wPB3c45fSRwCk9P
PATkrq53rV+8SjsL83AeG0cb2Ncp3dCKtwUgGwka70YFtILvKWuoBzlmI5usGE7i0eJ3kKYZPLOo
etx6ls0YFwC+EnWakjBZkwIJ+txRsWcXT1OgFIZOdoDOTDyStdHUXq3VtSTOEIfb/eYR36vD+bHW
sG98lq3mDIa1dzmW5eyGRsK9OhUza7lYZhrb7znH7DS0Eqnm/wMd8ku6F8d5ZIsOwD6StdlSw/0g
IZqsQOFsR/RDuH6csni1hWebtg/ubGe7v6GkQZcfdYpy5FbhGqG64WzUw5tLQyhru5jECCG7Py8Q
nRJhjmZWpmC+a9xKya9Ofh/c0YA4/zvi0IRKqhOrQEYA9pTm8REOkrXEdJ7vRRZbgKIvq+/9Tvgu
A5dRrAhY7oTSzajEfpR+WtAGKQO3smRbgrrcWLV9oLu0VdiREZjop4P8+OnGzEjd+D1kwtWM4HeR
5XIpWJvTKAFh9Zg0QOfFmKb0dJPtYBganP1kgi0EmP4XXNO7ozSmLZeIf5dtE0FXh1GTcKCSV+6U
zRQLOdpNPs1erewFiZI58wFOkZjguTGZRBp8u1kjy09NssJujerF50GMMZNgdFf629HSwmu7Gvk/
K6uqPoLGQxq+XULoFlpGSDDeYDWSNvzqYTP3Fopmj8PqTnkySAeoo2jKyQzwEVrsJL4XidR2w38M
1ZB1mmODUHf/zi7fdHK6Tu4NTSnFySPA6o9aBHAZRn/5bAvPs+4y9Zm0u1+jh9QRMN0DwPurE30f
jGnTF3sERSC5JuzAoChdvd0NDsZWni9H98xkJxIf78Bpb/Fz+Y5lm/JSBi6tSDfgWIF3mzQUnDMi
Z3S+JEZggtR+gh/BsmqB+z3xvr0oEslHbNuFHCq1Js+WGaj8uQIMONxfYu0/dGdW/ExyWK8ui0R0
OKfQgOZAHwZL21c5KgjeXHRJ/REkgfgkNycr7Zso0E7T+RBtzwT0aKp17Xf10FaYlSrtH96LXAtj
sUA8l7+jb4Z7F1yKeNGQmmIXcVz20Bbuxf30VxOwCDk0Vy4ZSBU0ZR2wJyjXZcNLOq2tnawVdFA9
wpOxwSm5sXQtfcs89qD5KkhtSlLwLAUT5YrmBzgwEOCwcZyLNqCWG+vtR4mZCczdNY4W/zCC/2kZ
h+vxPgIPjxjs7htTEDqSBoFX3TMXcOvo7Itwq4pNc9WXaLud4mC5ZN2YAHSLt0cmi9bnw2FWwEaV
E4E5s0PJR2G0rysFaxA5QDA16lUvYpPYmJEjxUXiR9qlM4rRxE1OCDrjtfFqVu2WmEl8iMljM/P7
N6kmyicFKOGbAHiQ55SFfbJmSk846FZw32JpqfenbOpWMgJX45hVhzt7QKAnGVI/uno5yA0Az2TE
2/Szd5nZHZKEUOep8WUbWjWKqFcUZupGFQyo5Kd/wdtIecCEzhyoFFKnwiw2tipXmlG40s2jzb63
JV5QjHbTb7Imtx1WJlCryEZj8l7bQDOXxt0jR4oYXXchiRaPIK+HvGzb1ldDnha/tmj6PFi3cOO7
D4PBay30hofdj8m99L12JP72hHqBiFj6HDhlFAM0XR3Vv3wvMNw8oImNQr1exxwr4FMMtfpziq/D
pHlxKvC+NXbiSi+B800zdgS025aPWgZu51zB7abj4jtmYaLlmLRRB+GHzA4hKcxgT2gG0b3GH8cO
68K+HXgWLBAMNokNEf5C949Jzs95X2LYLhEIOTaMh+XPSksNWnY6lghNxpwGwELJqKh/0QH8/2dI
WMnUuAN7XX5iDCc0sYdz1fmcUKgvJRzokMFrN2rPl5/xxQc1X+CovSIP+U1qCoXsVCmPMJ8KYemw
3khrIzG0KkHSagPYt8v05C4kXIHxHDuLfJaxuJNVyimIRWFH09ABFLkQddHm6MpCZQEbbNLNdxPZ
cCifqi3YSeY5XWkGkPKspyFfccrE9Y7DZ9/X8sdSVkJTUxilirjieYliRd7fVx84atE2vVAB3Aom
11OCBzIcBejDSu6h/jXejJkY11Sf1tnbnIF+WwxnZlr7fXRWFhrATbyDxOei9AZeW5mq64J0plBs
QsKLG1jWbdFj8zzGZ/hRYXUrT8g3BenKB9K6cP3xFl7/Au6Rk74WNgNfD50lcyRDobm5FxSnfLF4
+ad6YWGoR94BiaSXp8zDPezdhOB4nnp33Zi3C7zbZSoRUKl96KUbq177R+hdAxDPjIS9emnWS1ov
sEWZwbfLIGkGlqu1n0Rf6DW6oyKy9ds9tcPT7UXI6uDtmYcoye3xfuT8cYSNZ4YenBMPseUajAFg
3OTy3iik4Ip4BYto2j3mta1l0Vxim7Zx48VCOw1Q+Gah4NRVoJzF7B56PIoErQ5xkhDhIQYNvpZw
w/3rrbI18aCOF+IeVbFp9SFTcQKLMGP4yRyYEQaxJxJYaHPiBkr2iOPCVFjz8OCVUVxVVBh/S40b
TtjhIbbscdw0Mm/Siry1qs6L9ENLhL8hmxWo/iQ8Gq4x/zbLvfm3WYwtVr5q8eVgu4+ClMZd8WRv
2FQ2zDZuels9lmEqao61tlXZwb1Xx6ROBTkmZJMGihSKg1LKGONl8SaWnHAAtPueioqFumt9Prsd
8jW2pX7lItNbGzKkQKMtf1hELWoopBRwV4RlumgWxJwb1hVLP1mX1Z2Dwa7qjlmXLWBRi1pg2PEW
6f8q6zaxG2ai6/n56Yjxkhnkk9dBC/2c369/vIl1bjE2JH4wLZrMtpsvCMIKf01AAZvRzID+IU5p
BScdFtEetqlfBvz6FlzTDCqNKoxsWlY0xkKCBRcpNP0dI3M9C+MaXv9usS2KGoUzDekwaq6MEDfG
/iac0gSFzQ8owg+c0O2w6MrcNIX89zhbneSJ9o9i4bKLmT/t0erTz+0XNIAwACn8q1ksXVkwThl0
4b9LOpqoVGEuVn/KnY+WmXhD7iL1lEUn+SQ5TxZxkSSGzV+nC19c0mCW8Tjvvv+0+JTuu8Ec5ZVA
Al/nQZCZDjr6Ny7J+QEEO0Dsc8y3OMg7oBMamUx/b+VRMaYuBV3ANetLK9/AR+izogQ34II4Fm1C
huQmN8WvqEijtrFry+ckX34DANKxRSSGZRmg33Tq6DK6pWp3drDkoYTUU4MBZu6Asmsfj4slD/Wi
Xrw6YndEsr7CpbdWR92l+d3MVUqbsUU+88Q9HIAqotb2jAhj4vkyIFCv1LGmESRpLeXhw5AfLu+l
cICxs1206HlBVAkUIhqJgHcGqT2gMxa3M4EwcEnzM4ADgHzOMVuuSy7QrFS58hpav45Lz2yvTknR
O5V/LEDM3IGzOdfa403nAdJC3swCjG1GRSk2jpU0w68/vNhukx/0n8RMIOTWhyfE8wZxJXPJlnN7
EG4VD1hBP0yCbGjd9ScAY6GH6stSjLIMTK+XK3IfrSvWapFAAqtUG6LGDKaao1hmaCclOCPb0GqG
Mfv5R5o2j09m6eia1eFdMKb1AMEVbWIcs82uWWjSKU0pKdhWEycZaz1X6UizfXewPjEAcAR2TywR
hMdP7D2QIOTk7EjAPF47HHwoX2FUw7crf//WFdgMR2gpPwu1AyJsZYYAao5RE1SMfCykgYoRfjxl
nCaWRoYwQYSFiEea6gXmbazhUnJUL/ZC6Sknu/d3UvS6Qw/ZPTl7P4oNfrLaiB9CIKHbMQonzs6G
Ll/9t3bW7vCOlthmrXz2CNv+kqbZgWLaaJ+keYj4b13lyjV5BMv6Ur8kW/fjYHjuqma+//je6lpa
XPzh41n4KOUVlRz93AsY5vJ6/wqUf1uFR2C2nn/Eqjgb3UBRO06+3kHgnvjlSpJoMOu0O0p8FeKH
yfDyyvdRx29MhEc4ojQlmzF+etvhho8H7Fkxo1Az70eSOGxJBdt9kFpfaBt6mQhLTVk26dgTLvOy
fd4O7a9Z632MXdIb4oicgcp0EtqBbL6UCE7f1Lv3kGvKMXZfW8I5mxyyYt+oPVoYYYrkLD3mMXVc
y4Fma6u1nj8Byl9R94Fg9juCgD4DEld/++Y7aWyZOcM20TOVIlXbvs40+zJPacJglISCEB+RmxOx
uHLbJ39qqKnA8h8UTEt1nfnZRAptWM18p0ZpdFfzusQEisuAYpRgSpuzKjJRoyVatAmAVpO7EQDL
lPI6S2ZiLI7C0mL64gdZU2JAWZlojXJZvSZG0wPzWn3CYFsMMYg7qQ3yrI+GH7mTQto0dsdHFgwq
qGJBRAH9cjXJRQqvNh1+hfWkNfoqzuVYpUhG9nzv7x7BbwdgO4A3Z9Xxu5wflrl/1axCb+lILH+/
Lt/MEQ1yS1syav+X3HfQlRBy7CfIG48gqgHBnWBa2xtxKLcraNlbPbxELSAHv9ZkU5onPYwfZMBV
8rZEeMxijoyHqpG1Vk4qN6oqai82Y1mzOJ6moUNzJYVl5ffOP/RVfUO1FaL5k9X/zEeuSIRMsRBo
J83Z5NBg693Lh1oo2QGb8G5MzsXEsdgQctLasC5WF6/oME4ROuG7EecxvOhmK9nElRS8lBCMnl07
ssJc9aYqRq9s8L6B87YD2C7EFZoRijRwlJnYJg2cicvQ90cZNQbyxQeHpvSYZ8c6yVSaCzQ+yanW
dykRzXTWxJUUWqxLjr/E2wDMWY+fhZB5I4J8cm3UwCrQlioqE4yKjhNT6RaNuPIN/1RZr3TFWc7/
6w4LcKinqu7I2byEEFydM9qRSYx0e0/qIq+HfWcIYJcTAvvGBq2OSIGdaW/l+M9B02mNFwJzATS7
E0sFolMvXTANGDvCry0fYtK95Sfm5dcI1xsAAwqPmuLaiSTwKal/hgRvac4orSsvrrNjSojwYB6f
R9pSawJgT2YL2+PZI4s41g12AeA2YFJwn2/R+VINUhhVN+DlwLEX2mu2Jt09rR8SZItR7HpXeGBq
jcfVlpNeMUndvikKEKkoLysfLzS4o/ScFJKOdmhFU6LuX04vVGlM3NOMOtfwp831IrWmAdoMWS/1
WZ52mnZNuBi1tRpQbz40Fl/vdYwYo74H3UKrXbgprl35sNdoHj5RuDqyMynE/XhYdwd8QHY0bT27
dEL8abYiSx2kQAifpM48CR/3OGDES/P2Wllv4cBf8oG983rq0bHCXBZuD8SDLCNnjIFeLI/iecUS
l2wBaK4v7XNoobwgMhQ6MbCbUUDCplci9FY1a2YBfFrHfmTAdn59pTeKIyUZiv2WB01tSeqKaTW0
E3cwmsr1OsTVaDxKjREnzYkVf6+91NCrfj+38dmnS/l8OW6v1vtqXrYoSR1HVUIutaUKcSZdm7X8
f776Nm/FxyL6iiYc92+TbQIUpm3rRSegxME5QdiddjgKB3FxPxU+NvXtYHVTboqQOD5BMYQPZvlF
uZZnWirA4y5t32Mjvg0jZ9bNXUssPlgEESR5eKqzkGmW+0aYirKB+3sLeZjyuPRF3m8xAE+y8zfC
YQaixgwdhQpfyExRAjXlOupbBfPRPSAasNqONa9pgG5SuzmlVEjbUe0SolAvcstg2PIo8xucEHl4
bqhyT3euK+SR6YmaTUJ2q0nxSv9FXBlhYSo7n4en2sI4C+ypwB7B6GbSyLFPgNlMDMScrPfWun4a
HgcjZ7DQb4l3h2Nc9AEm8JJMS4UDSOX+/z5Or8oULGyyTyidrolXMIoc+X5ZyNvrdn7qkRdIvXrV
q9OyI/Fgos4qR/YUP2z4dFH66/ptjkLwJIHXjh/9Dm9IMjvriCPjeTdlRuXTmGK8W1Ykir3EdQNn
+llb9XsqKWK1U8kwvHeMx219OF/QDcBuZGF278qnVu0OTPPYSfLKgId6TMpwHfw/66EJj8JTb/VH
SJMJV9nRDJu52ZXMJY+a7sSS8VzuoUeXboYRjsJoUZ+77pyQcJ3yeVm4ALvrUtdEj22YA492sr/7
PmcOiWduWNs3XLgJTcSummTUlQRlZWOPInVrSZQ/rGTc06Eb5Lt8QymVMTEvFtxu8qB67XTPNP4t
yajVYfHEuGhffMU8Y0JHF/WXO04B+0W99U/Sa++TXb/3gbb51nt1c6jipdHyk3k+nd7G+PSIHEJU
NYagXOp6EaG8C9Hu542S7zXAvnlkUEJ2xWzccRrBYQqW4yVC3PmcdGvxJyhvZNxRlJq86sx68jRY
G+7PW5Wwucg8UXSVq5YZUlFcxOefuMmc3ClmJ4OAvcDvYeQNRI+At1ElOnuJKZmGxEmRUAYxrZfD
uUF6pUhaOkiE3Y3agrhhc3sVto2zTV/rgBOTtXLtkNaabR4NK7w938Dj1KyzWAJP8PVbMZoMRcVa
x9Xqg+cMRAycnlEyRgxuT408T401xh2qGaNCfe13hrca7jIgz2mVHFdzc9okERcHORrpLcqECEsO
5eBDA53fFA1Jk73WVe/vSkdpPJtSCdKQgLRZ1Lh5GCuCfJ+dWmCwu+ZFToc7N1pEP00isNlFgKWx
24BVay0csdW2dl6LFHNRS7YTQDn+n+nd3meCAFcfUZ92jAYS448feK8sOfnpE01EwTW1hwuPNXaf
Ego6EFdLu0chldC4Ns/JvKO/dslyshd+3O/HN9oZBoFMKkNyZEcM+zH1MYYZ6fySaCjlPTcPftyF
TihnWj2mkSsXT+ckKZVHko9Zl60GXeH1ymCXcJwzVJ94qglGT8CUpwQVExt0/JhYYIjTOYlU+NVA
GBpoqKSpIAogYrDqc8cIJSHVoxxWQbzt4wtnRTxpbguYmlRFhdO1l1fTHewbcp5toP/cLOE0LM0l
Hspr9jr6nS0bG95NtESBa5g0wsJbLKkgxJYPRsqe/3jyAqdDDBFvcXQksPRPuMEEwOjRrhTSbIs5
N06TzptargOvbFdrkEsf8TL+wUcdJGgS4bjjSkBTJmbgJGBj3n/k9JY5G9SJS73ePYQrPe84AShE
FEHn63kaKAUvznhhfe3Rh8qfmmnCO2V5MYoHbz1cGDMpaeaiPVHu8TJJAFxyMBTlLXrnGDrGy2SU
CpgayXmlQjVkmZugqhi9K/7W6X9Cns+Vg6uBEEYoqnotzsV4ChUeT6Cw9js5wTOUgUnKtzDIZfBL
t4vkA2IsKaw8u0LvBitw/yZrLQhZqK2/dupKXx+cjkWBdpavn7s+jGvXI9PrUL4IluJYWuTsBDKv
kGI44GY3Jj1xK9P4u6YeyLRQKWhLsIa2TUJMIETW9D3r2Fe6djDC83RXMOI5621HCx5rRcuPwyH9
P9KWRE6jJfiQeaAD2+fx7Z+Wlz8MPdVt2GNQQ3wg76lMKWadqFRooKIdsUXij3POAD/mEcgDMOjm
ZDfme1J4Wlsi/ElqbJnJcpuos6J3WvXpg4FNDcVqe8QglRqbL0EIFsu7odKZOAYsyk4fLYnWKX3k
bsvWRbT+JE17lk+20j7ZI8afZoyxaJvYrIKcQZ8ESgqYq1m1dMUSh9Ca7cLV9tRslfkPoYFjD+u+
awt4o53qYRmDszY0qVGkFwfUheGl8AbT5JQqA86M4mVk42qWDRFtf3ktpwBl+JVKDf+dM9sryVrj
Rvy/HP9RCAPgqZ3r0jhjOINKS7gtxrW0fOVzgHobokMs4xo2PWYJ4vfhwPdoXuTIbeAf8vjYfCjy
a4EK2DsQkCfx/9M1+4mjHgXJyyjJbTN2tv+ENpbIr94X1yRp4SmfsHzfp/IteEoISDrEEWlTpLYr
x2orNskt41VUmA97nt9LXr2QEbf4PmnbpTCYlRs2saWDHxBhwNrLxrJbcdbMsyhXXSmkA08Nsqw9
YBuyIoBoVtnv3sQ9saUO/Us+O2Ywvf6A3FBcZF8WzrjDxBQbmmoJyncuwPpCzAlHjODFZhZFE/sr
TYn/ZtoNht+rzlh6KMdmII58UaJi6jSVfPjCmLeTsmGHpGAgp1wDvdwiUkh9epm5gILPnX27abhp
JYcPqX6MFwlKMx2XzM2prf6eb+DZARo5OfBIn6IEfKZmjCmxzYJExej4pqkbuvexJhD8L1HC66wM
HS/s5ZH91DFCI3jKqL3cQE9YGFyDT4R2Xxihvy8lyF7CgQRMDmECqSFE+X5enQWOEsGIRqj20cFu
k24IiXyMAUwq4CTrI+uFW37IEjZWm0PZMYIoKBKfVrokuzApe04sk3GauoO1ubtjEI7Gkui3SVSb
TduL5nTAWAtfm+U8FJ3fgTznhw5Fvd0UwrfYkwLVoyouD8hQsq5SMT63m2Yhx8oth01cjGFRbsE0
YqPYV7PledKn0WB+pLk3Rgq586uQL5OIFU7CrhsQ2VjRRntlGN9YqG8yVylw1kpTR4NFXKX7GqUl
5ab4gu0Vac1NpjJT5a7jg2FUVt1kzgA3DUpUrDCwjfIAYQpe/V0fy0HImWY7bf+IDc8bm6628UmB
m+XEJPGAnP7nuTJLUVCQZvNc0a5W4PrSPbnXMJ3kDCmmpGwDaKvFah2Kw48+N/+xpXTt7/OvN02c
2wezccRWf45eRKtYjjGo5/7pH5fEEvvZr11eUoeQSz5EWoXYlLDF7MhPDalLvs6AtscF7QhqX2C/
xzJJdxpXh92peZQ9BIDhdUqA3LR1Ys0NNacP3GjKjM2RdescnSEMLbbQ8uVY2njmdvvt6XvlWG79
upFt4YwWyktLEwareWn0uqjPZYefrI42A7ZqDifVbXfpugj88rIj25wr5iu3mY6d/eq1xbeR//a5
YgqZKy9n3pJc8XukNR8gsvVH9dcUaWodqiQW91goy4MruHqAzVvX2Wm2AnIkD7T6Tmrpv5xSM84T
vp6Raqwvs5/zFufGXR94JSkMiPiCR5IAE7X9Qi07kmoBw1nKyLHkZaB7gHE2Zm3GTv0Td7N9qp7h
GtofU+Uw6Mqb7Bo4VNh7P/d+NJ6MWiYwlfplftw2SGM/+G8K5dV/8RlYgPLknJglWFGETbjK+rmb
4uFcnuvolBJsm05Ssi9/+/T+PW2RzlET3Qck5CFUcn+chn6HyefWNqKAnFttH5Et7X1gmEyHFi6D
f9GAjxMyY9hruHG3xgB/G33+NEF4t0kGEo8wHrO0Xsj0IBSbRcG4Fq/mBwf/XZbkzyid8oA+OsBX
lw26pG+X2jMcGbZd8dZU/E0EEklxJSzEjZbTdiAzri5YwFSsq9rx9Mc14mqEtVhziVOV3oxYxdSN
oUS9tCW+WetNhT9Dvd3glBo01SZ0NuiENd151Ws09kxfzmdGs3RDf6XmHGFnFYjzL5F+GmZEUXZ3
5TFkokwkgDQDdt1vttXv+GjQL5JhgrZxM1UOhRj0sCIpi8vXtxo2WrWrC3YvCx1EnuyEK6I2vp7e
olBCWDrMI+FzwAnUELNwoVm14MH0FdiZYz3QcmyWJzUigItv0cULr7DaqUbjBrMpgtvNSrnakCCH
pqnXn/yEwj4O+8RHkTOmGmBk6ov7yfi9pWPameYoB3wcdGwWQQ6Mgo89tME5MqqeFrTxzO5IOjW6
xxycI74VGqe07z53Jeh6AUWUjel2hMRtvVUZMPcqsn/cYbsgiyTRuqsNw5Pm86ZBKkjNcg80fcp6
xCEf3LsjNF0jA3TsmoRxxOcX2UlNDdJfJUYCbDuCMS9QF/HjtmXfKhw9ZSUAN9IhxOB+KvPaxO++
HHY5pMJIWVcjyB14xA/YMIKJVWELzqIp/DU3RvapWoexGiKKEfmhinZXfOmh1LVLq/HNXFhFJnfo
uFgQQaBQicwUMLpWIiY6FnEhwqcXxP/2RRS6w6nMLO7/7dU0S9IrdM2x77TFBEsugDRuyBmr/BN+
FzOMPylqCuQiK3KZLDqZx4en/uZzgNIkS5DjNB+OHgcY1ReiYapBITYRtYrZCygK7hEYVsRwbcRk
BMiQoiCGt/GeB/3Aem0H0s5RKd9GeywZj6Aeh9ReU2zGPgGRCtJ7RqG5hOFklX7/klJJ8MgELCeM
jgGayLj6rCsMpK6WpW1z6xXFhQG0pmNE59IHFZISpO7wSKfqB55Anz4n/iBXBRLAi89u0zTOOLc+
XkoA3r70Xdjiv+TQd7vEtJMOBL9J/JXJ64dnNEr8nV2ByvPAUYZxNb7z8cdSB+E4j1ZOV23LLBjx
ndChIrvDmkFBywdcq+MZ98r+3l5QKEQZXLg1J4oml6r96xjz4OqWtkkVg7ApQKiflRKWL2t3cqpW
XPE52b2UqjJzSh95xPBpUy/ovu70aMgXIuamzLd9u8wvpuDJQdVfwgMuwFEEFhVFRFjhdzkvxC+c
hFYXTYXlyjG0FJatRlDu97FuDDs26PV5YZoYOGK1/6BOa5LqtXRKvJBJtF65a1cz//KWIy4bGhfT
j7aNw42CrRZRQhp75txhRI1ajqdRVLSzbYCvBc4hm0Dl1qAC1+O0lHvYyxFy4eviOh+el+vXOeDE
Zr7ZFCc/IeH071obZzf2liWoVEk9d/eJLg2XOzojRHYLr4LaRYkxsSxn5Kq/03crwRUBqu2SUJAQ
rubVXGRiwhRVXm62VSQMxOmhZSx1lkSEtUyx9SDfADWHGtRTJFdxGySi+WzE5onlAYFya29Z3oHX
nd5snOrVibwFhVjdkmOl1TmkpbV5zAFDsFGR3SiT8SaLwD6hafW0W8AOsQYk69bz8N45AuCYK+dV
QmitRoGc2uAWZMnK4eKYoRH2MZxSJmtZyEzibwIFnch7RQ9fPxJSFP5ms2BoC/2yhBLOHtLUVuXS
Wwgcb5K2RJGXUx0U0RcEYUeA90rlZhjgCLTDeJ1KE8n6VyJZPTGENwZ+7xBKy96466K7TDGsThmN
zrDNvd9e8+l10iHBFNnPqnB3a9wQJxizQkerzKA34zjtWo5DQQA94lo4hcOj4Uuqkt3dTiMecqYU
GmDxLvHdk/BYyVT/rsLIfgvEzCUGKwlYXKDQxxF82azh+KSTn2BTDpdujHnKGblFeH0eAHgHBqzP
3yMVbJrd+tohP2Na/5AOFlHr9o+oxVrK+QlYVnCjP0hbVQW5sYWokQQIxMpOfgm//SXFNm9XA0iD
+qZ+41NiTbr/at19asHpTIPs4Q19ILT0k0FxfeZKKJC/Y6+rrBBlJZIUQgFW3iMATfohNlJ7wkBv
zWjVPmjUjJIU+a3x2VxeiKW5s5Tfs0W3j8bHlpAfaE0mmBMku9htLdVVxYl7oFgGcdgPwI2tVInc
y/X3d0n3sBFKURzpL8EAjs8Wly6TLtFc3Cnpp2/6nFCvEjq3NMWpNai6iTWuAPix2A4KTLgtQRH/
zShhrkf4tucfyAxxFHrhsEMcCzOKE+8Ddu9fLVIZpKl367/035b3vAPlhEYTBn8Tpv+KdW8d7Cl5
GbpP0Tm6wuWZzDef/x2b5MgLzFVriSqk29MGggZm1bM6N6EpVsg3In3g9szHg0eL+ETpbv485YOq
0wvOOyj9ESemWmXQ5iqSGI+jBN7/reWs3QsufeMZyo9cqB/goI6f1eAu8DYbvgw/Qb6WPWKH83Dv
zA40t5/pCU5oWagnpvqVcymCusinqiFg4dCG2dNO9AlqmOxmaDomC1KMtJvy3UF0WZq/v4dwD56r
HXU5yj8pWwXHvhHAttzAUPZIIKGppHgth3vHMZsj1VP8OxaGbyIHAthG4k9bjWk0nqx0J4aA85dc
bbW599pv0dpXqUOf9EodfObVb6fA/tKhvyKay4VDnr4tGZHilrTXnmjDJiU8ffGFTjNel1VEisNu
RbDcuZ0yvsi+/qxvPyUOGS0OvkLN8bU/VAdafbfEGSxYEH9TIOwZEtw/luyDpGiT0BNcpUo2PDJR
yRLFZsjH+rKfIP3RqOX1SPYrxQsAPzx2EPiBI/vEyH7BeHxqmCVPnELP4tkzJdBwOS0XWmzoG/BR
KTGjbL2Zz5UQEwJjjkTDrjGlxzo3iHSNwEAbyVITcoqfG4UVJzq8NcOJumkSqvzcKu4IwcdvbAL9
1KlzGSnd1Iw9pgdaHygtbmVDcpTbfCNBLACIPZJ+XMRzVfxDebpt4b63QlctbOixWCWrVzY+ztNZ
3AmjtwG/MTLoyeC6xHz45FgruAt+LXXhel06J3EY4/FiaTncHtot5FfP0LuGE3+pjWj4quwDM1Az
J2AXFIwpT1r5STuz3RDb36Vvel6+XSxtqBC8bDAk6hpTRyQdMguKM0vuURbX6aMfRMkdorYSSil6
3V6wBUPWyje3ASCjp+fMZhedZew53/NNrcVCv6b2Nwnh2uMJ+yoKkR8PU9giFY4uYAyxGuJ/BpiN
RmRONrvbCeaX/zYYt2Qw7vcJj0L05D4syINfUQKKygf5M6wJYbx3EHFawo6P+5obGjTrnrAu2X7R
hBrlRJ4MxKUBw7taQXj4JrzOJVXbFudChDV0VkwtLszJO8MUBn/RY5ELTgtuHe0U8eqNpn2KcXj3
fEcg36kE52wASH9X9P8zH9oiXbwI/O/ySAz3MsqoDuvK2fGv1RxDzONxSIo5nGUqHUV87rKLkOe3
1QtGlsZGE8RAV02FVcmoUEubKDpzPfbCpIEUtdGuICn5CPgeZjsxKTT25AJiEghKGq9T+qG4tQRz
GmQlxecUl0MdfCSMeP3jOszoFOmQlwYqrvaAYT7DUDkI4YyzVeSpilctDQYDU3onLXP9oRFkl41g
BlELdBSEWebZ3JcjTGgUns8Q3kFxWBf3EkIOszrPAf/HItKjJLYlSdhIBudJ92qSc/pa4q4xsfuz
+uu1FIBT90xEtdRQmVtrIuMMsJ5hJUjb+TRY0tYR4SgYG70MDy84vdJPLvrxYgCCxKPH0XcuGjz9
sG5dQEuaA7PD93YLygOlKYIWtQp6Xz7CRH7276hkAZRsbmYxWzsButpHNhhMp4ZW44154QzX4KjQ
pAFYFjrMwswwxsR38eURiyGlUarsjeEhivXs96Y0Y2VJlN5sg6xljozmie2XjWHe1BHoP717nl9z
yakMvihhGsRc9474A85z+F5ZVqtSfwxSXbS7Xl1YjzUZs7VoAe66XjB/PglRuUE9Jp0t5CT8KU30
+P+oNnbKIzrP0oERygSxjg7ihnEHEvgvdQ48EhYDEd3jEjHT0VeInkvV3/byHlMBx/t7VxvXaEzA
e8Gmw97CooJdtJIfr5MLuImEfMgk7XVc5ANoxDmBkeKByiNLzxsYjWYcLmaAet4oezfdRVrdEBor
yDOn5mI4lH+3nIRCdeGDID8SIpZoaHPyBKkdU7MjB1oGKesft5u/hlrydryfxZXeRcK9zW8LXLv+
bheJUQqReS3IBNGKrLZYGT9GmnZU8Rc1nmjgcmOkUI8Zl2ASFJ58GWJyrRcC0eG1JopjW8ZbZaSP
Dh0GOuQ4uLSonIUSAIJb4olx0y1BGQSAGoh8tZnRkwLgRlO0TI2PF3II3VUN6WmNX6u/TyU+hXIj
yUbmOL/UhmsuxKlSpPgnbZnVTVqv7fftIHgQVKqgq7pctXzlLpCX/Cw+64XQlGQSiNPrhd0evGMA
y9k0mWC4zoGGB39YlQZqbRONja8AbDVbYEx3Nt9GCVIQlTDZyzzrkbO9lP+HeZibcG+eKiFfztGF
K7erUgPbZAnftCg9267teiynSkWeDQO0ddZK1571c8Fl3MONy86XwehMD9pMKoCmMHmJY9Jbc5PH
XhM0DnlUICq2e8iQgYLtMLS6zar8dvnGBhEn5Og46LHD3NfUW4JwIoZsH/h2F5GKuAfrE31VSyPI
3bhSvoszUGv3POHdXqnAt2HTNH80yZDNe/Fo+92MEvTlK3TBRePduFgYWgb5uGg5VsCxBafdkhaJ
KBxE41liitiglwyH9hIxADjtgrLxGoViV4VCwydlADTCvo4wCQdWSITC+LP58okZtcge2nPN3k55
Y5zhiplAA2b2zCCjcRmhsn+LyM1CLH2eS4Uo3O4ZkS2kCViBMAxbp5mQFQ/9TCxKZYEQwnKoCUwg
+caMb6Iybg3PLA60uDGvrREJBuAJCgJNJsfpZNSOqyrDNamE81kNszIF+xXAX0Ck2B29wb+rHB+3
MND1SEB8BhyIR6YrF6+y7NRo/YFl4x84w7ItaxaiFzVUsO+h0rlOQQiHLvmlF/7hMfwN6Mc5xoNb
IFikN3PjMc7TtdaeBM7Ju8WEZ/2ZX89GxbsWWI4zUIyCHcUC3zjZdTO12J1w8W3THMmf8hVXOX+y
b1ZvsH/A0DIQwAYjbYFSyLueewoNsG4r42PmNIE916XbIZfm3wwJss1NwryR8RwvA/HNBC3wDYrA
6OxFrXKToU7WKKxkYYUctlr9CFDLhxRK20xagehnYnz2RzYjox9GNdPX8la50gJ9UIiKGgJO+pCQ
f+oQml+53P6XvZ0lgdf3pbAYdsjL1iAwfCwecbmQlC91+pTl/PwWakyNrU6l7XdsDdgErIocvcNm
IBjG3RcjsbzF/2pL2yjkQq4UusVGtxVayUnEiMJC+H9TQVDbpbvDiYmN2Fox81Zbm9p6i/wlj514
0fhScE/z8dW7Xy8uytPUIWf2OiuZOLZU9Dwp9TmPaearr5SBzpDjOQD7JjanZWvH7KWTpCqy4SBO
VJ+Hv4AkkOSPOfufkD6Y2GwkqQdv2qvFQ25xmclYx34VbKXBk7vaKiY0pCqKP75th2pn9ha45grK
1ntW8JcsW3r9C2zlFR3h4PlbBDwN3urCKrS8YsmC5zpLjH6gUjzQnptkSV3exj+6T3EMxFaZNS0H
8344qz5NpQWgNO4TNtfq3WeJhR46iiCPFdsZFMjqO02q4HVGno/xp2E5SH6S3f8Fr7TgyIVIoW+t
+RvGCQimU0I/+jEfptQISYaYoAx7KyanwhncUhzxKCq/M7prPXbA6aaUzW40UuhSH0zddUjPqDfn
s1EaUguuMXsenYKJjur2Hd4wtQo9PjmKhlRPHJDVZ+AhtI2boJay5c7LnjrcOYhjLnZTcelFfwA7
9+q75Ib36u0LF6e8Fkz2xAJrGIhbgItSawKoJYeCOvX89amFSOE2dBpL9PXQOHIcrJalDZqAH6wS
oXpzUmWmib6p7yJEZ5viYS5vgqj2xiUCh66iSwWiquiR0NPw27sGe+XSSrh5s9t9RfsrYvtmic0H
BPID4ZZyGDkHWOqtV4gwpmCh/LYQwMmyEs6F49JcTVpfxhC4OBg0MowYLiqPRQET2oyeQWnfqJYG
G+6sGxUOFJhIwr1OI84AguKl828e6l7KDfhMIFMz2jtpebkooGIdHh4G4Cxd2DDl0BURD6CBtVkJ
4hfYRuhzaCFLmYlZyjoGnhunCZcQtwQflu9JAiBrBCcSRzIDSnNoPVRTUdkZpZ539iVm2H0+Myxt
SsEQ3KjNE0unxSNczaeMF2Y0HKvUCltriqD7pAzobioqrTGvaATR10hpdxklVd5phnNpViNyLDPM
IJvN5R9ZnmprkSARU6w3PZl9OGTY/2XcpDm8e1BPQ8i1fdUHMaRRXkZk21PNby3EfNPdwf0W9ayj
Lfh9wn5WG0NczE7HZ0GaqR2i4PZrmZt1uEsggl41c4v4No/5jn/1KcN9grAezKI+0F+eKtMFr5vj
H54lJ0l5/g74PuZ3Ig1KRqzTjEwLfz/dPVS/Xj1p1ZjCm3p9gC/Cyzvjonabvi2vrTLuketAFbgM
xcOl1FzEee3XwQQf4elOzP7opO4mN76E4pg2PwIywb9x8pYL/AWBPXg/7rcpxPdSt9knR3WRWPHL
NvLSRX3EEXcepUdgqEqB+uiNfUnSisbhrRm3pJJxZHLoPauegftIB//zLCD14inmqxVIfIHG0G90
XdqtEdrUT8STM3+oPgemOxZ7hf1KrMIl/yRkdsyZr7jJv7i6CaRNiLldctjq5aoam4nfpP96EazG
yKkduwLN+gIq3GXPP3vquwMkqoTEZSqMAsxR2NYZbhiSFyYfJuju5+ZoJtHfePJpdCNmGLr/Ij8p
a6ETv2Txif1FsEP6S1IHfOYpzaU3RhPPCHzL1jIjR4nut1VADRvJOiDhswXtKpX+vy2ap6fjUVQJ
QeV8axIb09e8H+rUjcvlXhKxaCizEbvdurFjzcjaR9DZFYsTNG0W0ugmKZkj7nWix5Uk1cRMA8d8
UfyPb3Pj/IG2vYbXPK9EqgYcq49Nz7Ii7qjKZdF2YzRXyyqw5WT+SjnD7BjslE4lUuf8IOyt3b3D
zsby3D36u2fCFkWxveOQcWx0F0+tPGqGW7BiiRaLp7roZiqV+xrgahcOOS591O4UY8Y5pWp9qjrw
l2+YiDlv6lan4GRidyAEIv7pJ2h37v4fv/bkDP6wxg6H0xitI7FOvJWNyo82JLQYg2awlsRyQGUX
h4mQggMVwhdZHdNwNl2Gky4Cc4w8cx0HphicgCP3idqJm6sOneI/+acl5BX5Na7YQQOe6njfODR8
haINeVX9JoDKp1dm99SApi8ZdVcYTuYryLLBqpurOlzqRcOGcQhzof2pboKPXNJdS91ZJAS91o3Y
FqEEXnTdBvDpo1rqwVcs03pw6lLGQ+2fBssOTmZznMybgnBoEvja00bghSt/8O6KhEXu+ND1SYtu
uGp2fjj6bHePI5Xueo0bbTyWM/uDG6lpOdZtiOMA2EVmHsw6ONYaFL0Uncaza/zpiHm93b8eRWzo
iGTxO4m0MZ0odCEe9ULLPPspkcqAEqFJVci6acAPE2qnOMDPXfnq4nP7YCkMjqTQ49sl9a+Aqt40
28sg2sPKkixH/EY4GidEqBqMuV/iXLam1Lc4qpYqezU8UVsUR9LcxMh7h7IX1j6cIP0bh6sghKMF
IHBqktURuijI8hCxbjRGCvQAMZdHdbnqKEg9N9T8gQWz3vvuGJxryQinwFcpIPQoMUAAhjOFErUS
bFtcO8LKyBpOYeMiN9GohGic28b/Y5GejBduwONrPjSprkhWolYUgfyqDG7kDYja+nUuSDtOMeNV
eShUm82d1tB4mnYKWWB5D0LPJkXZhfqqWqS8EPcfv/vaOkdSn70Z73j3C1xkfaE86lXndBHajaZR
Msep713kRwUlnjgiiw9VUd5eiyTXKXqvyG4mBItG9HOfYZW1DhT51pTWdqoQpusMrqxZgcu0dD1F
HWAxIHuYoXGvH7tGQLYfkKklV2Y1kSGXywftiLGCFM7IK9QZiYLdWO/PudUryeI6E8VlTMR56gd7
/QzY+YzzlOzaZhK9jZqGeu/2wvGGSXxStnB0ZoeCRp536DjEIhcZVpveZiljhBSgnGGQLuv0EH3O
vQjrzoVFuDI2zDoly3JBEUyQXHzflCwIsiXDqDPvPYWWKPlLwrmbMWyHTCkpuVSSSP3rVzSsu0tE
rk6w1DXqB/Faw7hS7oYPx575k/Rf4FJAI5VsCcjvsjrpe+5SYGMK+PgQ4FbseqBVk3e/4ifbGqt7
lF/fc2lYABlLOMkTmr0b7fMqz3Q7HgwMMlsoXo69Q03X+INvfiCAHwrZwBVFARCCCG7SYG0Kpklu
FKQJV9H+7CzJV9OWyIgJTPPQ0IrbU1WsiRBgCWWwFisXPFFslxDFzgdPkfMYpo/UAz7QaK1xLog+
seTIXeUoLb58C1BZ3Gsm83sn23RXJvxEshuBF5ZBntwuFIZBPTNERHarK+fTwJ/jgnujKzFEVp4h
tWcihRxSoHcPUw4uNuHHurTilYTpuWjqa1/qqI2/KMQVNnB2TK5i1xSc/yvs3dApeUZSpc5QJDXB
HYcrbZTvRo9bA9rsRAQ9LHuS9zxNIitmCq6l+XY3nI7bJyvyUW34WzjhfH1BkXM9POlkG75fznp+
dw+Lk0fKDQVlC5KEI8nqPi+tDf2cBR1jssJuXbjd9o3NLBqE6AiYkJ/6N9C6+euXaJGtdFATHjLC
9K87UqQCehN+ssXa2qnDWPqtM7FJDs3o02cdcFO93SlaK/dv8rBRrTG4tKrmZ6wz7OGvZToA154u
jl9jzcGYWFF8N9VN4tT42E2jiVDLKDQnwfHdvmjAB+bFdila0jARFOeTpGW0WG86W/o220o/RZr6
/pJJOpbLnycykUvK7RsAgEZrqlAw+ycWREEMx7PktC8LWgVGoOMnaFHWLu3AFNiH7fZ8Dv4k3F8S
u5QMH770aNPYZyZY0uv4hZXyzP37cErUnYQ0kwTtTMPoQowBa+HhZonAgOmeUwWS2dlYZDLVZf1A
IL/lYlNNBd4rRwT7fPs29I9/j7Jap2/zGFPl7PgNOG852gkLB6Ru6sLH1UjGu0naX5LMZEA4OjDQ
BrA2okUitU29Q3pQM7vmP80kUggIxDnpzLKW4Ub3/gvWOlqT1m1x1VAhRwJ+hMTutyKF3TmrRaHu
YTOCZ3A8F052tzUelMOp7vr6yRXUSFLh6qyp3xpNwsTxbnlbZuGeYoGGxQ6UXdc1ujacAUR3+SGv
J4kqorQumO69TCQ8T/I4ArZtKtx0xOCQuzQkEs6+4DDkH2m5wPMY0ftF9i4YzFagBX3DU3V6379N
0aSnjxMzjqLbjQNgc503OU1xZGMS7urRjkhpt8zrxVGiwmlDBUeUNr5uotZH0vK5wP41KSnQ5IIs
Zf8NsfVqFTPx1BKnfgSkp5VxZOu/hUJrWXGy7lRCzCepMba+FbonXa7YTNyJkXltd1BhPhANcCD2
uNeMtx5Tt1LMHx2S1bThvYoxVOWtzXa8mjBdMAUSK+8p8QDAXhqNz/RGpC6JQs6FoNuwbFLaoEwb
4Kaof8ATSpbRBQ5TgZXHUrW4GLgNVFmMvMnu4Q/1jug6zbYPsTUZ59YzUxTgPBI9dSFZDHPujpBk
GWmuKdlcTFvVYnnJ9Hn1QouZE0nBsh41qFAtsvzGkX6dAyrU33PIRp2EYfrIr/KVTFcri2kjPvKm
Lbx1GGmNuCYKObATqGsPJ6pt4zpDBP6AZNYLZHevOi9o1vfqtMe3Hb0D9WOP61jYOo7KRE+zfVAq
zUznli0b3CYwWjOwa5hL2RXQyQni59yvlJsIZvjarkyzUxJ20WGo/YIlTmaQyf0/3qMdfRC9Znit
0g10uWkhtJ34f4KrhOkfIbR/zCbZkEJt0AiK6HOc9vLew2lKddFmJ+c3dl2DSxJ0n/6Y8pabO3P5
psZuEROveQa1m11vegZzmntDSZRhequfHN12F0UQOSVZ1+sKj47+VJzYsIqRXrjoeIfTEPK1aGSp
swt7VM/TjloF50j8dl939K3W56ERaA76vyg0CRMeVgIJK8caPkBVneEmIdjiKR4Nl0CA37pZP+z0
KWbIyrRXj9NmEu61D9dlvqGbWsinnAYvrszoxufy4CBuF5fN1ZevkcbOryAYmK2w30XFOdaG5gzo
LCGfBQfRENMPQ/Smq0MSZ4y1hR+nelXTPKgGHefzXm52WF8O+hTcA1f/GGQsQMWUSUL1C1hVtWIo
P3VjQEpKUjuulPHvSb0QemWUJ85uCXKMj6iO9e1iz5XtAEk1ZxxiUfP2gZP25Bfcw+hnqH+6zL2Q
wIF8pONmYF9/RRpD4RlZFkQfZMb+/qYd1CIYvH3X2HpjJdlIS/G+EJ/6YN2SfXwCd4HT+ebuRyqN
D/F3/qEdRXWREGTmsQFtHnj0MRLpiMTeakhXjPG1ednztLfCrTeu2tTVx+nvuKm+2yIDYdUoN/ei
gS7S8dyCdaF+YsuxiunfCWId1zDvmdW5uaugC2eKNLy1NWKEQTsz7yL4VP2lzZLZAIs6fpPCt7F6
Ycfpx8roXZ9zS+d1ciU8MZXeCFg9t2/B53NcOmoXZDb3eVb1rYZPwlm/EEih86+ZVDgx3RWKCFXn
wgC85HgBrtJ2nQnug47l4vZlfRl8N6mYNHKkVjHlZpz7hSNhbrJXXxE/D+EeQaIgRgRMxtoQJ3iD
RSof7E1c2OYIxAC8erbETjGjk+ng0JpZ7W6j/1g2iCUCMWaodlXDnubYckIJky7zTczF8bDRbp60
CAAuZAgfpny9zgCITT6tlczz06WBIyZsSa+clrzN2aUaiauaOIcn24DOeHOCr3abY/ealdgbp8MR
wGYRMOH7Hd0xdVbKEdKqmrxhtY8NaGQ5m6YN8PN5FVC594O3gVUQDse/BZW58olYF8AA2i/89VAr
4JqVGt5Zn4Sy7Yqv33EI0+jPcLO9YyDYyFmuJEs+KUKOMZZdxLZ4dAdwtblBN++3ugoq/3i3wcVf
NXyQgsXPQkFINIgDO6IiBXLKf4Fnsx6azNHUJ2kW76eHQ0Px1kVByAdQZR90hhZ9hu9wH3zY6KS5
+dxEaG4u3HCyZBMfllgw450mKBGNEwvPaow/EPtBqmLHlNSiD+8BHEyoqzPrZEecK2cbLGm6nDnx
pcSFNJKv/ft4aH7pAupPl8XU1HU83gDjrKmJUiadSgiy6cgXI8Onc3QrCRDTcF0hAT4UvnoT9zfj
ayxp9Dh6n1kwhBDlGVlHb22xrJ9jbR2hSJAZpSM4/QmVpmGlPVOyGQPylpblUJLjOlcMkBUOIP0X
1frx6xlOMyZNkzHViPYI/wllfk0ZiSdCJ81PJ9iAeC570xIbKrBiZiK+3+ETNei81is2hboHljP/
dHm4Qqf8lOqCLGsol9sQcEeiyRx+5oxu331taZ7TceTyPErWnq7EZTv5iblvGQ579SN0JI7Nrgh8
QW19RX5syxKlrMcAiV9b6ZJmtDMZLc5QmMuwxWZsEPzBsaS1B1xq1ONl4h/zkfawcEr5VjFe6bR1
8w2pOWjk22E6xSqmuKjr1dB46epV5pVzVkzuTSbaCFt5tAPalH1CGaHwZGDtHUorDo+w4U4NwxXM
Jc72tEyRPukRbUhmLPIaTKE9lul6dl6ENDbgO5p0HtYPunq4N42coSwf39JdzdYJpDz8StbclJFA
/KtxN1YNoa7KYJBTDl9uAd71bIZJDbXjtonj54U1vJoxt8Kj8UDImrsoJY7M6W8+SOIJYZqU8Teq
YrYnEqWePyMIiOggIFr37ILJdhE3CM1uy4IohTM7P/luIrj6tzwjdwtB0M0GWcD+LQ9wtC4rnhph
Ivgt4F0DauDVPd74PL57khN8bb/BQXnMWkerGPVIdcj2ue3Vk1rQu8NuQvHF27oFIOTD7HLAAnEs
LkEuWKsOCKhbENVEyOAR2Tkd0EpZyv66edTkvQOGjVoncyO0G+8nTJjB5rYfFLkpT9ZBktQgvFiL
6QetSGUlepTFmFvajOm0Pd8tz0NBAjz20A3uDMWWs0S5PpIo/24eu30GgWd3Rp7x6aYNBuuA8oh6
pTYsRHYTxIOlDAzhPwiF4SEijZYONMO82mxkbimsRXjdObEhGFMUZTQywaN4S2dORqFjjy8pMNxO
/qyRThvkdNP7k7IoVMtLO/kjDUtD5JGoMyI9dGwvD3f93hivNtthJ+wVFiqWAj7IgPHzHZCZtOFl
AH1K3u30e5AMkYGTWddoHImeUKjXJG5FKscC8uulPDW6FRLBqe/ZcpRVEoKSuCVwi3+CHqapyinL
1cIMPAAeCc0zNMXWw4XRkNtTvTtLBpqdstJgx7XDVSxhs3vKWFIoV/beCOd75qoG+s/o6zrn+9+z
JRhGnhU20FgwYDcFDfqNXuRUghzijY8EQ04PMOmZvG/829aCNkklWCNZa93YMwfEABgo92MLT9Qd
goR4kqLVVmMtiX6xg4Z+T7arfUhE6TIg0kxfhNiCX31mCP5/geMND1+M0JO/93b6usoGEtLMjPcL
fZJUwk54bVclA5s15fUTAuGKFoCJbzNcbQQ3BHIjVAMR0j/UCRlKvmoun/TMlKLl667GYYrxb8aq
6rU2m/N5d04pFs6ywYQV7dJcEoyU7QMFd8k2/vQrYHqYZWi+giNNLng/pZWgXmsqsPSNK4XU3OlV
39dBV8+Uo9hN4xLWgb8aCuBMBCPoIWd9uUJw2hBzlrkFXr5EGyeD0ZpiAiAeO6Bb2qmvIRePlWq6
de5rYbCTTVvBXeSEkEgGys/p03cxFtubHdVRovjpaQ81rBVje37P8X0gBdLGS4xA/4rHTLRXDHUB
1N6eteqeUvlNGES+dLet1vy+HajmmRnwhEkuMCOmgwifcS685OasXHVdk8+rXGalkJrUESKNT5K8
KNYICVF2mQ669T5WwK3ZweYxKAPPCLrok4ywKjDwYQxVQNSNvSInn4W8NToFSxUjNL9g1e1Efcfz
yY85ov+0IJ4MgV/OQGVA5rX+mUR2NT25HYxh7W0vEovCuoMXamg/UOBKhHwUhmKzxRHYhcFFIrv9
1DGOnWK43KYb+3oUzHFbwMgxoj7sDy5Q9duJ/Cm/NzxERqwULt3+JfzaP/E5i0FyoT25rX7NG2UG
Wt1SV4ZqegFMi75Ah2NUEt0Ro1zbbNYBV+o61EW3hdo8BKWPOjkm5/3Cg3iyaya3HoU3XfE3k0nN
utALo4O//yyuYtNXNCkGj625WGnVHo8iJb68p+Am3vR17G2QGN8U9W8f5lS22WrtVZdRH0wulnmw
4oVSh4wCUwYG0rCbOjQtDZQBp7XCnR9j2JG+tS2ewcuUjr9rKZ4lD/LrYDYOCU9BxI7/EoDJmYow
nAfvdIoeC7lpBLjkInoXPoFEoPFqfd0VgBmx3Qs82AAF9DF0fMYg9fP50UPI+m+rW4Vfh/CLyo93
q6G7/3NMRJ2vpgzTdcRh1hHH/3EJPz186TZaEZjNGQ0nRTdZiY+jIwilKiJRvoaw1eoPMM8IRDx2
g4XV5DV9J1f5slVU+4UeMPRmpE1KntkYVNN3wUhCalfRQQQWmoB+4JsU7QvRPtdqZAOHu13K3frY
/K/bjkKPLJjpEzjaFYEfQ6qNZWp1K4V7qWD9Irnec87E5bWnryWEER+V0AYxFJRtNUlHN8Luhp4R
RGVFBdYagLBs3HiwZL2RwJKjGSqcElBQZq9rZ5paKiVFq+5STH4yTvrNtBrrX5jblr7UnuNq4dTq
pNkbTrWyaiOTTuSMyDTNQr89S+X9kAsOn1i1t/sToK/LrbRxDRKYBKQCYfB/lminvZ2/bzEXsNzt
B+ZuAKLGlIzAd2OgNOiBUuhT8pz74wQlvhecc6DdVFXdzot4D2v1iTjp4w7npu37xTcGMJPfUoW7
QzSViZl4DbcwO8hQ+HrxFloXsNF1En3xQud60vNiPxhpaL3HjTk96iuH8BPzxAl+JNVI5snZ2xXM
JL4A0P+nIwRRUqDgSNyfD7/o80l4jtmpgnjmI7IEpDWqCbZ8rkwX3Z2C9XbTa3OT9v8HUnwVJ6Uq
N3KMjKQULSnE9cEyNT7fhrnhVrLmcTdGfXNbrb+dW5+TKcwdD4DjDmLuR42okLNJKFltWCWCFnPx
VbQMMqZLKdEmoiptvvrD8NM+HneQTfiB7paTd8GKbSnNOBpVCTcK9jNFGcxDN/4GFCIwaEh/CR/E
IXEPv3X3R/6yoU/4cCC6n4q1L1wTUkBDbC2kkb+yS05wF2/jbPYj3J8svmU3iHbmbQFhod69XS6f
2adZy7ZM3MEVt6UcTSN3fovVHp9iJSK3GWOraQjWZBapvpwgnxr7/VrJB3aUMXBrH3Jb6hYguYek
ocabVWD6PpPuCuvTvJrvN7i0YOqjvYDi/jAqToZQZ3KghI8w+PgXY650DjQpI6yby44tbcWn464G
Jcxgj/9N2piPXxlt7Lbil+fGBAsij9vhp7KByoPa9aGU/Y2G/VHquokkNRa5DHZw8AI4Q5Ur/n1g
2++io3ew4D0W1i7VA2poC6N5ry/22zOvo01Q4PDlztzIPyBZFaOLMlCStLdh45+e5IC0MAYxBHNs
D52Kdc9+zNW5ejpKSd1xJi+I5pgxe1zZbge8GWGgpnHGRB7LOyK3smRnAatFHCMYof+EKp0e/L7+
+TarBj0KwiauBAS58dK5cdTfIfT/5GnTcybDbUrT/yygEf+6gXLNIPA/aqsrSaxJk1cc6NwblKH0
Et17CoWtB79TyuwOzZ6goNQuGVSOs5TPDQFa4E84DGCLIeUFeslA0lqdWxxthbvsY7l8RGz2J7Yt
8LLAcTl9/507tfb5YR86F5nyrEzXLogQX1hR45tx8C27G/6z1uNny/eJ2YWpmfYlwRPNAEuXKlCr
oUsYWIjVOo3/8YLUc/bfclhbghoV1jGUBmkj+vkR62cziM9pYWSafUy/8N/gzlmiJyjohZiw3qY6
4E6FExZbjsQyvksYRq8/xtn3OC6DdrUqs+l7VZ6m4mhiBbq6A2bmXWy4Ik/X0ZvC+Dr5TiIUhx8d
taFThGz52XoGhfBkfVnS1ifC8xFytaRp6adlRb/hZOwePk4Paobqxidzu+48uqCDun5cDF5b53v2
aL1cZ2tEP3yxB5spaZfA1b12rKNyTe1QRS7QQMRTN7cP18LF2cCkpx/Hdu8oRccuYW41dfpCUQvL
uDqTzcoRdotSP7njNfgMQFafyd+a3vM/ey3ADcI7H7di08T4999rKZDKOROPIqPG5TRXMTdtFyvb
gKSu0ftyta0Q8N0TlBe7M6CUo/C8tMw8LawQkK7gO57XlC91vVS+gNr8vhlzahMZnF1Kmdpp8mZo
3piAip79K4A1zljACWqFMmTJdyowOq0Md7bwcV51w5CsUUj4PGWosKdHIDaU+EeVpEQRX5LZnkBm
n0zIbGxWY/utq+nY9jdClvqHVEG5bo1n2GkOwwGyl1E82i1zsUl8GpT9Azk0LjnsyjFIip6f37sS
0Z9tJkqDaWAWKMZtqkpy+zrwCN9suxp/iFoDcPMwj4KJtcsFkrMsWeTgmQeAVP6NDLt3eqDdbywy
X0PPwxxPP38G02uwCp0PFDehlvxrQrt1Ufq0KJkVeGvNwxH/lsOyh/8EAopfGAkWYjZ0boW8COaK
z2E2ArgPYnRekHnA4CxV82UnmyZ8Ww6Jy+6B2NcyrhKo1PjLimjR2QNBAz65bUrv3nkN1OtElMh3
iMpzc9yqjiNbxTX29H+Fgml2vvKZM34SKQ6HQXDHqyAmT6k3WGBtv1QALfT7lbXiVgt7oWpL68sC
j2cGMUNodt2yrL93Y4tC+mu88Q5oD4IDuSlxriv5mbcoBnPJrYpBSrDbYlDZTj4iIAXHEPGwytE4
ibbaC6fm46w+cmKlU+5t4j2jRb14+5OfH70uzC3QZKJr9DyWKxeDqluOLAUHfPTSkVNFLpBeX95K
j6Ee9S22CLRNR3RcBBnis/2/GAevPJQU7lFScC/cbz3Wh0BBZPrW2+IPcmIF/xbigrzXam13DXKp
fZPHRlcUumpbj1Ywcjo8xzs2451ACNEiPVwHSUdxhgHSiWA/vhgSYyJd8GZftErRD8E+RqLGZ7lP
r/6uc8fdmg6UYRi2nPNMJh/END6mCemS9XLy4v/h5ezLvbcytd+TEnisC4CuPaPdAyLWs4STpyqo
uzdC+s/y3Ikg3qwe5v1SZzYHeT1pllnxnVftlxwW/rGaEuyYKXwuffyTFeFPvHjCtcJ6JUgI8erN
bb02Cw6J4qG7pSNGo7neZ0ZYkfAQ26fF5AtvYMiFBpqNaOXIEnpaFstoBkkq9WX9GaQFobeFOJr7
dZ3leMtt5rP/VRBEmn0oaSJIb9iOKCmkEvYoMxxtEzw3qv60YO2A/K1oZdZrQXANapzp5Sdk8vLf
vfQFw4wZ2k6Ct3BFDfe1+cjuCSdVXuhx3yeRwAPzDzoB3yUXytT12OcqePbxg2fLkPndi0amWMvh
YOAgC9nurX5CQtF35HpKqK/LaqiRZhtnis8SMSrwRgkGJPInLwxIC8mkD4pmWtdqOvPfSpMG+8o5
4/zPA3msUSJbSuKY2OcOOqU38iYyX09EHpJ/1Xr6nskzqdXbSTF9T4Kc8oM/HZHTQAUcNBGQwu5/
Imvy3TVbnvPa4n5yc63U3SV7qNnXFEbU8gdQFHzyvVhsVAWd07Z1mnuHFNmGzNQyLbKGMUjxqM6n
K4rr40U3Zwgsik+kpnRo6YJWaZUF37XGLj00R00x9X3JXCt9KRSxSdzYQlqIGdbIAq58EemXGEqv
R7N6PIHzUq9kU4Xz9ijfi4mQ8L5A8kvElRw3u16HD5rzJlIDdV13Z72JAEs4cjPZW3ARquYGSj3v
aU4nI8l8oizgJHBfl4ziKHTJHGVpwd7RXqXim4IqzqBOxTdCbtBUVG7rZg1nKKzogq7E7VtGTs7l
ruZFUqy43n5WvkYM7C3D+eZyPCIsrHbiqPjGVdoy59faU9ZRycwijPWKxo9PSoHmKWs0eexDsAcP
tTuftGCSqdkGixtGk7ET0etXvCxDnl6V82O9MB0iAtp73Dmy1Vlj83NRtpqiupRkqUS76j94OCuo
LftsQklpf/FYyCblrVDHZb+T5YBXyEb0SNfgeCUEbIRyzYDdSpMhFx7X7EWg3TRjmzWn7bek8TBm
5atqzzMLwdGpDAT+2TAs3IaXk+LpuYJlw00CzcassiIoSAD2ucRXQ5B9uE0nFZgbeoUmafe3sCDe
5V0Bt4/SK0+RL8lgCK/WOoLc9lwVsCqZ+uCjQCOrHRoXfcJERITLk3W/pIBI7+1cQhCjOf3OrrY3
6y4HpKMwPgvRfK8Tz09j5ZHn1aHhj7KLB8l5+WVyMOa2q3u9wEYjN1cYMJ02wkqmNCr72zjCSCT3
UjICNXY6xABSRrJ+fubU6I4rQgGwuA/N7LLZZrIc2Ddu+cpismhEILVD6l0OqjLRQE20Q4nyqOJ0
4etC7q8Uu09E/QyeCSgngQ/++3milHIicTh3dFpRK0i0wXWinMwYvHauIkR3JGdgs+ZTUx8S93HH
TFbUNIrYNTeM2Dzr18jk4MaHlcS5s7S7+IPZMt9rAMlP04+YWcjMPvQxF7OjCXEG5CVSQAGwq+1/
gU4e3ztNykqKLkrC5xb1QGwn2IgwWg1fzfI0YGJVVeem7MqTEVQ/p/utNV9yC2dTU1hK1SPQhh2P
3E3J328hfDBWsPouD6S06tyL10axXGcMHLbjYpHziXWOROtfqqa1M4MNAz3X0ZdPxEadmQXEOW2e
7WVqRelDs0b2bUkAl1zgURSMNCX9Wf5RXBfs67lLkhiXGp4i29ZqKeT5Ff1eQPQ2YmDPEKPFiE7k
jNvSQbyn2w1NZ6kIAlvj97WD6tEwbe42Ttck3Sw8X1M6eelA4PftexLnZpFBz4j5w0GLL1jJzbaN
PtcNy3ZExjlq3nUFQMbkw9j+WQuwOds2qg4RFcL+LBzlRS/pplHWon/ikdIj8cKMC/24EMJJf8e7
N3gVQN022p7z1RPWHG72F4Tdcwm2Hg8keG6e33y0GqSgBF+Oyn5MFh4B+2BAkG5Vlo/Gc+l5Ok9e
FHFIR0WF0J8iTsTdg/LrhhqQh25c1mWZLCnPZF85MmhuNBjjHtsPEfp+Qpo8o1lOJX6pesRzyI7f
VKC0OfDyLR82uL5+lAnc0+OYyERxquC9iiTWhsipXA5WuuxR7NBQw3OjY0a0QzZwdUP3cliCCKdU
oBvSeuYfGkS/2h93vIyix+K0LK+HLnyraYBRw971b5Ve/eNXNIBBgo1wIHE+0d4oQWH5Lzl1zeNz
bO+wNFJTjOD3eqSCL9jw65wSqRVQiUPPFsWgEe4SxcXWRCB6jPc0Ly3ltD+1HaA3QX+Bxg/NvBqU
g0edTFrHAisgDs2E7M5KIVDIZfJSCnMmHQCTU8h0E4+pQOomwL9DVMHVzgiv9BSYdlw8ILNV4xFd
fe4bpFXVtDFwIajXooesr8ZDTUL5dH5Ja/c560CnY4ltnszPf2Axk8mF4N6tJtCq2w7USSaFT+q8
kCu3NyTXUlinD+P176tG/LPkpoE/k2Q+EOL+GHgpZtFjb0/zkF9vHSJ2rcrJTWb8gYx/kxTs6hnh
4tsGbXmvE1DLFdYeJ1hbO+oz2HcdObI+yHFIU7wbTQbWvTIN+Ekdedj1P1nBw/2s03wrAUgAtYqY
9VD6M47YPiP/vyGGEt8xvJjiZ7O8ogl/xKsQveSeVQj9dv02Y1PNvWWj55Oho2DDyproefJwHyRz
GsZt6qDnZZI4lERbf5ywPC6G9gHtmVjHEYlniwwvlQum6NIo7h6mT1XpnPAtlSX+qiF282KUZNhs
ieAEP0IS3NxVKlVSDDe/uVMhpY+lb+56Ic3Y+pQdXBggrVOG2JUiLUq5m4UxXzuCfLT0iSX4fqEw
ZakVh6JHaVX2pxiPaM/cE1pMM8mgDHowQWQBMY/ITQl2GjnNPGKSJTYXpZJeV4lCZQEYZ+pfeHWf
9pM+w1wj/DrerZJ6W70F1bf9RdwQaYyrbTUj/Eg5dgRDwRIJygZNymcq0VmVLe+IKvF0c4Dh7vwM
rseK2AzG+muXnxNDjeBxSd+GR6O72t3EWuWrOZRUeH7nIM8mSjqtW92WcfLqwUM5p11NNe0JJj/C
32aD/juO/AuoQPPzFlM7fzXoZVVKvzgRzePSStKuzVGZ+UXwZTWOYY0wx2EaKExbX3lgqRGKnx5C
LI+Vlb/IuVyYjcruCTzam72NKtTqYH1noax7r56BNQMuQBqiwDu8pOTGZCaziSmym7Cy/BVbRG0N
eGJ5l8wHaCm0XdkbZ5HYroq0wl+MdywvP9RHxcgCM17Es1wpPCAbilSTnD8pdO2CFjN2l4Cz/uue
9hLqwnDeXHpDWeTyAdrkn+G5fplgpaqE7vDqpBJMFD0vwJVo0groK1mYLpXTqKWw0xEHnBTodG+j
OdoCaVJRJJKeuv2Bbkfmp9dMYi3Au7g+O2gLFgAG+RPuUfMmD2Y40pRCxnMNAfck5T4LeCgsTQGD
gItM7MUo/LvrSzqulLYLrU85gmzc468frF0EYdApViUq3u9bL5lzKdk4N0zEzAkRbAHzk055SBFT
Tp+gZ/KV1hYX1MOOaOigS1CbFPp94oQ7Th1UakK5XJfpBq3uCHH+jwWKTg2fjIzHbzAlGDREPFwl
s3PVpgSQt3N3SABMu+ltpyJbxV/PvFMG2CJKi2VHaYJgAp3EuVxy69s8/k/NUa+SiFTGrEqFU6ly
Lh7c4JDjwQ2N3E4+FofT8Gs/gUU6VFP5WZ+cDmNBIwCiKfYCTU9cUq7k3WHUZANDu4ZhEcIOMoA+
YIu+UREJE5IuUyoMaWM/CoL0ueGIltg3BeTdTHkTW5Ku+icwEWPmIIQCHFIUqOHevUfbqoKV3SbT
l5HGF9wVr8dt6zRshmHNAW+LEGhUVyFh603DF9P0Yf4lt9HKTw/ch0W0kwGxyFNQuzE0t7gP6kML
AewhM0W9+3p+HvPR/cyZP0rgIjiTjl0quG4//caQMcSsn1Fb6ZuPIxN8oiigWqym5CJ/ocbP/ycN
6HXOXs270AyhtHo+r3KjhfhIf0bpMmF2jehS3M3NkxaUNZobJ5ya2WG0O1vK9SeYbBFIlSYG3fRN
UUnEZoR2+3JfZRUMLMCGYZipspKoGsaJ5lioLloi5p71UO/r/N2caneojHSxDyUInwoy02drB0/o
rMeMPxzfg1SZPantKZzGaTONCMj12Nr/RsyDJReGmceWHXbbeKNk+22xg2Aw+8ek5be6/zCfqN5A
9NYzAPH9nVbYVtTKHt3mGTD0gFQDnPC61q6i4I77Iu59t38rXVwhvqeSan+rIHSPLAYVJBRW+TvV
hiSYU1QDGTJXAn/FLJfFofBk94ymmDbVCNj2gsfblR8MUDa8xcCkQM+1G6K+l2BtGSwKhmRY6OmD
xlmpNFCryRzy9Ovxn+j6f/EUdVmwtKPVhtEfKeqvsLqgVUMqTxdewtLtXyXIIt3oj+HXP44TDpT9
MAvn4BvzmmvLgjX1g4MPsyotCgAE+6UPyxh1F9ixyz8KRjp9ngQufM8W0bpObpqIDrt+2KoSjol9
kRTzwitNxhVSGzCkXhI2sGwyYDIvAZBmoBpG1lMteIEJ392RnV04OlT7L7ufQo4j8TnEkHGg9FrW
x3esAQTVoRg6KClWhyWsxY6UiWGau9xjys6cSwl9GQFt+wSveYoObXsDQX4Op4MT1i3As8M/Pacm
maEHPgWtPGYVvwDpb1szGR424FI+LoNbBY/TXw2Rbd4hg6Y2tU8+AFf7LHDeMyroUtCSi9uY8OW+
TIUUCmmOmFdam0VFsgt7bxoQc/A1RAq5iDk8WdtJXst9aQAixNGM4pV8+WmbMxPdkS4g83Fc35CN
TzqSIlGx0CtaaNr3wjFdpHr7N0IIl88JzK52Qr4HuLqwbLc9pWA8s7M95HzZzd8qCXyyM8y4SC9V
yTXNRWYNU7o9QCK8k4ACRlC1F1Jxy/1uO2pxt9LDdYclIMuXQ5EFk/f6zLs3yo66rhutZ9nZK33T
0+fWotFFq6LFTf14TzeshAyqjKOpySxPIIzf8xm6sKJeVfox1ublFdYLk1q0rnHeCkpKG6umZFxn
v1xbrLRt8EHMDA1AjcefHcSAClZrTxeBt0rqMKbzyng1DiqWh0/F7rjQ/WunUXJS3FSsr6ewOoSw
+avRLuX8tIJPuvhuCqy6Ps5smItUGO9YiKqQhUwmaYyKyslmCXmOhSE91yFjPW584lw4CjQq2G8t
wMDbWhnrcNVsN/8H3iF8ObW3vspIokbpxPCQ7DulrhPhZ6UMZhSIzCI5WbZs1oflAnr8iUc8NvI4
pogTkv0vtPdMPS2aEOgFZjRke+cMRb+EMXvqLurEBEM9nGZOSrqoR4NzvrvVKrFEAbHQ/KczL3vc
DUvXxUVIXDNmmf2uv4kT/DxY1A3k1uHM4pQurjyDM/OpNpx1XOvUmueah9/nPkOCVIA447D8Z4bO
hjAhRLdxuVO5T3N1FjMYbzZLR2yC3Dz/ABJaZBNBqc6X5uSbkBA56JNRsLiarkrmCrExCmjgYoao
Xa/BlXLTRU0qhGS6/mCaP9U2913WX74oCf43l1STxJ7q+ighj+8Y7ZbDM3wI/cFyMce+jYglFL98
grJvOiEHjF9K2bkq1tDlDgntcHVb/EgiV2xePBLGehykYmDllsOK4+uOUOtkuhVM9iRuxw7P/i8b
Rv58qgrhOBFeLheUh8iT7oXrd/DbkqINcGSnh0MCoDb+C1csH1kxVzf0M0alAYaW1AMwgfvUsyqp
poSTgnWoP7pS77Ix0jyL8CBvdheinwD2o99SGJOICOxUNXyatz8h2RNlHSdeWEcAdzGUwIh8hOb2
FcYwI87rMfWXgq56aY6eofh5yNgAKJKvWyBtEzBIe5c/yoc1vsx4WRIAYClX0x6PE/k4RDEEJCW2
V3LOazX2rZIvxbXVv6HQTBBICainTvEK0u8BFK6PwrVq9ZAK+ClrMfxYppWWy7nfzp029GYID8Sn
41jhlDqk7VBa896ZLYW/c9qzqGkDkDEM/45ZFgMWrqGxFSWg1mz875L41FVhia20rGNwGzfznBWW
kFkAHesZ6GJO3SewmdcpBVwAXdC7GwWuWVQr9ReUFJyxxdoTSW9+B3d8ZNKzC1PKzf4otHGfpK8c
sDj07QPU2Uu9nTAKDAxUIzkNAmkXzmsgHNLpweq2vuhzig6f8hxOk2ZocrFyH1lKhB0/x5mdLe1K
n+qLiu9uf2u4cKcOTK7jMN+A326xdTxrqe4qoeiqlxrS07nyIg2bmWkVDxIF/W9HHNXwyMM4aCh/
tPJoXy6zuiFioTOf9A6SO+oMkR7eUEQRGog4hygTbp5QjWdgsftGuRMLAOuD4wugy9SDtSnNUU2q
ep49GKmMvF5mHuZqOw4qAja4Xrtg9nA7zowglwrGb2MHwFnUWNa5jq1c63Mrr32g/hnbZAhGxFMV
hnur9jlSK76rG0Aow/VBPdXB7d423XN7u27HwBgvmsWdw5kTJxZ5n1oGd/dP7HWtiCVInjUU6P6T
DaY6+xrfQ0jl09J2ZyptUmTt5L26kA+g0cNRB04Sq8UPLmSSwN3eoZhqetE0Ol8W+CSQ6w6Ev4Jo
fUzBELOIYjxtnyfO665jMWm4LiD+DhLALcYuENCKrKQ5iHTY+VDiX2MmCYExmMxd5YhObTMiDEcL
uZ4JYLZNU42yAnBX+1Cy4wi0i/SfrkLUq/nWvtrNadxMPSsD9kYo/J0GXu7jeHabwrDHeHFpPhXo
wUjOlnafGaC+i306D88aGQE8lHOVFhLf2HHr0eZlwW4T55DY5DY9C7q/4cOKgK9RbwnqHufh0Ytj
m4izWe0LSXYXTP6VbAvE5oMpCYBTwi6jyMKdxg5dsaEsIxiNivuN0lHXfK8+jlpTTpiHpASTE5IJ
iWvYN4CsYn2MukVyBdzC3hLaotybAphlWMh4svwCIROD1m4sNqiWgZKLO7tmT6OROnlxetPjyBuf
JBz77JJ89/LWudO/CVjRkpwXWyaHOTbgKWLT7SA8VeHiveWtLvqz84J4CPFSUFI5o9XzqmgM18F7
Mz+UE+T69RKqN3cJNoH7l+yFIEeaGxHes47DHjRQdQ9DLnVM8zSdCEHde7/CXRbhgae00xxakgqv
Gp1tb8hgdtUIk+UAq7pBp+ZNAK2mI8JEshXwU4VUxBGhNBqQGSEMDsM2uZND/qGV9EiC/oq9sXg2
QbMkLWURWkLn6DMAYzS5aQ9XpsWu7eC5WpRz1GlgCGd0YG7izOkRRm9J2KbcHk1ZPgysvFaVhX+E
eEQQ50T4acuGqOwwhFBLgl+62/THELhJ3XOf/tDi/lIkhjFHPoo50W9jQzJzBCcbw5BYfcq3ebKZ
DqW5sfRi4L39rBefpiqTZdZlP5Ps7t6DjSBCytYjOEausjn6LhDdiHi9kudVqaK18dcKTb/LCARF
YIA98V4Uom9gjMI3tSO29F1Nmn7V3yjx7jMmqKeiE+nfeAl5oiQxjnqS1ABKvd7ffQ7YucGmFjOk
fFmJEQyM+YHIIBfQx0fRg9l+YhnF6bs4Z1lvrMqFqkDqsB9+0aYaBb5IVtyLz9dOCx197vNyhbXV
QiXiFHE3ZDYpvbr5kC3kLn1j5Lst2JlkIsoqTkkB16CIGkVfnlD90huTlLvr7CHaPzSJwgVQt9pr
Pqb0BA8z3kBW5i80L2STyLUpt6RzbMd7oCkXmojziRfr19zB4x2iFaEmQ3g3YpTr0r2dtpKMZCm7
ZTd7uVazzWVh202taQhXiD/s98rXoo4M6VRoDasKOTQVPvw4G2ZUDtR+iPL9ykcCHaRS9GDWs8qP
ApppA0thvcy1L6QkZ/eJ/Uk8QGBfqJVTafJwQ59IUoGhD+Zysgf/bH/3ht/Fu4RsEPUXzRb1Tdi2
/AsMNs98VLiYDiH1Eu75KKb7KqDorG1tb4Dyfe/xxBwKVD6KCb4+ooYSGPmfByfB9/LgUjAql0Cz
mSk1itv3F0JrrNCHZu4ky/3mbnurjbSRtrcQ+xpdHS/Bt1P60AVkNxoRkum8ZUdmBJYSRD3fgo3t
XXfG5sHawuiXG3cFpZCegyguC5LBi8/tOvtfgY7uzff1vDKVrusXVN+M9yytyaCg0shcWqGVRipR
S/Tbdr5ggbM0nLzvDmNEMY0cjqoagw0P+oljj82pDU4rikxL0lGTLXG3sUbD+nkMNKzQAj2j8QFD
59cyP8WJIvK1lgXBCxVIgJh63Zj6xJ9HmhxRkyb2oT8GPdxDar7dzpZedSLFtsox5Cml3pkmkrtV
UQ6Ve+xsIzmVDLMqnmaG/j4JkCMMHyutZw1Lu0fOiBcP2DIkv4a288ZsdEZji2IFD3VvCsO6oh6F
zySfnoCK5qgyxRayk1iYkTgZnoSjStPGUtDBKxJi3n4g2yHZLaCMvX5VMq04Wg8AhgJ2lWdi/DoK
0OZY6pEZvpTr5NaSNRCz7gHLSCaJtRNzOqMrRYYQjvErs+jOVS7/TwNiJ2/Se7/Wme3A2J7PkDFL
YQEV12Eod3GX0v6WbZ9SfKW6Wlpn/Rr6OyxwqeYvpzH9aMCN3x9DhAwFXYpcqkn74bMD2UG1ohrS
3KS/KGUHQMlGtcYAexG+tQZd0z71HZarJi54mSfi6uoZh3LiIbOqKyIP5gIIfazSqgVaIDWk5yme
CUPScr2TKm6DurBn1wWj1tu1LvujyRtMKNvY9HOx4t0MNvnY6Zu76RuRNkbVtj1iafDD86gbtpOs
zTuEHG9oYi7T7hZ2Ti27nBz7r7vR51Lu7J4eRaHgVOvZfr5N7NZkCz9dGmdqFONNF3bWzQHptBbx
LSpNAKTdESSj5rGnKhCQnWR/TQThAchlkddf+xFj5Ban3JjRRHeGnzKLqaJFoE6wRH8aoDzDV7AB
8+85H9caUk3LwbZPAJHu53mxaSNTc+2Jv/yRaU2tzgZdyat2YDlidP2hl9aruNdt91LPPZ9RgaU0
Esm+qlvqcz7/yWN9zC1cswOJ9iVpQbv+RtbPdRpht+UiERg0lUhFIc4OhAFl3KTXVGTLi5Rk3WG5
YMduZjSUwuXjarkN0P9j8ijJQXB09ZBvNAsl7c0TE2sLyiwN8yMH+I4dLj1nAimzuUoRuxP8oCmS
gQkChEewUAMeTJIuXO/ip8YnrcolexEYN+jqyAiWJCqmwzbdhJa3UZOC9wpAeTWP5lUnx+xqYpSi
J9A57QeT5ZeaetM5Qikyk4v7wKTdZFGcTQEHAFeqdbjVHXwc+3aKnde8xv1qyu+FEX8mq57GhtXs
R4wkAm0zltSpMcs2XmF/zb9N2gvjDIOoTSi8HQWa/flVQWmktdAP5/YcieDJarHwUmGFzVSihj2e
atvw3gB/VoYQT7JisDiL/9MrGcSUdX6KUgthnmfGU/gcz+0M3/V7UDf2PcUmPrIB3RZGeaW86sJM
Ytx0N6WTv30LzPGvrAeBHmbmpiHFHDa9ZN+6dzEmayP07XuxRdE2inpJiipUGq8kkizJjgRwtppL
wAlqMkkgJNa9c7kavfbo6wAay7O6YxQmvxTVVcOyrTHtJDZvJVyyDm6z/VcPaKtGmx8EYLvLoNWb
2jsWNs3EzAp2fHBr2IOvM3oYnLVdZSdI4MXvBzy2FaWul5+drtPDNZMDXUUmBxaf7TY0qYMzP0hJ
MIcX/FT+2jIoC47GanZibG7J04j9WzS2D+bd6f+SUKGZDCzQ9ZHtqqpgCnwuHj8Wj6NFk2YtonQN
VE7BnyuCgUhVkj8wKJ5A6S5nYQ5sJrEes5+vAc2YOzbOsSnJf8ILgSC4DkSJ/9ElnPteFFjolrzg
zYKyCpTRum4opOdlMCVeCxfI8fsL3EwKcNGkoebYSkFgnZQjFE8LKjfWjb7PsVbWF2M3FYC5y2gh
c0MLna6qN+SjZF51SUJBW/bbI55Z8zEO6SeoL8ahy2Xav6555hwS5A2teVwsF2D+zopN9sTTKMkT
8kRXG2rIyRFTnmtjzuwlzVX4rwsX8GYMwLjNC1bSlWEU5b2TUEq5qxa/t/qvRl//xK1VPs8sKnpw
XYDIFLIq2lcblZS/x28fich/cVTSny0hsgbyvaCmuSkfzZaV3Y3oS+DANbF1cr4QhMNMsdp00Y6i
hp7BNBGNX3VNymXueTdFK/pgWCAsyVXxOqLD89lxmZiUwTrRTeh/RMvnG4oYUa4ZT5il+dXNt4LX
SfZTeAmipNYV9TJMxIA5ndorLKtXUJSQPx7gPQ5g4EaYOjDyQepp51EhZelVWn0ud2Z4OsWGLjhw
gYI7MbsDp/rEGCG+rzTjHXiBID6NsLi2+PKkO3KcLb4vi351D6X/nBSwtS1DXou1NkYaqpsZlFgg
uRLqLqOKsxM+fc/zg14IjCRCmW3XFlPmDv7zrBHzU0nvbRUeOOJuuzVMbcKqRgbppJKq8FbtJCIL
n178fnaeTtiElBwCgfqCwqgbmpHBzuc9nSL0nx36NHrQE4IYOwKUbrbafUMQ2QfPAvH8NibXDDqx
q4qOcZ7m8zY+zmsb7K2r+3JFqfabq4HF4EMRRvr9d0CzGFDEqnpUYCJlrqdUkgsXERP4JL7GKoSb
yG8ihXKzbDGp0W7QVPm+AoCE2NsFrTLB7zSu/s355H9MaRjnMsKVTmSqy3WQyia/DuxbE2BA38k+
BjUI4VOo4myE7YsrYtkMlmGG3uAQZ/9BXIsNR4nnWMk0VATDDLyfwMmE9sRwBBSIJmw6+KS+SEqR
u4uWjoy9zKjAacYUm6VUxIp3DLX0xNDaFuVcnDWGODFgkdjfLjVRwss2Z1JEhChAgVC1tb6I4PJw
3BPwl5DyrRKID0rNsLa3fftx5f7v72B3VYv8z4Bh2SjeV0Rzji5YXqVkEObsMsWEMdUW/1lkCKnB
HwRZc7cS0kcAcne3Hkk+93FjZYzEMjyiWEgGsi0PYqHFKDcFslHw9xJ9cguanm1ONQtN3wmVSIA2
oY3gbgNceFCovJGJGFPE1bluAwaAwGUVuPNt4np4Ak8R1aAnkTIVKZpWDhztKgR24lq380A7JbkS
wvrQheav6oekcx5P7dYiyZTdmgq7fxWyuRbC/fNYB8ntpq5JmBZ1zGIC9RtuTpO9bayHg12wKBb4
+wA8TYRYjIiyerYkqhiRNaYSLVloCt0QM9Yl03qmv79G0Fjt2NWuq+opkQ7JhSBh1EqnNgllXxCg
ovCFq9Adl6cROU99+X7FnBuNwg+qux9sUQ0xjRI240Bpzl6N3OWRSeiQlCAs8EhKyviKyEHNoN9b
Uz/kZeU7XRLe+m9FBMJPECPS1HnP9XV3glOjxG/jO56Ygnkv/QRsDU9Miz7jKpFcdGXtCpSEXETL
dKT4nBnJomRkZAslFbH5TtdN5ZsP86NBW9aBbmYW87/K5zzbEswik2eEA9FhhRIy/hWe9Eso8Ztr
90S8RRphnmDgFtqQfTzmD3Vtc65rq97I+dfx14bGhsapvx+MOWBfp8AZZPoouYcKEUVDao4kUkqV
YG5tT8DB4o0yeYTGzey9CXBctVNAdvv6WBzbI4YGtsoTrRqACDD/MFvQQ2KOg0oyZOgOa0nrLroS
FKGG4dXSMN2+p8LuUFYclnORHNubjsCEZycqM56XaUBkE9wqjyvpEG5QneHDccK3eK5iFI/zJvAX
Ve2D0GU5xZmzyEIGcvz4hpgKrecZpEiGLRubz68U94zKwZtxC5QVt1QGIXvLVIsKivMlpkMvLEFR
+oD9feb7erkZKe2mxBUU3eKBnUB5Lm8KM/WHm67Y9a7o/ZIPf9qBOqdtC/jIAkCQ1brH00URFoCd
q7D+3wmDYLt0LUjxLqUyMPjcbLiHVOD43YpseD55RFhqt6pKsHfox6SEb+npQABMiYTPp12uI1nV
7eHUWz82gQh3w98d7MNGPpi28u8yz49v5AxgOUhqinmHuSnxSkRsJcQhYoKSpgvVLBNSNLBDm1Wg
2oWyAWZ4dIMDDRlolyx/Bh8OKfUE/T+ZLztB/yyMcz6+Q5vXJIfLtnEZXqQF3xj/0HADEJcFh3J0
FGsMbGVtM7yMykBRxxXrqvNRSgHBepbe/FijcfK8e1UfZq38Ley73peXlwt3OneFpPDFJKkyo9qz
syKgCmaxs58zH8eXSybaSXYUQSE5S6OrNVnY11Y9WwT/pgq5bQX8tO7eEGClFr2u8w5QYUoQNh6/
B/XcugzgL1uzyjxJBrYMfFlaEXoNoDEzDM01AmaPxzq5is0XzKBlTVIjuYFWw371TVyxWeym77K+
iu1mPf2Nq4uGznMKdDbyWphpZVeV726PARTwDv5+5pfuHpj1ETIvuuujpxFyxWKiqLJIuUP/hkcG
AzOodbjHPAsHA7DPuxiQJ2wu0HYnRkY3wW2E3kGbPIvMqltjnYuxmhXi0nxPP7dceL38+Qq8ItOH
xo6sJGqzlqA0i303IcXcj4PNWZjnWuVBb5+nYVnaW0w7WJ2xVq4XOJRgcQRpQBtKpRHdA3HSZy2W
b7jknW2zsA5BdjkqgX22zecui0kPXEZnPiZdTutjk21nZt9qdItDS0F2gyVkgAKnxRvn2rSejdEk
YDYP2NE1z/VXY7zyuXTKBt9glt83n++Gr0zfuNmBc2JIY00asMytZp/WEvVeLeEKgwx7I2NolQDf
iO6ZWEsBFgjdiMS0S1wrtBRdpxXNlYAHu30i8rN0otjMqzRLbXTsWBSlCxX0g75v4ckOcYz8T04z
lb8MLqU1iS4uMAT6tNl9Bspzx+7aWrigEEjm5kzpQKWi8Pk/zqxtGHwKbKsFMjJIW2viYFeWv2Zv
XVgEW7qNUU7+u6dFXV+f70NXBgSIwXuzrBLh3w+iR3kZSP3WffxU2lbyjbuMMvBvFF+mhjJyfDKH
IXgQrK8YJzTGtPdrHxVXoC1f0zTaPPNlghcPi4D1T6e5sqkEj4UinhfdlGkE37goX2ZOVcTuY6qW
9EbOysfsvOvAPINNHZAT5SMCIv2HXACBP4w348CX5nBL7JJq8CSeVSMJx9Q2bcupT9/ka5x6nTxY
xfM/nlX+WVo549zg/xFSRR6R9omKzJV3omRnhI8LpZ8VeFWZuBNNsFucL41+Ad0JhP5wVKOMu0XL
2rp/TlciVQMEYdci3nrehTCsmNmtwVw0JjIQjdvq2iQg/Ro3JXzM5tnUGcsyHhTYSy2sxWReS6ZZ
IesVn0O1ha2HfJoBCjH0OfTV+ZbBPmVFdLQrzvT0kHA4VNQhYn8G+R0mTTHxLuIEYZHkdHayUV+2
clbSfJd/tdp02d8/NJO3dnjq6cmbw4tUZFEBF0y0lKKXFotkOkCrhtAYIrrfrrhkM8thxaDR7wM+
R8Xq2QRrUDs0JeggmsYbDH/CBd6gqsoNgPXJU4usDNc2F3zJ+nK1LpPnk4iQ7Dylv5bRYQm1L19I
0g0bO1apvvhiOI8TvQn8PzhUglnxLIq+Uc9BqzkGkhcFRmYpYTVRg95KVSuA2vT2vHItumKicM6I
QYDSWDm1r/9Dr6x1bLl0JYtX13Vuu67oJN7LLVIZIDe4sLJTBlZDGYUWhV6uXWDagAcIQfV/5rIK
jcaDxXe9o4XCRDZqWwrvWbbZYcQ+SBK554xrZCtzl7ttoOz7SMQhj9FfNZTDvGBOAgAyD8YDXX7w
atxd11HRYwMann2QUeZxt2TUJqGd3yM6lZIYGDERL+o+Wkkngkxj6/OOQvSQHcHruycVFOp+sBwE
ld6j/0rXgHCdNuf6zpS1CZjhgpo12pcfN8LzI2jQvuhWen5hSX4VoImJeY4aJD1zINpJ6nERQ1ug
LGePYzQ1aq7g239m/A8IPJCJ6yft5xQj/o1lS1D57UlWMZ4g6nlile+bpn1sF/F5QlYyqsaUOZzE
ND7O5Ttre0+B+d6SE6uUqo78lSBUeq10TE9lttDYlrC/GMI3LNKR3dBCZrvHlwhltObqhR2mEBIF
SVck/WqlAo1qOPhLsxEnlB2O7hQDxNCGUQI8VKSn9OgGJT0wBwihBNJxKm/f213vp3PWZX0GlbNN
rbj89JkJcJnCj6qFsqCFSQ/yqpL18/V5XsJhKm4VyrD//ROilfX9f4WsynYktA26tb6nt9Stahs0
5juNrWL4OrIXAX0SG9V4IZOyxMogzf7VU2d0zy/OXGbMXrL8LsyEe9yEohw3bxjoqueF1n/FuObm
fjc6X2eCVm7Ni67/W3KRhYKF08vJCfx0FyTL4YjNIGQMi268HR7Lwy9NGvxkwm73LILphBnYMfbj
ZmmSqtMGfIMyW7JXHo0fU0Lytr/9p5qGbKJAo3tIT6igrRyDw8t4k3Y+6Q0nWjDkdilW4SjbLLOU
Ayc/zab79udpl3FYNp2M/NnGi2F0js+WhugCSLFneWYXKYX2Uhw8wLrYG5Pkt+H4m/C3nV29cNZs
P/3x0VwWp1T508KBBkD416LfZqEPTCSd4T3sl4e6QXyGVC0RkdeyC1EhPQvWbmLFOQH+cMU3zATu
abOgCIlGkwI56KCVUX8XLrzS4sinvgQieuUsp2QRiQeYu1aqS5IeuI2upVevecAeJj785/vubg6n
h3osPvg0lrVP9Np4vYGF/E3V7j8VYkQSB16f12AaHx9LdtbDzXR+nSSotDNujDr5U8D0cfDSOmSb
cqpIq/wfiWBxwcNoKO68JrL1gPWGND/dQz/2NHwEn2ncxFefsc6AULhq69edSv4/PBMR7HzZpWN8
Q5GNi0sPu9qGz+tGPgS1AgX7ktpk64EeWvFy6x54W7Xoo2PaPZSwDbjhoSAD1IbLjQYar/jKBktY
m0OOMslaulcj/jqspkmg+JHpjS5vovr9UnSBEOaE+qfiaNTtq03gMKb9GDfpHeBfg7TLqzr6A4J/
a4juez9YzpNRt8bY5b2e46edXzHcjJFtz7rGBWY+nl43EzWE088G7S5LD3O52aDqAUjBkQL/z8rL
/BM1SvW+cdj8WckzLdTCfO5/77t7tUCJjkYra/AXuvu2s6J1oFmCa78QNvoGtuJFAZFxLMLeZXqb
gZ/ryNj/hXPfYDFjlbVFfSEYO+jrU7adKkQ5j+uGDqCcJUn2B8J9L3Fpinuu51SaKoGFSZ6Ubxmy
iyzFnwvHgARwkOuyf2gByppdwdBEM8uLX4ipdiQdjT6BZJ1xa2agy4iPYPC1wTNRe+hvVpPiBLsg
oyc5L8BvJ/mCs1tWxmfe8ulwz1xbBTuceWxvoFPJkxMcdEGUE87IsIpGrRJ2nc1V8DXy8Df9247r
+8M658cBvjmJNAb8Is1rZVFlK1Vw6onmalv+znUwgQsG0LC0oGNnsmo9Nk3imX5PIZZTdXe9TBC6
g16fMRXN2ePugu02URD7W9i2422YbtFL+KwwIrgNOOrmGDjDOcXcivRdqaGs/PobhXhwguHElXSZ
jwMMHfEyMFZIgfM6t5lmIqlwaZSJy+8ZogVgua4nfZwPcEqW+wXY37o1AeQ0C9Tw8LExzFFV7YbA
JrewVh6Ttjwaf9sNn0Qwo7uBI70VE3F+Z8igVez9etf485+3MlArLatGHRh1IeS/W1GvpHkGSY+b
qqiayXQI3AJuo/XiJtBW/joMPwRpnxU0vVnaZu53gBI4sE1EvfYOY1Zr3WumZVe5mxh1UfZpoF/U
DFOVAfRerZdgvfg1me0hjI8RIHGLQTNxcO3vubkZslXg5+KDgY1xw5iNlkio/hW3Zdmi230VEjkm
wjlCkgP6x8dRnvYYuB0tPL9Vi8OPJ5yzVqPNJvUkrvpTwfp2XuGiZV/T5XtHRa59krkn/K4k+jVX
93rKs9dUuaZNYPhca1dnKFAwMtKjbplrzTxTfm3041EIYPlqfDxtOv70fmzK7PF3F3RglAHO4d7T
UzzECgSmPqekRbxRuAjAT6PQvGAJUj2A/kyF0Y9l0V7l6KS7ArkeTKlAsiJBA4tLIEsrlJaco8cm
QMMZ2tBJ0CYwLfMS8x2DPxVJ6pscOZrXArShNtkVrGDj8mlZ7DPI2B+wlQwdoOIxHFyrix4pxxEE
4iqSv+NpR4l3iF+JZlXjTn65gH8vlY8LdsCFQij1aTi7Ig9X1XjxGmP238Scjk3MSVmmikpmiLSt
PWVv0M0h9M9mqq9KJvyW45ctproekS+udeMLkjl+jzYadQYoiTlIikBTinwldaZho2UJso388fPO
E+ti7XqM7ltpU+5M1LfwK49zqX/2KWgfQPLwTMFO+HLPvQTO0Vo1v5QupMVQ73dRrP7LJfv/OiFD
rZZKWZWwF7Cf4nZeVsbAIMgyr521IXO0SyW50j9v/pLmoeNIF+I93fvHSAH/YToo4BtgcpNw9PEC
a2s7URjyVc5wPexrKsNwfitfig+CflxGLdw7LuPnyuO5kbKm3h5iH+Qy4dKRsUrvUajr7qfMnOT6
LNfMVttnNPSf+ReogUfIxa9jjUQQoTxxPI8XujGUE7GMkJQ+7mwO4YhWatIhD2mjJUArXgp25ofP
2NRfEs+yre2gSTrvfNSk6uU8Z6YYkwwoXRPfQQnVYVjetzU6bL9ndVIvLNCEa9wMwjAeZ2Fls0eY
7+GgIe1Gkndka6BPBGZAFIpvEgZQyynp22YXG5Y/qk3bTY4sIYJQZABCUkGO1eWuBb+wOkv0Rc8Q
+R/xlWcrRsWxj7uMFIrnz1fne9VNwk7Xrp6rpekN0PVxUcRxyp6d1Vp7R2VDivND1L4JZ9JC2G5s
vShxP9Mh6+/xRhRAAY7uOsPOAkd0/8X7jrS4p4XylyH/b+iyx7jVDlo3C4ksk8WzqPnUsWD2nnRu
qbQ072QwjqG1b7Z58pSUMIpIppf706wL8F8fmK6+l6JxYAkra5YgeUlfN4hVCKvNbNw4Lat5pfNd
tvu/K1R3ww7c1JekTvmVIkKK4QpOzC3iVe+TDcKlSgUXeYiPqd9eEyRn9GIsmFC3kpDksaeIoSTF
8w6RQ9JLQbok2gX/+3HYpnPOYLwFk+v1aTB8+hokH5n0pjFyUAsr7KF7UJXl2ZGQUJEb/Ivnq/QN
Kr5xZqAokBvf9RNasBMxlK0GCLRIWXLsPsnE9m2nIswyi3ntqSZtp9pgjos6PRnwcTWxjseN9iec
u5K90zb/ulbWdm6Z9AliXsgjYYNaPjbShIhukPxT5olZLaWY9zf2cDHRQIlrLnksTc61gmvKqiGl
LmYadcSB/pEeUymjxMHFnc32hCh5qD0itxslcd84qytofcAQj1d2QStR9oOrsY9Q6jVEUrA+WUL0
pS5WloR6ONk+DFb9WFfnDUMNSsJYPm1ZAHdFcXb3yOxhrkWVcH0ZeTaqEFZd3GnOgF/CQBjiUiR6
ZyIRPphRGF8WYLUa959qFwLXUqTmYv501viQzW7cwCd/YxQbTgy7kA20f8XYIlwbz4DoemAwwXkS
7o79IW+ryu83sWktd99Oz2xixw9QxA6shc42yoEEWnrBCRgjCpnLJim6fR0xxhdcqHyvwhGwJQLw
Kwrf8Vh1oat+MJr07RJlQpjHT0CH6fyMgc0VVs752GODQ9rv9e8GhMXYTohPjkLmD6LPOTU/mWQa
LeyA/DuZbfWsqibV86T1zAjkGCFS8cMs6/vvQAR7jHp8eM1D4imZL+e7HdhC6IuGUhdYvAsQo7AV
7u086pFpDoKcoTIdUwisQbDaFl8EgWgVqdoZ5icohAvKpZ0NRDGUwYH7k5V0TAshUJTkOkTHpleJ
PEJT7qbvYmaE5oFEBDs09W/hTgxIszgJlVpruQp85vdoP8tNw3ZXpDmgAQBrOv/+0aGUs7sNPVAJ
3lvotub0iE9pAW4FkhfauyG0HqczfnL1OzWu1sJvJ16/dqsmflTFNSIpokjPcXrZ8dlgHhgRVI9T
56249dvYH5QD6uIVcKkk3pthYNEF72PUhqsY+mv7NKoZmO2NutC3qx1envZe2y9/it7PZBh3piKe
tepdltkpfcSwueiCOTU7Nt3xIc/5uO0PyOsg9KRIIStTSoEumEOOYlLQAnIHacmMBGZd6AihFC1F
CwK1ZEXXrcIqB0X5zs9wtOcQhhsxkY3ocAVi7u+HzPfvYcXTu8bEDCwhHKiESL9bO+cGNVeSlcil
Hx9I1pueNHnLVft7c3AikehG0QsfkrbUkE9fKptM3Ld+a+qb4rbphwL2TRk51DlKgO6zETHI1HYY
/1aW+nDPVGwRQAdzCBMvMnwdWmbKaWPHXY1b3X1g2BP0IQOXwHD+lCH5WPM85zsLRl4Z/nk6QyPW
XdeTWXrSy2nLFfy/X4k2UVFmQ5ZSUSan8rMLsTIsLBuIjMHcIwjp7JktXKl8KKKVb5DnzWD09rY2
V2Dfw7PoYAx547Bxx8C4vLmd5lSG7KYoj+jfeLHGK0+SMITKd7FGhE9W3s9PTLrikFmxc/0vUKak
BH2fP9VUEdkrhi4LMvPR/mcnYMsMDKFLXd9dDvE9X149gwJxwmAigxqxaT+D/i8xZJ2CtCruWscd
RdPHqwMraeELUGMVfZVpMGLl/oeGSprMXJPlXmLSXib2BDB0/3D3S8Dv/j6E69nmCnzya1r5GwkN
S6919bG9mnRlYqOQx9U6sKEKXpHvuUPzlLWMUgoQCs3BC3aSkHrH7NLZ5xEH9mKgG1ml/+6hrT3m
JPdthlobm0/UMwuYxvmv/ZBPBfhtgSeHokPrBTYBkb+WuRof1jypg54Oh4Y1WfzTFIdB0NkpBiIw
NWf5fsmkbadf/PE6UMyu6uxUxjReKgbAudBdDZqiYJLzN9/lrnPOmFv/NUSOpSbV+VxvTRo6DhDA
YmX+819wntofWfdfeGy8+482kbK7FuIm006qv07Z2IZg/Xop1x2G9FPy7so4k6KjgKPu5Fgoc41o
nQcia+hZFB2bnywMQtc2WcC4USjsimAFpe+ebjP8G/MvhAH5vmbuF9xZwWFp3opn5VUQBI5Frl4n
jnfZ8G7HVIkN6tIjzhT+S3K/M7hcZR/ESotgfJiqdLdKH0NPy+nWkxO49DgRV7c9ETgidOXFlBxT
rYOO9RAOUcvJ1X3/AM6ed4a06VXme4QVYmPAcxr49a9MdDz3Dg4Zv+AJgaXBSW18KqSwRM5dK/xG
fsp/ik0jpnmbzd9FkzIhvSqIE9tqseKheGVPusB0bp0Wimc2yFc4lTnQdKbr0VJtma95kfFmDox9
zzWCZFn6OXcX8hb+Ll9F+e77PIRfqvS9hhMWxIy6Aupx4Tx+fs3aJUtYmWSBVnq2z0+8ZqRQ+LAT
m+04ceuyz/nNk3pjjc/+m3vYJiq7g02ZOzxq4QEIbeZFIdKNqgmo8LPE2vZ0UfxaZvBcJ2xkE1gt
ddVI6IFyM8XeuB+H5bMjhqnBP9puKlg9LyENOS6aOAprxcSVf1BOI42s9Z4Z4mD19IbmAsGk6F7e
cDL/R5nNxfBzbE0LiMpLXGPmkJVqMv3ibWF4Fp/LS64RNcJZ3nMBguJF2GP0QGkihyWDA7vkUqBz
N1zjp1b+3MFtsjprf5DxLQheO5obZfsjdX7CN1aixnq5LxHmlIVRMjex7WzPnZUW6923qI/CGSQ0
7sZjCz0R1Hw82kLMcNSw1ACSZnriu7laaIb7NzXtjaR+PVC25Y9EsUqR4Wr0gj8N1er3/XSBaBTi
kyfuaItMwlDdO5YV3HSq2OYtFI6S9jUfkW4/oPSwJISDwcxikhNO6lSktRP7SVpgeTVJVnUl7a1S
BaKfx+Xo6nv4tmBsUIHASRyHgrHFTOBT3EL9q7gF++VnD7oF5Kx+B++s9vUIeNuk7bhLT4uR6PHR
ch7c68bzDU/KQHf4FCFIFbheL+9bljrSukflLTxUvL1s1ctW4qGZXNFFlyEOfWleI2wKuhM1S4Ig
TgFARxNDSO46nTylz0uxV9XMzZe8VXQeDiMz01R4h9RY3oqVclqSg5yj+9jNBK8vMX3v19zxZ3kS
UUysuUTykZfAZkgPbxU612W+W13pyRqNqOJ3hf8llRnpknFEN2Zo6KPt7RaqkhbxVQpI1uKVs2ZL
QPbpdp7uo5r87l4t0/FbGsln3KrYkEbs2qesj2sRYp4DAE2brJBRZq7Q5KJk2dgvXZNiHzXxrZb6
d/Xx3Z01BZQit1SMAXbbH7e69uXxCodMfEtCAyKqsH0Am+Q4jZaHU03kS2vJIy5rVc8k1BEgtQkC
+2yrNzhStl5e0bxU5aeAsMAZaG94oDCtzSqECVYm6nERMMzNOEbgN33zReV8wn6MecPUqQadYmEk
VUBpqMhg8+WY9mYp25Cf5+2No+/kJsEO5ouJ9DOXHmFShk2CJF24AzUVBaPUUHFVd5U8rF+7r9BM
97G3I831NsFLSk3mEjeyW74SQblb6YiXgr17uc13baJ1lvpa+BnNkdkymRdf1PXmMhDjQQ9Yhvtz
tFdXpU1cP4UvQqznIfKFF2n/flTkvSm7aWkql80gxHaf5hvFvrnPyL4I5+30Ah/1NmfqmAacDU0W
6aUeVZq8IBGhmGIxz0eq/R+azuhNw5j2AtP7DeQ9JMO8RhdAVPf7Zo1Sy3LGZ+2PajfwikcpJ6v9
wFjgXvdScE8OuNpKLGlShr3pqfaVcWUV36pzbsJUxG+s9deggYpID1Qsida6OTlXT/EGUclBH06M
2XElpuY6kdKVMBMBXkG2Es4G3I+yXk7+3shO+LfuUPyKFlmceYrCUpww8kyeyiaoc6WiHt7+ysIC
isrZb9st0riV1YCsiIzH70PEwxirhZuKacJrR2y4z8ZR0XPfROvUvYXw4M50bL+k3i95l5RrR8Ds
qeW3U6QrJz/Vop+c1zx/duIsw/zQCWe1wkdjJDx3GxL8tUVn8opzaziHgkfh9QxPNzfpfqrBAFQR
RkI5RmcIG+KvNWJGa82IAGKCsgLR2p8LKD//LNJ676BmWcyN5A6fDwkyr7snM0z5ACx7462VapT6
6wwLssDa7uyAOwXJPjN9CR1Ljhs1Gk+KGdIzNj75ckxkH/jA+SHtW+tfoR9/KGwkkWKPczVU8fB8
aRDCI+zi+iGdq8bgnVVGzr9q3VDL6MFT8ZSecA6rOrp/qB0av4quW/pMxASIJvHpETlysFexpMH0
ge1axweSSbhSzPH04dP/IpirHnyLDknrx5D5NAgMYCK7V0lZl82veLfVI6vHpVDynvk5UNnCcu6q
3zJpVTH4ryoQARqIOop2gyax5k0YuW/3rcY+qqQd3HNfdMe2YM+5b6jM299Tha5cq2kdX0eVbD4g
GftNwa9KgIF1IY0f83FyZ7U3Vvd1ZYZxp2JPrLzwhRm6W0sVB80mVW1z1Ea5QAbbqhQhrjlw7FIP
U32WEv4oFxO6wsozPX3SwYP31aYAXaDslwsblelLayOnJ/N6tbNrPoUb5o3dHaHBqaXY50XonF5z
h/LTMGlXPKcl4rvBKzErM6I0rvLxRzukH7+4tipuhTt4Ff/stZxvIu+I11QFRFwHP0D0EfszCiOq
Cj8CeeU7XCqQnuyvGKKNl/xfi+XK0yHLhLvtGKHp4tQan1UCfi1uKQ8FKqJ09VyJoXdDpCAvYZiM
imIBhR/u5CIf+r8f0GRQ74djkuzYYJjIRTrUyR/LwN409vfWt9d2WLJapRKKEcn8bSJj3tNI1s96
4b6cipl4Bub949B3RxXFY75VPYudBq9trJqBkeKv9IzPd7H0af1dlL3/bmt2akepSQC8hWF7QUFO
wa2mNcx7AmB7bVbn78xE7tWyxYlKJ52rHvxecaes6N9E5SMe6osi65JZjh66VJi4OtysMyIzjxi6
8Da/C8wXTAW196Br7smttDuyuhduzO57DBNzduA6DfKEJoOFqdZDwOi9UniaacRVP+H4TD3l4LWC
8XxwfN++W4PNMeN24bBSKMPcwU6fC103iV3fl5zt6yVj66b0tc34fF1XTvemG7aKHxdVOtP3HUnq
x69UgMzL2W95l4yBwPm+j9RNLTOowzrVuK5WJ+ZGEqFNSUxch0TJPe/xNDwEwPv6Y8owN9zCwW2Y
U7kHU4V2fLZhO8KAFpp0VNN5NZZaCtknEO/IfUUQW4t+FXR1BpTU2C/5/n/UItrHyv/op1/XVadV
lLbwuqQPW7edVLD1/GuPSY7/Mr4/6T+T2yqgKOhjl6dLlKSTi3UIOwrOgwmwJsokHeHs4bPtlUeo
R+CNwib6fU407reY3RzMvqGp8IRaGk6c//hXELYVFXUpJHC2wqEmutqQMYrRIpSfiO//3m3J2/Aj
pMAMbZvGR9PuO/U6txIUMuSyYMkP1liROlsiqZ8cUFjaasCZuOHeRXaVvjLP707bnNjv0yFodCfF
DR4S0LAirQw1xEqhMvQ2eKeS8dn4cg/MYzH1Vp+jj78FsI9fuzDa6HK0Szp1ts6CfzZ0EkD9ynsh
q6Lgab866OkmCVfJHZV6QBgBxpRHQiWFdczvspUJ6JigZnde1rqdqrH4bl+s73jGjSTJcStZPBQj
fOCqfH9q3lqcP/hBGTUM7XxMec9tKZGmCXeMzk+rR2Ke2JA/5LFgTPSEXYXT5ZhhKIBCVvN2aIR/
4Cvzs74LY/n9dP2zH1tMCT9nJMEUk7lznu9HZPK6ZhopeHKxfKoGjMRDGLIGGOEFmT2GUuaR/7fl
ZklRXWsWKg4R12per/yE2rAEr/BIASnIlonAIBlRNuwmaaPAJmmPwvLIgw32DwNBS/0oXmnS7UDU
XUZQ/KLcBmXyomFwRBrHKjdWvoSJyKTnB6y84D8/VtBbCjuJ2mzHHnlHKlKPMc9Z66T/8y3t9DSx
avlcgr2LyLlza2tX+njFgOP/i6nWBrvlsofdfoCCd1bZ1UQppZa/2oK/jK6z0b7mOO0knUv3a20F
niGrqxBAO/KVXVq5KzemZj0HS5Y/nO/ZLieqw1Hotd6hNxx1+iefVIIVEjRXFZVFddzzfgG/iRuQ
lMrV+NOAA+S6qN0cru1KJOOLY7zLFxTJlF7rhggNdWf6RRlt6DDUgrL+J/aaiP4NCefhhBQQ9aQk
+T3UvtIc5qwb2cBb+bDmWlrPXb20lNFtkXJGHrmKVsL6prBBkqcZhDu2nNY3VoVCqPeCH5hUfNM1
MgKprDET5/jzB/Ql45YbE+m+h0ohccDfD7+AwQ7cxiMAL7Yh7LLSkXKSSOHDu1c/SffPa6mnhFh9
pgJlYM037f2fXBoCRVgT96rLSnUCQ402LnOtUXH+2mzTgGXe5TsJr0qdHeGmpOx26aD6yok/lVSS
j/7YQ/9tmJso1dU3FnmPvS1dyqbX7mnl8pR0B0cq8WqrI6aRIQyWGTQJnUKsQKmIigJ6tw1QNAaB
JdP7f3ehxbrWtLZMthpTULsVaaxp0E2t/gAXjnqzUDeGJD7Y3ws75B8n7vtnUPEnGx0Eiy/YUkQE
nSS89fouVMYZMZXrELl5N0u0JsxQ+SQ10o65Vzh7ZlveFBNKmp0B4brnXqvxHPDM9NqbhJ/2vhJH
nJXkPZGneQTlqzz/NdLHS6rOAhxyN596Ortu70nkZyzFaosNbtcjQZ8EtkS1/wBdD7Qrt8DEQxPW
h+KNRD0Uy2yUAShszPkXiTnZtWgYa/dTwYZgK4MI+lRXQtfXrBpDGVGzFe/d9GyTeyJ1BGbO41RW
b6WBMrV/0lLtR8hg/DIht7glrNGX/Ma7Wty3qR+nDv7bnZnxCD18fahuT7wkO1gp1rwyRyoDXhgm
m1Zz1LEADr4WZ0pGdstRYfDHfzNwg4A4Hdfk7EF8cL0jNLe+AbHKN+62E34OEfPfSgF/oePC5bjW
OgvYyqr1iarKou5KiiALrVybUIIRo22QFLYO+1LoyfgqwW6HVqFlvXHqz1GRnrBMtlhifScMK6fb
th4AdA6amQvxxT94CVroO4qSZwLQtXdx90UjqHcD6MxakQ4tsv1mCKh1wMVLIagaQtcJ8YHqfXEF
VeQ4OfNwaS4IgtyIyQ8/CdAlxYhJ7SHDJYrfHEdGHffNGhRZERnWJom6Gc0181IqY0OVejHdIXt9
Y900xGvf0d6UT6Bu85zLI5PsqacoYCerbXXU/1zZuAyfTwKQk8isTTC/c4Q0RMaxhufZJzIVDUbp
J2m7e08ZgXVPIvxTRfMt3u/sgYiLjKJNhL62KR5SlK9PwXDYmF5fvOQpj9TMC65xnMmi8GE1WApV
69G75mQFndrRXJfA2wu2MSrDsYH7Lmy0fkAsKpoR1ht4YK+bGWdevkVCuA9SwopGUMs3hkM4HRve
Xaau4xch1Z+RG9FhU87UjPiPAerLBr4lj2X5KvRsuNAHdydOP4gGhLv2RKq0M5XqiG9BWRwcFWF+
yQCcqDzfo2fFB+OOh0SkWlMSm4pTHICcdleeuYafjfg8CDYGGJYDJ0iu/PxbpxKdd5vm6i94vR0m
NGsj74YFayFVAu5+QPifvespTC3Fz8JKuETYfQC7mh32Gd7am9oPUtR+Z9NZZ0vBw8RYhsgqVR4q
YuVE73qCL8aB9Y5Wm6YSSY3MYDG+UFVKjI2lWi2J6S792MIFxKjOxtVyRKnYOyUdn/RysCuSOGX1
N3ZBVL5t0BzwxnXYdYm6jQ+SUo52280Bsc9DLDXZw3Ft/vHHDYXyQ2yjB3DI5gKPGfuf4mpMkaP7
JoTuJ/qt5oEwagi5chR2+JEUEQry8vG+2q8SkMm5h9/A0kbdDhfaw80lWnda/dv6Rp/tf12jhl6f
sNbAK/9EYBxwDT8ipGQVVwqqDMA6NGM4fAlo61cHX/KgPrO2vaXCcgvsQ2BSHghjZoQIdH6LHXdq
iXs789ZZhzaRVFibMQcEyN0Mw/h6/b/NhS/FmVP9M6E6arou7AOpGs7BgG7ujuyYXAbqCmjU8zw6
Q0FPqaM2umrFbwbpTRPJcVUQ6qUbXVNmWGUwLpSdLpdvVE6T9OQszpwNy2fnnxQNfjWkOzAK6TWB
XlPvaFWMXhbc2gzEbJlsyPeS/7CqylOvrgl+qtg9wp/2sY3q9j2MpOdxnBt0WqqSLEVj2sfGLeP1
b2MoYnbGXMwHQmnzwwhBa2bBMmda4Tt0LNZSYR7PKauBiVUHF5MNDZ7nDEtl3K/+yeHcIh3+DchD
Kx9UZUT1r21NDLzKUVYLZX1O2L1XRdWLAxiEe3TLkZ23sdOkoLGaNyWgmBxF6x8hEA5GnTMviq2l
a5bZVvKqPr/fThmB48tkoidEAis57IGMATDPZgd+bdM6psiFs3dzePMLeWniU4yNHb4UQXfFBBgO
13xOSULnEBl3RcaNbycG0RyCvl47Yk1RazkBjSii1KErx9BihU3DQ4QzNScSprElYHR8GN6ZSUy/
nPwW2qCaylJK2hdG44cORUB0QHEDF+AlcZ2QZ7wSnZJ7d8QO/v0cPtEO7B9d4Fi9cN9yS4eKTXJ/
LE/U1rEGDMZadIJmPoLi/MnHqcnxFviQF4zYEld2zkiFHTsV/0MUMAhZJAKpgwv9Tm8iuXMXWZvJ
oXxQZwAADhUgkeRaeTfhJnVhGvbVvA7PCqVHW0rw7VPU5PT6TuK/ao3uTG3Qqve/Xmvf5jjGdMOG
UzQ2G09B5QT2bhOjR7+uOTsIGI/zYDyDklSAQjI3OHF5tCFZXRnAc0TrrsJFr814DC2g8Eg5NCqJ
ePyROBJaWhJgy6Ppb8RnQHAWSqQhDCB3l22APvTgg6+VF0S7b/bbY+v0HaZikIf02inBHqbKHoWv
7ZLRNbNJoDHmhw06EaePAGuwgHNLnM20V6ghyKGXuh2LlXDB0gGLj1Ae9f47ir9W0CAsVyRhqBSz
kbsjQa/HbtHnPZfURSgJk9jQ34Bm+a5ysvSkKZHfLwliY9a4zPv23EEELnhzaCHkK3VhMeDacTUW
zhgpFFseJWiGYvgu2TP0d9xBLWQp1mZhlkRKTmU+SBKz8RCqtZFy7HLYy5CrcNmMvLIXYaXQZrE+
Z1Qui1hD/1sSS4vrREf5hrziYiCjImt61+ocG38HU1M55vLpugJw+iZXTn0qLhejXZQZs3j+xYgg
meWeDDGzwKaCJdS9uzC7u3CPigI2l4jDGZ9+2SKC3l6xKj6BH6fbcdD0zQOJWCMFddNNpK/T2Grc
qLkBPZdrGfZ8bCum1BeZ1DhK1ueYVYZ/IGXg6vrVWvjx2oGORlDgD/N7LrqzG6ONMnJ2lCq/hBHe
324N/gCi7CT1zK+/j9fggd90pzGFrujQvRFjeiYQQiBiazJieMzy3TAZKz0CXarJDNx+bT63s2n1
FgTkgUyEnBuHiCml3Peu4GAMhFhCD2qyWUkRtlb3eSmBT+HQ4m1XHxJoWjLfDNtyB2IROoNcX16L
MpO9re7xpYG6rxBNd7hB7zJur2Xy4lJ+BRsUgfzu5NVKsaYDKxDcgQ3TtwPOidrn1SkixmiN8G6n
VK3ncSFzDCFqwJwulVG9bOhbGU/SGFI8lcmSmPzm2dX6+Ns5DHGagDF6ud9zvF8iN7R8TsKmnXv0
dJ9pwclbiwuscsyNtOMx4BxdKJa8vd1Z8LIK41WkHGfAIzGPHoN/jyNJ1S9oGiGzP0q0UBQSP7TI
iC86hgWPbw73ucLLrV78+OrxQsmCZT7aQRtKR7tDWBWl/ko4G6Q273wfZVgPcg4OPwQnTqTWhPdR
dd8o71gBtsi+L7G7qlLGG3032SvPbFms193AhdJ1mwtS1d/yOeWqS1O5Czg4VNwBDtMYNf7FY1Bw
Eh/8DrXzMoH4jCEpd/7PHMMcD9oPxwwYd2wLhIoG7R5AKhrq9GsmVqcL0MjewYfI0kIzP4rVwYXR
prSsGd3wAyrxxosauQC09uqvesWEyth4+jDmbueyFUhV4zH4KcRNPPSziuPR6GhZS2KzBL8u9nfW
8AQYSyMdbuSscpkGVOnU7DYWbs5qA5S6c2IcDShLnukP/gyBoe/P6Zhb4PNASlziuf7B0rshVp3h
mfBVzqzDi/4BluT3co2WRiBwrmLCe2YqkGAAuG8+rJMicPTu29kcBQxOs6byJ8xvKBcGAHQm4FQU
+aLwUgtL7ihTWvQGnryXYqLmQ3NrkUHuk9ANK3log+w/KLLUF8oWzWv2Q9LXFA3tRzzQpLRW+BTS
lMaQrt3cNgmDLnt86qsMEqjI8gx1U8TPL/k5HhhTzZkJwmdpymkR8uJkfScjkMmyroFKtI6Wq1ly
SsCZ87u3VP2ODLyHMrImm2ztnSCZTVCoNDJOkk8cK14d0gOXbrv/G/GuoWuqoBO/8p8eKtDmo2ut
a6i51TqO9IJMoNCh7nhio8KGFK35XkJJcVNo6UXrIXx4Y5iz+nbteo+3gzeDmXAjytWI9NxT2y08
GckSkGciRvhoP9z5TLEWKyEdcOhD+opGgnioH42DCw4JB/WTurJB5gd1poRWMK9i6kLakNG5auYE
KYo+9VzdOSm7CHNx2XKj++QVUTkEgiN6VZ2PxoXmdQAU7z5+aEcX9SbNUjX+nct6ZnpfqONmZwzy
MX1X34ZfRSGe1siX+VRhv+g20qULlZb4m2A4LZ2FDMQ3qdDpBmqh3VkmdbMvaqHdDkirT1A2X38R
63xrUkbOhMcJaQq+OTYIQIyCzU3DX81GAz0NBoUAJNSpNVf3e9viS9LMhxdAiEsejJtdoSfafblK
OKzLV7kg8WbW4g+FoNUI81JrT8M2M9rrBLI81tss0gBvi0TbrypbpvF2MhBO7P6B+CTs/Fo0byfr
yphliLCW9TZtef9AgG9jYmRkHyq27lYLvAPGR5tMnYKUD9xRD7h/GYsFYDUhcMpmQq2NGfH4moXo
qQkDy5AB5flOS/QWNmWme1F9o7wqEX+vh+Zsl7t8CIufOeJTOOBVwC4Rjnb82CFgnAneFLjKyKJF
bl/VgktFjlTfFjgNM1nqt/DEyShyEJycF+jh0Q8LMNV2qr+zLUU2pGUSnxjpa7YgEdrJXIk+RbSm
c5CG3UPNyS+pqJkGvhpQOpsl08qBVoqcsNug9StCi9F8a6DnyBQgxcC0VQrQ0/8DLNjmSIHZVLYS
vOQNij+REDEo3RKXzhlheUr+fZlG6m/3pnTHdOXk0Wz8DS6ghNzW2NL6IG1tBAeNdXQmfuHeLJC7
P2bRSgZbiS2yQU2FBSrEdnucL09UWD9UwM1N7L2dTKQgyTIop6bo/QOQbeZCXSrX0ue6KUqJS+VN
2B27r3jPGpGTqHaYpnZfah46EA5VcM0FhS4C74Fn8q7zwhivhb/fLDFoUSwhjLSJrLsN3i3qsIVl
hq4zXEGDkIC2VbXKjtJuVixV57VJgUzCcG6QGN4ER9BZYflS0B+RT+WHuWSp8+LxeBtF+A1wjH6j
IFVWc7vPnZmONnXLTIHkriwUW+X/q640ukiqbz3tPLccWYpTm3qvEIT/6bQZr2n3ph9BmkGzLTnx
jFpvJ60xQRj81KixD5uvJpFaScDpZ7VdeLsansGndPng1ySLnEDljaFN2nqLeEb8X4mSGlONa6Ak
Cdnfc+Yy49gX+5DR7SEJD/BYwXlMppVMkswlP14I+1swJxQ6wJZXsnY23h99ayGEgD8R2bHqJcOh
ZNB/kF/gt2Ll7NMUyvgofWAig6++IotFj1OEc7/seheBY+6NhvsHXmyL8TI5gcW+iBekWGNG+v7e
fsX+V5aDrWBMZ2Gz70UZiJidfsLVANtzTSQg/niZIUb/LQmr41ze+MIoosIsttS8m2qEVjG5dxKY
RkrEjq7/EdJ14Bcm8eRFRhlqQcqb5SfmYtBdq58NhgLxLBXQ7qPM2OdeBh13nr6T7qmu7SQrQhHQ
rIQvadpm9Pehga0CSWxi/xCgaYDdMpeKkO53i8BAALCMue6G/joYObL6U4FinwOzsIWvY7hCM0TH
u1698WWBQrKXWC+gqqwrU9+hvhQWbNbJCErNyTZmaTkWixTeYeDWmwPruNDnn7F8cwvTYKFFa2ap
4Qa+7a8VLSwZvC3qkJV5WzYYJa+VobbvYWBUnoaXxRuQDnR/xHXTposqEp3my4FgPVmR50+mzLmO
SGE1EOyfGto3/9nq1jU/XSH/eYHcS1qJBcKchreaQGaFhFNNTo7h4VNPJbs+VVBvhTor36gF3hi+
wlG5XxZpvNULrANfp8EdPZApwJbVmyuYJEVO16CADsbGJzJYXpF35+f1aeKjxfvwO7lMVomJElV0
IXxYDpw+MA89zpweChRCsgf/XG30nDw/jjpcw0SdnaMPW7NSjB0d9UoabRn008dhk9/P2boRwdnK
XrcdO1XYilcm12a6tpPcK/17xr6MDo6fJWpeXqJ0L14yz4UcyW8xqy7miblWVoPJ10qbEmlWfejN
XWiIa/SrxskqrPbG+RVSDtYTaEbgp4h85wbZAggl81+XyVCPQaD7htrjsWQ1PsbpwsrvzTjtRnks
8KA+pjbr/TxIFQgx0YjpHbIr/I21xadCHwIbRMfW8TAs5ohf76KWuH9sYa88jlWxjX7ullfL1bN7
nmRqn6yAqXZ84u3cmYkkC4GVO403sTshDH00aMlo0B2WYFr6aNBf61wjp7h9LUZB7J9lSwMXINpI
msY9NG/N3rTz6D8dvYw+CL16uXnVLBbND6jWDLeXKsyLEslYaegQeDs3EPZq+HSG10mcVnbocyqe
+rtiNBzSz3WNKcLgqZQa1YLNBa0/r8j8qZvsQhPdrPGF2vjT31X1EUetZNxmvbnUVgoLy1JKnxTD
Sy342Atuibpg36bsxNvz9PDt0s6clb1Mxy5zYz3U7+VF3AjyldIB1EnCNukbKW22QtlVqr1QKn8L
mAFHgYjmHGdQNlfDR60oDPyzfYu5KKtDD9PvOw1ZP4iDm63KlBO0UYbNRVrSeqqu9e9u7QvUUOm0
SQ/yeNLDEkiPImasxC+5PURT7yaffVjCoLCpObDBh+QHoMwWJqJMYNrXmCZPOv11g4MhFm9bndKo
hOEFT3J4EoBP5d0/eVp/8YGJY9jEC6er3FFlmB+vMJo2QBia8/9c8gjiDbrPzt5usgxZNWm65aqk
s6lH7cC1W9OVTN5RySnegVNgs8sJ5dm8887fTxHSAcYRJppXjUOL4KBvD2ozkvS/vIPqjF1vSbqb
QhU0V/gGTqPo94y8voH/qRN8fUounEWJLt74RPfZkVxz1K0GUvQAzw/8Drr02GVHrumc4UYuVrpi
AGdLa6UGJrV/XXgLDp09mVBoglZ38EIC9ofAnZMaRHGHFZLn0mhMu3tHStzH7kfaxEook1TXARtr
n1/8zS6X3bApSWE9xBxNV1E0aBjOv/RIWk0HBu6iKR5U8O18o3UQupeRkIKAxMahiPNhuEt6Dyqd
dcQTUsqWMw4YvBuzyjQt+cFRrcPuFayVOs4pNvVyLZmGUM6+pmx0nzf95G4Q0MNYrasUX1FQ0pRD
QOFJIjFbazf/1FyfNFB13nj7PVB9bHnyvmlUhDCDb1eh77cfLint1iuL5dwZ17UBsVFmw5rYPWeC
yv+mhtI1Hpme0rCmJN/SPs3vOvssBxZdLOEXvnQnnpzBhv0P7SErMadHXfUXqJWLjiCqm3VpjoNn
6WAQg183Q1Mk/FGEjG5OXt7P2OomVNQHbCqOS3FLXzPU7HUAIzPpHEhyphz+6H3FtOf2jWDtbR3/
PDeTTT/YPjf83go+QRkt0I7A6PkGY3utOpWpWvxlW/XTPEsBryl3B3fyC32hQ2yGCsRVBmq7+EYR
v4pZF2ez0ctyCtJ+0UqxtxOloSyfiLtv138Tf1VCtNCd78+vrJ/OgHvNNAYOI4z2Z0VzE20vgQFY
ymxrg7TPl0p6NeN4eURaax9CYx1LpdkoGlvk/5i+m5kmfXG/3RGuswEonQlHnWHlC0d/UPjj1ufc
nIvxRPbQz0kx06q32f/B1hIftCv/1hlgE4lZGZmIhaMDq8l+EwDc2vZtD+ihVyliKtGRt4ZcKhgO
UAyFb/kL2QmOggXD+XfQ1ttJhPFNVb5kPT37tn9QzXFoKJsUoRvpVbmZ0319vxmNn9VRFy/9wUkr
pszWflWX/XYvdGkpFMlvVunPzTh4UA9SoX4eLl2hTV3s1gSeKbbbaI35nmB28zSEFtrbpqeGpREQ
adLrmcrbcCn58/hVWDzWMMBdwUo0D6z9FsfRrkbBEAkxg2jbvjA8h98+zMbVX/fnqeeMtNeVbK3o
ysiNcLkT4iZnN6bad/GjQ+fLQYkrbmSfXyGBSNeZZsgqklh16uk4yTl5Ovluks7Ow946jQnZE/Cu
FB4IpifQO+8sMtnMVtyo7kAVQ+CvWO8EkULZbI9rp0/mQli/eoqKiD3WtG5dawwv2vNqqVWuUpCM
gwkQy0Evn9u24sSc0DpEOdMXtY7QWB1y3qxmUp94J5oyg+V/7oGeTVId/eAprPAC5gm3Qqos3/Rr
+rJ8vUhBCw04wqZRGsVXnXQOPDBON0iBCovun42Mw+6FnjwRxCufCjSvHl39RNJtgQOXgUqLa7r+
PNqtQYHUJbXx46TCS7HC1+LEV71Fc8ZCCzpvQFgzGFlp+PX8KYSm9Ij74WQ6R8yKkun+bsJunAUj
uFGy7lWGCeX/zmfOoLy8jTlRYBx53NrURcuDHe8em0Ja5wI8FCr6K8E6lskBTgZlD7vYGFgH6vE9
vR0yYijbNe1TPK5+moi/l6wLb8YFKHxAkNtPWd1KagR0GkCnbuymRHWptC86MpfowE1ktsLsOUYZ
zwyJdatgWxrn7XJnbLm8s/1XRSnzjGWGn6Rtx4OclxtX0sZsjJ64mzsu5PpfvlGthicbBBpopWGo
rRsLeIzZUm3+zbW0fGnNcX3bXhRhIF5rmy0/KIko3gYXzXUAwFMvODCewq/kkj8qCAIOoQvvZg8W
2AX2zwVtaNwZOc02HDkZBuGxM7A7WFQJbXsW/I6JF0RRxJtgz9MTtoBOz5tiUmapYIU+3bEPkpet
YnXpPx0dKvhGxj0f+cReixsYy1D3HaeTOr7LDUvAKK63pYEvaIPFXByprM+gCeAAh+R4VR1FNBsN
9GwXDtBJ1y1F9XaNg1/dZAmXJAaDtC34mX3aZWZYdT1YP99mC0wme67sE40uqTb2oyrZERfmjvrR
GLAv58JKniOZSCTfIpU/a20jiZTf6TzhtnfEEezVichxJ6jfGfKt0V6Kz4vddIvXPXzr3K4XlvGu
VmWiSuaHTbq2ilgbtJVZa4Z/GSi4/ikLGcuhBP6IImba0JaAelixWHFn1iStLY3Iwg6xyPehZNcB
NCqSPdRqFywJ4RCOD68twbBDOcDOe15pzOEttpx0JlhDVZiwbXRzQ7XptZEtd/DbNIa7q3nGJBDW
pHXUvaaYWRiBYbiDFSBudkyo2ihVcHSzaYQ2zJ+Eir+ahErZzHF/j+RMoqzOBL9KfrOm86m9eBog
Cu5hArDN48GSB1Ye4X2l8dxDlHxEKxkgDC5r9AMT2nR7X/aXJnTVZya5bE2cdt7Xoz3tx0Ci4CHW
846bAjPaklnKh9fasuDw7tfT8MGypYawtWnB6hJfmP6tDav1HBGWN60rhmfyaa8y8jH0LwnDIy6q
Cno4kMh52NM9+3t6P43vPpR6D5IyQ3cXrIq3zfnRVS9yhZ+wfn8ccno7914ZWvjRiKrkZX2QvoWt
eRfJ/36XaKwMB12JJ8eyYCyz/fw2AMenakZIWg7PuHjrLZro16hMVv38SmwJ0iInTJPdV+8+tkVF
E8auqdmEUidRxC6qzyYVfaLcPnsiV98pgIO1yE2NYaamg+PL/bT92UBEhAFZYog6DT4zW8wRLqYR
96+hTkDmEWwlF7/o4VLprBt0JunTyWMYlqrwJhynMeYR9amR+kGePwNBstD1DnFI0xAGrWoT6ra7
ZLqQkYJ461Tq6gP45lcR82sMS2mnrYVIHBc0bwZx1WfBS0KrC2fEEvEL3GDZn4mrkGnyCVLW6n87
XdyHwQS6zmRhTcLXAK0tkngtS+0TrWNeB5cNXeziVN2xrRiZzx4KOlmavS7W3wslEQSGizCx+s76
T3TySGkGRZVOH2QTaA7KzgQxS0vePr8+0rJfiN4vppwABfELcwwbbsgR1CGec2zrm9x6JjYD3N/M
S2eM0zeVSJERe6RS9eM8W3Rk+rIUqC8KAZ/n8E+206t5HQNnPoNsW7pE9I1+S0oFAQuwl9r054cc
lW3NQy3bAR/vl3PBm0m6FASD39hW242Dfy4RV/jELEB6yPDVr/WDbmmIMkjgcjnj5baJzSfzB9m1
y/CSSdzjI+oOKgsuFG0K6yMARqoXS56jOys+BqQAGHg/rjgMQTKr5Cf3sBHU2fgav/CZLeS05KN+
EbhLxH821eBf/pX3FU/2AurGK+4E5lBphKMaaehD61Q5ki1eHS8Ze/ruskj/R+X+p4M7YCRWFyY5
X6CIJDAAT3e4WKHLYb7fgmGt9s27C3YPRKgpiH/MYRgJzFl5IYlpP/qTYLnR2i59YuHZWJo7p/7I
lqNJcBs5nVEkKskGiOMe8Oye6Xc23V96OqJaFxB7+UCRSkwnWp4dKLBvOOfu0uFuCFTNBr9GSSVa
fmI3BrlKo7Wph0tjWvV2CGY/5Ho5l6VKl6gJeEoisbqpBrLlUb6vaHhuTRBzHfoieZ4mChcTjO68
mCTm5NT0NinX/vea853YMvLvyvK0w79qqe+FlEh4Cfgy12W+a2BmJITyAusjDY3DndmRgHTrhZHc
oMw9+EjpI3QD+baB/nqwzYhsw54Z2oqtRoS54q4oFhKg+u/aJjbZq6/Qm9BgolLvbxmQW4kl6F0Y
bBuYaGyukLtQ4fywO9DHqI1Azol5ZGN0eNmMhL/htyfP1BtcGo3uc65kWO9Il8/LwVDQ217almey
YzQkxS+VDvjPGPQBRotWd+iH04NnSNjNeAj2mmPrUNkalKjWxK+WtJejjl7SOlrn5oMJi+/3gEhs
nhFNJDvvMxSeyfCdIyxTG8sxU664B9hblF1+MTrSStjyvEACTE752WOAFPmPXcZ0wW8ne+K8ZjHX
4lNzOcbANW22voIzEb4o2fUpWFOI1r9gC2NY1HyL4+ry5CVtq8mRwg9SERI5KQBvGdklWqftCEe1
p/67C0bOnhSrwPhLv5V9f7MrC/thB9ntGu4B5XksyHs7WtZgsR7IM8l4fFQ7t3eYMbe652aNGEyI
5I6MQNI6b7/RNQC28qT69ks1XmgbFEpxdqMmK2N/7DFehvxaAaxwHb474F3fvzQFiGXe4lpkKYhc
GGp2BMRYzNiAimFRS2YJEpxDhTjkCK6+7ZVwAXxzOqLP/Jc7rsks8bNj6PUOFHaTsZHzy9vKFLpp
79zEeLylxFXVAOiU6a2JpGdnJQ9aLDDJt0jDoajUXUV9CgxypRDDyO6aZK2Di5Af98WLUynN1Zua
12WO6Uoz1LCxJVVevwu94Zc4IRfMaQR0b0J4cyODv8kch0ADSW9215fxQca2LYq6CHwqCmPWPtKM
bPp1GQmyGGL9m9NDIs0hC/YL5bjdIp0pgLXQG/owB+svNx8VyaGHBZUJHKJ3qt03jCCAsb9Ca7Sr
REYBH7IV8mGDlCj0NwBkRol2X276mIj0vrV2eLgSWAU21SDcwtugiC/wU271Y5xy9kGRz5J+zO64
+XofwKLSa12fFIFEymbqKS/qYfSvEJCAmVWq+hKMEWVDXIYFF4Fr0RUeNEj5JXXATT8IZ8TdiFPd
++cdHoVhbTKYwj+ztfq+aRGmM2emSdz3gV2zVHtOOynEUxZiOhDldsiomH2jNjJsTDzNuHa8M/Jt
LYaykDuHCEqUSf76wxNw7U1fCvUrR82403aPic0RuxFYRq90l7+T310SX0UTOvG/4UtoCCnHEPfQ
0MMSXeo/qiYYFXFgrAjFCco3NYx+ivQMaBZD7iyn+9YL2MTJEub+4NwLZioBzrIVamlcSNqLfjR2
5jUPH0HQQFyaNe8wa1LYs6GGbxT6np5wHy+zJetJ2Vmqp4XLRawj6vhdm2ShjciP/8SH4JgU0yQS
/dyy/Hy8xwhP8pPN4y4r9udG3Tc9iiY64KQzfMlkSUg7OfHjVixDpSF19imvxBr3ul049GtWiNf9
QTKHnhc6LoU6XF6QmkRxS9Qm9QOkDUCLr0lfzFdLuVzel+N9iDbo7unpw9OVwo9TGFyTEqwicaON
OeAtE1yXQ9eCvRbCZhwFM+xucHO8Bf4cAk7K2JDhvh4Xw7HQle/Zb7XFG70K0jQQXxVHZV1RHzSS
gB3934fqML3YuGZRrEj1wdi+KY5C2Zi4ZZSBXiJFMjAEGq9/a7YYtOb9Be1Vw5vKZME6GOU2RM+W
jbs35FZa9KKC4fO+gOQ/J9BesytRZY7GHHl43V/OodHE9BzK/Ee1J7MlfrvcA0mMeCG3jVwTlv1U
5zhk4stASIOs3ITMbpVz9zowwP0awyu0RQmDTShRb/p9PFiPkmLs31p7QoMaeM5bGNDPvShxOcRs
YyRdjTaxwLf6b+Nt8VvWwh0V8c8Nh9qId5OqMgVefSGwb/0aeTALrIoc8E2rOIMIlqMJsoGooXps
KWcoq1e473yjUcZSjmNJ9zpUPV5AjTriIei/kTogW+C3XI9oJIXvL2Buljrcm68QUJb1J/RWwplQ
Y4F1+9+iwod+xyQgAuCU6i5cKKKUQzFOhqxTBC6G7l76iopAkPMwLByUG2LatUFSvLuQX7T27gMQ
k8/B8G/8kI3EoZcWBLRXHoEKtNMuQuMH+FYIQ614vdrahAwZIVLw25KZzXeI4nveIMSMlq3uqBIH
7bJNVqQyBvHyXcbN+9d2uI+x2VpiJ+QnOuB9YMzSzbAhtQm6FU/01lkmCtxhpMoxWj5SSxDsiyQD
Rehss3RpzY2UHzH5MXKBFJH9/DIydbo1Bk8D2XdeCePR4Sv8U4/ATlPDE5tDSjBgGpql5gnb0KNs
Wr5DFSNuNpNflqOUWD2RAgEI//oes2i06avwtmPl97qACi2qJQ01zBOfzKdu73+St4quHzX4ddeW
daFKQ4NRwMAzXulLf3mzl/vwJ1L2NO36JoqippanZI1gRTO6wvfTDZGCoPv/wCIPu8d4X55FaLy5
BsXFtBi3zmN38yN10Fw495uv4QKeKwcRI/GICKVxHdSvio0QbUjJDMLJK5/CTDKTVr+LzsSRZi1t
KtiJc1YaA7JfX/Xhyjxj58cekXGfH98BoRVvimlnXq3iHj4Jo/kltxbFEvsM9ugKFZaibgM60QrW
AS1MZmvzHTqcbEmZkRYlCg2OX2CsRVNGJh/z0SkXYayLZcEmh01mOawFJORJiCiIHD2frq1KopLF
ldeOq2awXGd7T0fAH5KpuSIlM0QFbW9rRhDKMprDw//7d+U8jurh23GPHGyOYcVuf83Qk8iU4pgU
2hLnQBmi4CW6LwV5Zxuzh86SDWj8qF40D1VwNdotbRqc5+hDPBs1nrAO/aKVLpQPcfJRFCc/yysA
94M2Id6w3G9mTL3ROBvktcCRVOYxGZpIKDH61ue5AASBUaN1i5D0YK/PRWqNo3C3F/ZDV9DT7CJ1
EL58g46m2z9DBdUZXmy6Ss9Fng6WSK2TnFMnJOrN2Mqd80A+JlJNrTbb+S33rus4V42z3TumnEGv
IBPrJadq4lIzJDXAmJ69VPYth39gpGm/QDTDpfFBtLPgmKW+83hY2iQtOlnqYMpaBnjeH7ZM8P3k
pGIUGFmnaRHhMXGHW02ZtIZU0LHPBx6K8+TKxhd8Rkesa2hehnGNHUmhrSdrTDQhLPvVkYcmxpwg
VxcHtGDhnx9Ac3MIi3kJ1hUb802ZGG1E1No1FSPDrVGXctOPNc8RXHYAvNVi8l3n0Cjg+mLgCHGs
4Spy6CYDUH827MKeeNGO4ncKD8zNRRyzUvN1Y9n40tblhi+IEyEunCVChvVwLyLPzMjKUHHNQFBa
wiyeCuRZFDE/XXaHtwnoXDq2XMyfRY7BtJuEPaE2ttKk7y801+DLrln8y7Z82Uy/KqOXeYbXMGDw
S6CrRwvcfN+dEwr+o68Nrfc9WgTK7DPA9tujNu+tpQWA9eD2vfxGgMVcx566+JqGkSUqkBv4FvvO
0GTagp7nmfs1UTYEW1P4bsjJ922QrpZdWf29Xwg9q8iqXSABxIBbrlPjQAzbdZtJZZQXGGCmsJRt
a/xbXaNQe9O/o6vblUtYgn5AzFpifEigKaw5uhiukZkltbE+exUi1LG7PKftuy3eHWQsdJu6CNnY
fEt+DmyfMAXOjiB0jty9KYPSaorc07AbpfM1R5guxGDbUsC2s/hAkbC08u/wWzicEQlVWdIYlQaW
bA9ADE16CLvDIFbx+jEzZ+P8GmrpPvi1gw+rI+m9zLs42doZWEIcuxRz6cGsmXc+jUqX+Sov2xRO
L2XtDSvi1Ujmk6Z+DoO4t2MBgZkzMU/qCyoqGvYFvbGw4hL02ioy+les986K8PKlAQkv1bS5GnJP
Nc3BD/lSbpJyS6WCD2MIsC/WH7GNTXfxLCt6mVfTcj9CVu4hpPbCxpiv7Q1xL4KcHShI7xHD1Lv2
EMb9dfH2tZFdAfpUHZB3cQVvH5/Q5l+FdjnOBKbBibj5BdKGFu6x9BW3QEOD0/SA72bnQBAGqxvx
CKcRpJLP7DHcjZC0t/fPNwkhUlEqFNF4fDgZyBft4brbmB0i1un8uJiCvA8iPRNT+9j6S5NoJESd
AzcSHmUIFvwJ4MQTog6MQPDXshglOe9K2AYn4zijxFvC++SBxDq613/vDaFYeoGn/GvuH8/s8+WS
UYzYoyRUao1enkHl8mVuxTrnjxENWXjX7DI7eWJtcGybk7NSCoAycPdwl4pMmM9m2ovGKAWFRg0a
7AjXDVrcnqrY8IFCGpG0w2nljtAuIkuXWck1Z1x2s8D626MHsaoe4A/LYWK97vPOWDm02QjBhD4N
qHrc2+mTj0++gqKK6i0SiMPQTxHlfiXYw2FJ2YeLD6ag1XvKU8JPHSt5oTAUj3h/y1FTqaf5vgo3
PxM9P/nBAx7JpT0fM2wwpHj4gh1B97BIcRCO2zRcBPooMw6v5J57vRJTrFdEglx4GfYXLokFrYrq
bIRIGeMhl3x2Awmn/V8uMvNfxvq/1Wd5YMgnvYvYm7jGvRsWX2zrGXXBgn0EWQxocECxrbcd4E64
WwIu5bdSk21fh6uE7n08o5lsnRybBFhFG8hszU3LpwV2na8Yp1vpv21K5MPGcmPEHbQHlPXC9NTU
rAbrr77hIKDpnm7wnPVKZ48i1+xxu38XD3ceZZb4YAsSCIs2GQkzAfLfnfLxHGW5VppdyslFMbS0
3X2b3G9Qqu9Kw7AyIYgjMJKyZi28mZ1oWwT0TW7Z4mHksrW3yKmOQN4+XTsRMmibe4syXn+zdFax
te2ngopfKyYshdNvwq8qb+PvslKkv8jh9nQ/RFcy4c3a/+Pbdh5dFAN54OhvLifw5h0lxuk4HuXM
1j/P6vJl2salLhM7syTaQOOsTdFLnQ3IyY1pJAkpyf24VrUX0fFWdBxfzYLO0iI76ovNmNsnZvUp
3rp+BYABZMm/Cafv1XVyaT/Tkxb01IBA5le8bugQbY7s6iAVU+DaJaQvwRBi372lIwjuIcBg4J7o
m4XTm/F5DWiTWXK4h0l7PbVjH5Q+da6IhtYiveE+lHiw+lqMjT01HSm6UtAHc/BbTEr+SaUQc0Vx
vmZCwU2zi/mngaLApwBNfxId/xmS+63CaRG6aUnZgknAzxYuhv28DQl6cJHfoOxyQFIyNtlPqElg
biWLVdmOHdtM+QVximfcs00rs+jmqXhs0+e4UdQ80LZGc7CMTvdwQkpc1mchgb76vLz+SLhlKaMd
x+HDAIsCIF8QhA7I8Qp6Yp60/J36Xa/PbFaaz33IYGo51OYU39vJQ8729OsDtCmYQkJYcAWgLCl3
3QM/5iwFvCPf9az3oQ5RcM/IkhTBxi9pfv7v9ezsNXmRpVLgbz3qWnrSvemNRbwhdie5ArP8JOB+
8TAQiSdlfBg96z0PKwQJBrRfo1WlaptwwAEk5z6nLqX+68ChjU439nePq5+FX8cw3GQYrKfjUHyC
TMBNX+P1S+5SICrsWSeGS08hIlmuLCLUUXmaKUG7YLQfMpcXqroFSy4Jnexlljfg3GaWuuJyLgc/
l/1xg1TEv6A11UDNvxwMLPHPAPYwd3oFJAHJlvKRvwg0iagoNDIXWZOGc9lxQAI3xh3QZ0fMZoKX
D/zbuck+jUSpm516HBTzGI26W8zJJMHXzxEnsAYNyhDs0Zhf0ez8onywYKca0Tg8bdICAMsNbGEj
Z2soqi8ZisakQzdch/ZTR+9zsTLe4sORCFShNjT0aZPHDCzUkyHxTdtVCFx/3dgatv/sUMTFiYFS
ofVEh1eYkXyQGqURkR1M5D4Z5bwjUboJsnf1zprFRSoho0F7/enbnBSLwUVskeJgxW2c+oGnsO73
z1eBl+g1rA9Z8vMXTrWtn4BVWZk75NkBDNWOGl3cD1cifvDeBKl9y7Enz0WRtyd8vyr2xH1nBKV7
5SxytP2jsFPQr64vWpT2mAXsSRzwuLTR9RasyZykflAhV7dscYV2jAv+wc9qRwbOanDUN5GpC52I
mgVQy2pH1UAKmcAvrqcWKqiVRW878V1k7ohNP7c+oOOjw/Z5pO5PHDnhl7xVvreO5SBPbzb1lZPm
VwS8Jes++xof/zzyhqhURkN+IamJNVdVQ8Wi1nx6CS2Ie/EdeLi5EmfpJviJcFn8ys/Wm2XJWr1r
+WaBauTpu74ONKUm/B3La2Pl5MK9BMs26H8rHSteI5yku3cs5++eGWlB/a4NfSFjL8mx7Co5IB71
bCaQ7hry2HrDgCSmxApd81XbHH3hyrAGBT+dUgqMCucAvpZ5i89Tfn6FGYFIIoHX5pVPWeKUfXw4
Gwfy78/1hJI65oqmw8itUS/0F/2MEYpPvQnQrS3uUWVNJxJrxzfwH8/cuuzeNvhI082+p9Vgnt64
ahlQKUwlxsKJhTRe4N8wnGGVka8RS14aEI3rt5bsy+LHzudG2KK6v6SW+/YvaRLiI9XLnqVeHM8t
WAPgkPw+zsSMuVkbatDACmlZwM57bvwU9oTrgXRsKhfMjan96PJEFNvL6lNLW5okis9+caBtNRzb
yc02UrQ0+tUvVi1CmcM0ThQ6mBvu0Y7OjnJPUhYuon1YegWUxw4BvV0gBO7rWGMRPASgYkgQYDIt
L7mdgdbTxAOJddnzL5/pqc6hiKeU+YH4j8RUAY2Q51ErCE7ne6tKRagzp0PaJN9rHk9ZUl3xsMyA
rhdT1X+EWxbp0CLvmjMtflUy/MBmyqtldXva1qVzHXdVmuaoW33A2eD0R9eWDWFkVLnc3A7i/PK/
DeT+YZh/BDNGwKrQN8QGSQzSnOOG09Yg3+2bgU5lwUbRDMpjcwQMjuMWiVdm87p1osiYrrkrWsLU
q0Nm6p0xEU0rlN2qmB9/sa24jQtGhDyEerBDPLCgnyLPvosUSTX9CKXUb2hF2JIvtkmzUfAd5yjL
xU6+eElB38Q1r0j0TSRdolyiok1ackE3jfrLttxb0LeTDBaNsykMgIDAJ6d6i6Qz32gOkI13OrUY
TMOvnsi33qc1tKBz6rcyfMaKMpx0GiQxXsMZq1SYlFeIDd2IS65lg+ok0gytHlVSfTp5UIlxK/kZ
6GZSeEjtbyTvl72zWURy0SsaDHhEuAAQY6WmE+0Gs7TJskCAKlwWYM9tqLZJbtzWdTk3umWAa8MY
KSOqOhX5tIZmafyE0wxqEyIyOWmmVTZxUu51zuJR7M1jVJuz5rzFuSqAeBeBYhcYuPsX5uGYeuNR
e2hWeV8L+GxU8YASXdaQfVH3HMJr7IRPt9DHJrb2/OqC4c/cUX7MLEBS9EevMvOcS9MPKvrwHf8t
R5Z3m/+rV10h5eLsrK6pxh6uqeS3TAcSd5OY8CHUMnPvA2Eowwv2sPbg3bZe2mZ8/HtVEUuFJSnS
wSQ1ztT3vVPa+uigjtaMf3st4ojVknHydqCukpDVZ0D7E/jbrwkGijxHeVFlf0nq0GZNRzc4OnD8
Sdd11/j2rcBlu5uE18jlorPtLIeO5077B1alQhrHBUiGzIL8dv1TjbbVRymJwqeMWf4t81o5c38L
CyJ6DbGuhIseyJTwLPltLCXNfYl2vRm9xfZFBJ5zPFH+YiVeAC+3rV+BLpETtCJiirkKX9Zm9v4j
JxE8yBh9V0TaVz3Pom4yQxphp9GDwqd+1uvom1/7wKRxbS6WCL4jzh8agwJ5wB9dDvzlu8hnHHqj
o7mLQjJayhAkOkxoBJWO00xBPQ2tYoPFR26qwYwMp+izlULoLdqpjeJYl7xWycG2bLX1Ssk9FWTQ
tz7ZKKlbynDyD26OVDS7V9z1olI8icUUVoiESBswByIF0ZM1Fw7qDWUa0d3Y3Lo6jaHpvhn88ap8
Ki6i9RMrelb6PA8NeUfbM9YOX6U2EdAT7FH2sy7B728097OFC1nGiJ5vy3aLOcUXwNrr6fv4j3Nb
ZRVWUCvg22l0Y8sMSklI+uIFeq2kCyu/b5Gtv+apVRK6aZC51tIWf4gQZdyujH7J9Slp8fpNFMWa
T7cr2eP1+LH1EXTHF5SNfDbP/spF87f37wZqDQB834VyDkO18h5RCXq7uiy6buz3dz5B3MNDCJFL
gb4fhxz4C8DsAZssrFnqo6/U6K7jQ8rx6PDYStl7q3+JvzVu+yti+8ZRnjAMJjnhcn6xGFjVBi+d
QEzUyHk9lL2ZEL6LFmVwWnNC+rYU1KwEni2Bw+FNFO+FhVbOWyAV2yD7dz+OdV/Vbp+0++v4RudX
4bNmzJbDvRCDWQmCRsKQDgOJ4N4wNXT+z9nxyu1bjjgiSDqa6eKVnKlE6I23qzp6kibg71z7Ny5w
UaQV/1u0oEzH6JQocweHtmId0TZ5L3D2jQIzzrgfRrhuEAY6TwS9HksEXluRJOK7pQmMUv5FGNXM
vDJjZEz2mhRf/ChptC0V5JIdJCGFw+886+UWLMSYphTt/ANU9fZLGbty6xzsViBm/Ch5bHj78Uja
z/Xc75omHAxX1hndi410ub2hQ0N2UF1ArvuN0ZFurNIW4DpQuK4T7af4qKJasSBwheTuVB+SOGTc
2jBXx4VvhWg3BqtQt2wCAozD6oH5+9cB7w75zxUdytfREi4f7zo7n4tSEv4eC2Xol8DTTwbd8Kat
TnBaA5jcIWz9kzR5Wm3JNaOLlknhvhj/tVxJeJTqN/G7plFkASKf1eVZkkXSjCG8jm0TtqEQRdN0
xokfPUpjNRjg/iEPpl6jn2lbGYRnAtJNDb+gm7yRY2KLIBDDJafb8QH5Ur5H/A1rIQmc8uW3IzAp
Jd2EhXpt1pl6TU2fXei9+KqffBYu+j3pda8EVVy5AXdQu0zrivNx6QLbvQ/IUgulJi2FlnKRlfS2
FGjszk7NehrWdE4YW5y7E0lKy564fXvPiNCIns8/ycg6Rtb81rB4IXxZkCyOGf+HnTQOBlZIGio+
hjxetDFJO/S5VWGOEqoZ60TV23DB3EAbqMOu/inH8wNGcXOIh8dUIRr+mIvNGhqmZbKBGG+rxNv7
fsXegOwRn/I7Yh2sVPATf0mHFlGLCYjBZFSS18uMUQFUuzJTNiV6dy+SMfFHG2YgYF4KEw0OqmA+
NM0ZaX/e0nC2BkR0J99yxUgk1DKhyFqLIsON+Vyzkkvu7VGFiKZaMKi9+m9ECTOPvNpQVjGGZSZ1
lsr2TbS7+iEoa2rGrTS6+71yFBQj0KMLIX4LKiPbRb+iaRF5tb9aI1jWVpnkZeHZdJJWrZuzLGkO
QwUo3nx6MtQZZNeOr35tuMFVRoCi+z/T302Q+UhnOijvH+jQRd+rYaQSFl8AcE0l64FhrszQ8Ktc
CA2HH0aIlEgq4w4fpXZhA4NLZVdEF6/bVrpTmOVHsJK4lKyN4RddQybP5+4YYRLnvda0HhU1UFDM
K5i3c26bSygddToKSqkyTQknVf6KaK3IpPFmU5j4wYDOlC6rHbqpYiu3tV0yoMNBxgh+gqPfRxda
FXk/0gcy56gRVT+Vjjh+2YsLEYtp8G+HHZ4Xl9BP22XzkBVpMy1p++P+TdTdBTTT9ya3BGExjVZ7
60GeTN5QZhohfXeuLVAIUc9pabsQmwDEUNls5ls2lANBvV040xbDvg2f9mQ2XOb0Pd84r2wFfI+s
pdR41VNFS+CDIxNOk+CnQnZzZ91FKHq2IsVZV9uwHjnvlSAkeapXvF8JsEGwwzy6ROXiQkyXqLJJ
lr+lPjC4xqBGsGnPYmEffbS/nkcbMDp1jX5aaCe/1BAs5QcTF35oqLD+fjJDOxRWVoBwoeFBysnO
Lq4MupDUotU9+fI1iRb16ooZNckwfkjx5a7zPK4FQ2yPepzCgvqGlTunwE82MeoFUJSfS/Yip8pU
qwqBE3HfKipMLngxEKDmhcP8iTeaS/QKM7Joyrr7JJbya3iXTSg7421vorqQ/dRW56v8WMvrBO7L
KVqXQtUqDgjNMpDDogQBlNwtGNGqBgu+TeqXaDf1zH3zsyB9Q3IxJV2jqJfQg+/JfBoN0CGkbeT3
+yl8C831bSj82d/IzWVntWCRZ8FkVZ1erOUUv3jmrq9Y4O7994Ohi08qVZyIO2Zgu1qmqwrLjoZK
Ttyv8ONLQxdI1UKkSOWpoleO71U3kHfOp+4jLXjTuQDvKAg0cYOauLBWjKXcuotFeagbggmW6U1R
+mI8VsAIH0hc71GSpfX4xmZTUSCF0Bldd8Oe/D16qya5OeiPH/uiJIO+qxEIuEzhlrYZAHdRnPyh
IYUzcy5KGlxWOP2fGRLWmCHPFBtL2immJkZyX3rw5A8hPQET5B2aLp4SFg/0MZ4vKOSVfsezyqOB
q4X4wOKK/kdo0pUn83bEaNkbQXVojgpGOgtpX4fmHzjbIYz7DjJm1h5HdI4By1NHe2GG9oE78K7Z
Ma5JJd4UxGBaa/FEUKeBXLdfQalSEu/PdwqHkfkx3oYYetN78nys84j/omOieMsCkJpmuIk9TmhN
wb1P078y4dFVQMvZra/EHk8dy7GsuGHnquH8M/4BECsf8k6Cvcehm49khd64a2i05Q4zQRok9g9z
K91dVTtno7xxYZYP31bpYgLbVZyIdY+VHYKM97ClBLtez9Tmztz8yCN6t5A1KvuhIKVnXAuRhlwM
k2tqdFe0/dTmejo6+/e6YthWRC92csQ0NcwMB9TiN1UvaApC/yfzle63L3UC+COJJ/VGU0G0tnPp
0J8rsR2fqDUdx5MLG8UI6rfn0f0IwF4SsjyfxRMj1I6tXcVswL+fwLL9Oev4QzVUefVzEBw0xFRZ
hwp7Sk2etCpCrdXRZaTme6tU/zHUoXCASkU/qN0YD5Bk/yaq8dUAb8KnDJ+7JOD3GckcQOAVMuls
7PiKzH7fW15N1ByrbLg2KT5h+FMQ9MvMFFq0VsdYoowhHZ9fn0F6B619FjaPU8IrKZl2FFo+yMCY
g9E4KkyCb4aiyGIm2IT2YiHWcXMZnA7HE7SmNXGg3sjubRzTUXTjvuXTP57DpGtZXiUAq2PIxLn6
G8YEF57MU2EGPn1n6itH2xSxDzGlihGyKZ1GT8iW7xExAiWkpFNPpDLr895vNCQSUuOUuiwnHvKJ
OykoxZLCMb/V8YV9iFa+krwiq697EGL2HTMrryAcR5Ky94ZD2Tf4+pYH0iIhQMPD5gvzp9NT0dn7
V88e1Q68nQUUHGHaLuePRBfgU0B+P4pEYY/C7skVFwiRTAskvG3qI/sO00r/m8r1bX2UDsXLWIMP
6RBqeLOY6SWiIXAfMWxytM/Vx3/bczH5Xr3CmqehSAlBwdS96y2UPBybCpLsputg7mhRMjd1qCLj
wwCijucVaC9jO/+QwXCnciXjrOgMiO+SMIMNFO+4vJX2Xx7H8Gi4iYFXKd/2ABarUrRF27RPNgV8
LfUVb0g1H5HaA1G/ve+uR33NwyuZuo4iyevNW0iB+2FaHRw/QYzaUqlb4GBeV8IPxO1uYikn6yRw
VFd0AUDxYobGf3fEFwdRxkpVrHbwXr3rZFk+5RBvaDRDkmCezj4THYwxXEtj6ifZgmnu8tXa0QRG
E6iJnq5Z8auLExjpuEAH8EhCVTbD6c8bLR/dQMf85kLMB6pGZxBR93IAgoz6qHrDQFQHY7zj7Yau
2VWlWlA1ClfXRwcxepKJMj29RfCDrRxxdaiNM03UDU3+epCCep1QjQvvIQttnhLKo2kK1UMdnqsy
1b5EXcST0pnbCSk8+chKa8cDTQ/Q72gPIZ0wdJS+xjQhk/3y6wb5YVhZVzP/iznstgnEVqt0X6NM
BrXoknYgsxslaCBIut5fH14WQBp2bfkxRUtHFiSyG62q8g8u4I90XuLvHyCnhnQ8Sq9oRLY7MNWn
VklQHliGCM64mCEqIQkvZUJcZLlSt/eWiAgXD2lXzAg+hq3L4IhXjr8kXZuhUBXdZMwL7U8FEWh3
/l+CwQ+XsDp3B4Bh1s/h0g3IDgV26MLuv08eSfDW/XO4cauagG6hr9P+gu+78DnUd4kLVKW4ef7b
59QtRYuojyUeYraV+6U6xcQd2ztzEG8ManYy3ssVUoTkYxJ5hb8JMwmRvs+2zYCaN8sgmYSUcc6n
E8GjFNtLHLl2YIYkHbyl4+zj78sGaXTVg33Smmj6cDdFQfQ1TcWMn6nyzALF9Mm2lr7JayZthGwM
9aI+wRyEjsyLo704yxVQnMDzcbddlNYcKF4pW6mbTB9nGwU4KSif0iS+F8ijcXyknZwyCIQdGRwa
m6yKtZlfiQODeYKkDoULKd46ubYrodHkE8L+CC83OvSRe3zeFbjcF8drWru8J2uN/J+xAfrk85kE
NUv+DfIm2y9DBVgFyt8PS8Jbys3CeCVGYPxjzSwSIAXE4quq77ScQN4A/YXUlU1uJJb+A2/PEBjB
VUbCTCnip2MoPI9t3oXyUN1bBcHoXVGPbZwTAnjiMw/W8WkEi2KVElTbE61kHDOqEk5UUmRUNZCY
Qkb+zES+i+YLt2fxOwdXe6KDnpUfJC3IJR0h+oAHiOZsr2MboalUL0oSOoH4WgKaODAVEwaVQsSd
54bVz6iM9eL5gJDE7wHc0lFRnvxmdpBdrjSACk949F8jAEWnKy9qfSxLmS174JPuo1+uKKbzG5wv
MP5EYBDLnQiyXkai8uwIdFNwAmv55MTy5Qd+1Dxj2uqZKiQzpFTz3ne2KUzW+FWjiG5+5kOas7QL
eb0+Wg6bKm+2Txs6emWYBJ1X4Ficld3qdadCi7F4gJ7XuLkyYRC9X/Z07aurOXBsazQqEUdPAueF
N1FdH8CeLW4vH/ft9QxjkcfFLJCiP4R/LBN7dhq898nybcinvrpvZSuPgJ2cThtR/qMzQEaRlq3l
mbGQf3j9CHb+A4+KH2ErHerj54xPW/LEKwZAYsS0GYjzMHoIOinVKjGuQBXq2PGmCh9o1Iq04llH
ESQxHALze/QzAyokpNt8ybkdjbPA7F0iR8OWw2hwDmyB+Wq2mF0H8erfRrz9/mY5fGv7nW2y7xiw
p4+dNaYRymL/OxrhHemuP2UjURd6zKBxVuS8k2YKHzSo9atLbSKrX7KmL9rAnPpSIb78aw8sOUob
reC3qKLRMrqV2t7KqI09UoopQ8rZ2lUyfwK5rbRy6JS/p1VAiZyA3pBcXFwvIRtVdP7QfdZSq8K7
z9NSzuNhrA4TXTk7jmNoEcUgDjUJiX7Zxj8PAHHymT2/ppJoDbkgFGUe5CO34SML+H3c6ngQGQBi
KfX6Zq4jwoRApsqVTwxB9GxYhc7rTMcMollAzrMfQQDkDpkiTz5+54ktrwjQzhSBUyhxyKM949ut
ButWy5GPjkbf/hQf3bDSwg/vl6bKn+p4/wxvzNbAaRiQi5eFnllK9Gmf5wvkHVze9nnP54jRkeWV
qqd5bdULB/YWP5FCwfywuaSl0Of5dNXEbjnQmOQi7Hrq24t1Ia2VCNtLWiUljxVTVoVjp92EAd8C
Di6kfH73fR7yrikfg2XpI5vh8EdpL9U8Rc217m6PnFpzX5mP2H/CYqbWOGPhY++SauU8++KzAd2Z
ywfv8UgmA48REBUJCGhkq29PgQIzTVLYjZj1HYAvmTjX/apl5Q2DejVMsCfOuN1BLrIZBHNinprf
WXc5L4U1whEAzAHvC+BJQceFmFm5aaIsLi8zop+lvbnuR246BI6daZeuAEOfI+XPyllJu+KV0Rgl
Jm8izMPDbC+Ru36pOIijeKF/UW/hmYRVGvRgTwJfB5tZpMWxJqNXPfBX+cIhrX8gFKlpJcwHEFm2
6cPJ9jvXvhZluOHgb9ZT1fEPD/IggG0notzPVS2cyo8LeA1MiAqp11RZwZzz3zTTTTTY7djK6rE5
KUZHht8Gw8wCVQOTeslxulsdQqbhYNdeGJtdnlw+ImzBa0vmTma/UKmmblfm4+8AWSA1ZC/qxG5A
TjfpZKkAGqL16/B9z3FYl1DPEC+fT2L/F2gM7giuu07qNoutVi0rR+3ydKxTyc9kkYZqb841cQQ4
QTpJ0bvoyGE71lCcdDqMBsYnOg6biqmYLN1uktN6nnkAMjnGjjByi/8qt84GdrnoW1qdkb4SM96/
D6CDUV2W3YlMXTRTJDJM/1yS6J89O7GEK6RRR7EiWZIOhsr9qsew5PKGDP3UHTQXnG5HnOT13mYV
8kyjAG8ZhPg0qV4XjfIa8p0jp9p1W7FSCC808ikEyKupS0zwAUmLPOGBANhorECmBXuAl6rWA6K0
UnD0qHOV3efRqCFbFiaGIIGaWsNvtZOkyQw7egY5oEQeHaBetPgmvvdM7/wcgS9uDr88H0OGzsYo
Q7j3kvYTA5xsW4wRCVDrw01yuh8EriJZnJQL93sG/WDLy3KDV6azn2IaLHUuUQdbabQyeSWGPcFt
ZQe38nvHgH86Lgfu01tS/7HGw8EUm2KzGeXURCi1f3pDtPabcKEsN0PCsSDZTM/djMqsgeg0Xeit
3WsAC2lS54HsA27m/9Iolq9lncSUPCsQfAKhT2gwySM9+X33sf3RYHCyMzAYIaUf42v27GHBEANR
kKThoiaKDtfY3z5SlXMVHHE85YQNf5nkIMRGpA8TbkRiSHCovGdoUF5zmsLJExclg9mHVJx442US
eQ77KSv2GE259OXZ31ki6BVwESSaTVbH6oZZ7CV32/DLmCeGPRKRk82Opdr+kvmyj6ScylFHC1pN
h2W2gfH7C4kvUWZHEkA7p3RS4CDwuhqBY0cVbEevOcQKdJZwXSqfTObxiAa2MCN86Roha0EusLuS
MZFzVDnPEouzmso7GjcsGgy8AtXzuHOEeJ460YfNxTVLXtVKLso+/+q4jwGIEWo7Bu23QXR7K5XM
0tPg8NiuJDPFb5AK+JTr5F5Qs+5YlLZYHSofUvx1I/0CmjecpQfsUhT9Hz7YecywgcNWfqOctBBg
NnpIeybNN9cOauv8lGh5IWuBVTPIcHBxIDNOj25Nvpdswudjfr5ZKOCA/1vBD7cb+GVP/G6qfj4i
q74QVg5QF0FPLWWSC7jRGlaCjjMS+EUyV5dJ/IuBK/oHUapnNwVc/SdNSIsZKuZbr3Le/Uomkjom
BX61fLuoPv+/WceDEu5KhZTw4kSX7S1y99Nw69A5+By7yhp9A3Dt2cTnwpjw7dg6qZ1hnErAktNS
zr37kX1x8eumpeZCHW6ldVzTR092H8oQmHvYTapckjRWKPhgMfIPsREQMK/4rILb9B7H4TqQaLFF
mSY8ontC4egx1jOmavVWGl4S/AUjRksVHV0EtztwfEP3lMY5T87050uZ65qkGBBwIcAl+WgTuySf
ntwu9Wr2B5uo8ytj8yNF6W7DF1Vz2pCyd1dEPsf1ZiPvO0H8nFVhAFQ4W2iCj2aVHJSydz3Fn0/l
qHSxZEKdup+v1wWDEj/o05L/5y0m9HHi2+L2Lu8M72TnlrVoaKG2eWhNVL/LQjddr6CugqwW2zBO
JdJSQWL9AvOANNQ/EKuOxzr7BpTz0ehexJZwIIoY3DfKkhX7yx6wOqcHdSOZFlKY9EbE0iSmIX5M
tYwWSyZYuLCsX48EwNtUAR5GdZct+iI4rsEOLECjlpfh8k3hiL0Y/NahP7UMPOAO5H8vrtBcSoDV
F/KK19L4VQl2+EyuuckiFjDI6UOlwXM7HRqrtu5zuFpbnK9+13nt6m44owU+UhFM3eiiZ3cTnX5e
UDoNX9Huu9DVd6O4QDy3LE/x1PYcCbZ7YT1wQp4uq/4RB5FBSIXlBn6JwJJ5ybokefYCA+g/OpX6
7oNasvmflg4SPeDKa9zCOwYmnVYvDnE7ANakuVJtVP0eLe0nf/qkw1LMRWXmKvwb5EI6kUgrmETe
xnFLnaZkM88EXWCIJ6dBD28GVSOERcEckIgG0KnAvePNyNzrqsZ9nBPAvJCS1l5kO3oL5PJdTn9y
Ln5Dy+HEG9ah5PIKLHQ4lzB+JdIXHdOkdwscmVHIWa/Zjw/Vn8m05MrOO9BjF12fdoNeMj00b6N+
2EfRXiBHs/319OHEobjxWyOTy7l0ORLITRP06U6hLRs+Wd4bRBjfO+xICl58KTC4JFhLatf7pniy
+gkMCdkeGxXs/i99evbvKnoUxpEI9S/NtQqANOF1XdI9F2sxcmOYl6HC3tJUCO1YDqMilIyfeAcd
sjbN5HcNNgdFNbVuZu3fFsHV+XPuT9uHdjzymmogzjdyH9V55pWH6CZbYh0y+LXVZsygNA4e+jLe
ofW2pxTA6saz499xx9FZ29qCL9xz/4XmqlVcV/vuMdUYOGZNO4M8W4MrCAKsM7CAkBBJRKi5NaEe
uNE9+wbSi5vJu4hMQI7AoV/x8HsBaqaNs0kmJLFL/MfbjnVddKologAwUAJ/3FwL79pv18KdOOmS
WsYtxGm37TyPWgy7EmsgrSXQ0dCehz1+chDTzcX6Dtblc3P7+mozAcIcYH9BIorzwq+XdxRCKSIv
rF1IDa+3TFjjA3cab7+dbb3eLGZrM2iEYjvJLIsgT3TelhCK8mLj6hnK8p5AMIN+b+Hc+aFVo3Ue
MoLcT6mAglobAHe3+y1gJDlfD8ak1VSulyD7hRUwVaXZWAHAawJ10jr6OO4E/IPPO5B7EUz7ysgN
bdHX2eQOf+i5rG/REc6wYOqK51yOH7lLDk9BuNd0QzwbVNdxkighYnzzh/RtaPXbCzRT9to5LGpR
ciCJ1XQzMdwbR1borak2VrRjRXMJAGaREEVYemCxSQcE4jKFYrPb/Oum9kmXUot0/xV3w03a9Qt6
Fz2pnkCI3K7CWa9HlFvj61J4U38pT5Nk9ks0tqEMHdp6V47Dv/l9z/zi0EmoaFozaFFVydC5IhXN
uDbXHPzpHktcEkSFcbavdkXr7Yxdaq8TLbHR3UKpHMJgw5SwTQ5ezp66BHGaUFx1cwZyxWbJyqCC
gcc0iYrjf9HSm5gfYMUhL1NV7o+sp700IGr4aGIQGIJ/QQ4OFYkfpF5CtChZXIeovYafL+8XSW0j
CZ/v3UOsj1LHX1G40LiyjkBDWV57dsmShUJVfQpcfWR8RLmHhqmFrZHW25VCaC0ydGHGEFIcSIY6
3qhDTprlRTSFW0hNziMRzAjHM2BPdeqLY/evtfiijJKhEMei1YpixieF/Lk37VUmReXn37aBk/vh
o8Bo7mjErMrCzo6H7eSrkse3CDIbD6pj/MIe7bFI4q2avYV7BDR2N6X7E/JxN+zLV4TPskEYXDAK
dnkLwzk6izMSk0n99wnpUdIOC8OOWSoCeB2gPRxBlQau6NkhspkK7jVBHOk9dxEUrhr6ArVcowGo
GWY5elTCnWhHkUpXb76NMWKB2hFKG6DE0YVuGtF+9MxD/jt1uxR9nxYMrDfIGQdCDMG7imUNRe7d
C+1amOBXbqiWRS/arT+d+yTkdSHCa0Z71Bz/Abx4RCsoAJgcc0vVHgZXQPrTCa2lVBClFmRKMwBk
wu74R6Qcf9jbgZR3IzGe4A+Eox+55qljuY+95qKoomX7EecFTez2kcFfqUicXzmyx67PafNs9/w5
S+itHNfxMTVZgYF6Ynx+E/7oTqM5spee9F/k4k0yxT21WYoGEA+fg+ZfyrCFsA8+GsCsrDir5Y07
Bq2cTPM1dB3h5+W6nsi47Yanl8Bn5CwsGCM4wmA2/PY8Q2zVWjPLwA2FYzST8Pu4CAZ8mI9sOrpj
Ujj/baJJfPP1+bu9bMNE5l2GboVs87C8yqZmbGOaMpdVqeIe6GAOA1Oqj0Y/ZYjMTO7CCD1O2ZW9
Y2YuppumvngSWwCsWHi9QBfDPgvWU70M5UaFJW7iaQTYv9d4756ptUy/aJkCFk3XYuKxnY8GmcK7
JuKrx6d1GaPfhnZkEEzx5BfCB4qf8vgeqQr1LooVsqNbEyXRx9ypRG4q9vcZWJxSxr0zwtz+sWSh
Iq6U/xA7Ucn7rkRoxz37baoTKSi52jZZS4E9s7AGORmBRHt+CWciggZz7ccyrptOdvzeMIUGSfkv
z62pMqp45/IFQ3s/fSxwum65vD+dgoCU3g9/V+78dBEOJr6n4KniMiBIyY12toVqC3w+99owFup1
JiNzSS5AidqQ+vSRINMWp1pLglGtnxTNrst7hX0+9Kc7Kg74Qj26n2axfmPu0kHL4S4gLhqmKdAA
wH5XLyqz3BN41TljBRR3y5O8gqSp+H7wfNuowqkLehyzDb2K3im1N+iB88NmmIEF6eBSPKe/i4+/
ya2zqYtRre8CxuseFOMlvr7Hdm/Y1lb+lbIPmPZfLv2wCkJZcP48d9hIjB1bi1aRy0OXG502+ECO
NDLMZPAzPWkf6YvSGv3cAiiQz76ouhNGkKZ5Sv82kRSI/8BjtitUDmf/t2Ik/Qsa3Xk0rgCt3eDs
HjyskCIwbcmFJxMAnB58G3uGyiK3oycupVH0MioSFGCiuc0l5A6TLVoYo0N5qM54ztlwathcFNAm
K7Hec//9lEVJAEVVUSuS0giG5O/hhj7fziGikdcL8KMXvmcRbjd/ILRoazEJsYfPfqyU0Jb77o0v
AnJHXzBdD3qnT62kaiM2N1hCHCPA2yi+0SulEqd+9sZMfTTvS1n/6WpjRCQmyTSY1x7dvZqbpJ6w
3Wc8yT4kCfHxgy0wjdPFwtWlVAmADYZGKHDFkEhKSDumOPXlRYoHN53qa36Ek6jYF1rBM+P5Um28
/sk7XnDvcbEJv6F7vsO9WO9JAdjh9LdXggOWUVHCHdiN17rxO6922ugGeMDpYL4mC+IWHVn8aIIg
UIZIEqOdRK1pZ/kl59YY4bk6s4hjQmPE8NkK+ET04evxJvxoWq3KUO9g3VDmN9AUye7F0W67MsN5
BtaDw6Pw5SmxeWAlMq6KISYgoR0MPARogyEk4TfjvuSfI56aLnt6LKI4wmD7XIiWwAGEXoXY5uiG
2CasdKUsAdZU/lHJnQPOYkxwCoVNO9Nr01GYYiyTmEUH0EZyYNlJtEM65Q09IXLxsHVdeTCVi+vP
oMlIUKhbOodlb6pWC3SeYPOLtDg22EQBQeVbRvmAj+T4aP4wWz+Xa5a2hwk+/WC8/3bBSHQSvut+
4M/Bf+vgrjnStm8QYCHjlAyYfbN4TWZs3JgRmDnVkfBM92GRynnxKT8IbkzVRsXAAl/22cdCtwze
Nie7PJtrfvZ+PnzbE8c+oXbS9jQzGNHPQIdnEHfDQZxBySV6cbxJ4/FE22dSKEuTJexCF6rec+G5
8NV1avc7oC7sLWX8//ycdXUSfHsOwMvSeN04tRxxDcT+KzD4MJmC94wMvVRbfVfdvkQcOraRX//j
/GBajaA5ReVswCpgILXX/jGY0CY6rZZfWAGn9ajMOTfv0APVfkZbBDM8P1DFI7YSHFzZtvyv2zNA
Uo1QjvdTMfhmUFKsJIo3G7VwgTG5lHlEf0MCWZBIuP5kTTX0g1mJAs8dG0ynrl5V/P0SjNKS30Xs
TY8K3m9tYsabMSt9/K1xWYbwBvTQMetnMQ2Yl3GKTPmoUyS43Aowo756q0VG2mbD3K+nv3ikJPR6
q77HNshwzs2SYALcaj00vi4N26DRgDA8HaXtkJyJyktNO3qQ7RRfM5hHUFihkwYVZrrcDZNymShL
Lrg06KnIF6X+Om1RujxgScVTVVEeRm7vB/9twPW7roxoreWcsPxUUKNVh+ARj01yZGCu7TEhhO3Q
Svh0t9HJS9fpfrnvlsZsP/XXqv9zuPIdA48L+otrAAVbcMrr2Lx6rV4t6R6E9C+vpJkGXs97V5E4
fJLzky4JdHOHYrAfYamsm98An2Za0JIUEOvAmRlX/3uEARb4qRDWUWHPHDwfvau/GRjOMtx4vHwM
vIm2PDfxzmwRJ818uofdFdVm09vtw6jq+7pDVvIldsoijOtdWgb2Q3ZykdogadyN8lBHOUkV0EAX
ROvPSS5eIPaEqFb4QOFz0SS/tCfRaFtSDcW+/2tqtUbyAXFJ/Hw2lc9vnaaERM8ggMaFBuOQDGfe
y5bQxw3AXdkv9XGXYqgXz0DAcaxYwc3IwIpSGUpSM4hNtbQEvMJ2HGxpmQemtyxzrnO+fxG4HmBT
dy8MfY8IuYP1X+YsJlXyMvJuyDc8fHp3c2fnMio1lZbCsVxMgrFY9TtRuCozOx492VYjWn91cy+6
UD5Zkc1HIaj7+VHzeCb/kLmnahsPfc95QUHfEwTb9SEqwc8T7TK87MTvrLIn1q/hLMv0dSklofoN
apV4V8O1lff930aA6zWfpEg9d+2ntRYCcrnvG866b1kNGoRpLa73bPvqXg2Cibz1mVi/Tk26KNUT
PQGj7i1ye55cC+Gl7+AVqvyKAIIwpEom7QwFn1RczQFFez+RBZ0mSRe9sJtQPqTAtJOFnBAPZ8yA
Xi7CdBNSyCMf7OsSlfEm29H0vZ+QqxtImKUr/WIW/Ni4adFmCYMyl8o7E+mBHjdZr2czjI7iVo2U
RybIuftLj8Fe39HOiw/+DX9KOjGkX6qPDTd4/VkxA9syZiF09tOQMgVuYtnJZa6K32VDut5YJgFV
NY5ItjAqFv+p3NqAk1bHEHpQPXaawEuNJFeTJMaH49kgLfmYgtyNV/eU4esiFkGYiQbR5xVun8RB
ExCltcsTQR2k6Bq/BNtVsNdxJBErvo/BPwSbi8sAjkYy4uDbpIGup5W/P5pJqwOwyE8LaiNCkcoR
/eywJWgSOnqoTswzqwTBveF4384yar4INdItS/r/PzijNGh7n6UuefSfAx+7YEJOa8GCrapwiCTK
+io9buYxrS7Df0axKh1L8dUuEfzb3Yfz/+0wEAvwtfwJEDnlcVkqQeKXq1Lr+RNn9UYljhPvJtXZ
o7he577NVfQk9LkDgWo4+eo07YrxSXYg1d9ao4MPvmAvDBF+6mPbmcb3tgvV89uaZoYeWnJ3Zyca
y/n7LxjTAHgktyrm6/MkEo2CGILy0pKTFd1EI/BksaVJ+DffHtC1oRMeECY+8DZkXl6NAi33FGug
qvSAPelGYJt1snIgZ86I905m6GatpeU7HLdCwHuLMtYdlqRdnPgqpRFpNids8XFAeY9YhwFA1gv1
CqpYYsXUcJ8+xoyqtnNyWOSre22TNGgqJs1uFLVrbK+aXxNhw3Dy+o4nNI2pyD985DHlmSnWF9s6
blPiMRSSGRdTNotFth87NJQj/7PYHGbrKVz/ZolaNi+hhjR063gUcQFQa9kGTQkeWzgfTg/EOiBy
89sliSU+qbYY7nPHYBym5DgzOFaf5XfXHWcZMABn9epHhhNL4Mb6GlD1m3HEqRGXmKZGcbIu5m8A
wTqToTmYVtFBHjx0dnmaBZ2wd8FsJWaUgA/aiG0+c5YI7Z4ucpFutfwJJ7vqK2shov2PKl5gyejV
+f66/3GnK8Z2JvhFXimgY2vhiOhfbWDlg3ED5CigGhjqbXDKoOYCgs+nd/gtFFX7C23UAHAcESab
zogvkvZ1eghCzyDHoot1wxu/JynNb8gxXG8RBCuG67A1R7doEgLCfOOgf62cTFacu9hIfvqxlcI2
uT6cJROvjB4KqyES7s83ID27Z5ho4XWnLq83BbDGTHlbWtT7+2qwd00BRA4mYru5HM2JJ94tgfjv
b6v55e9R7bdIV28KBhguy21O7/AhtkyT5AJea+w6ZU8iMJJNHek5hsR4Ro3dZfYolHhhQg+gaxR7
7c1b5BKU7ZwkafLo+o9XOjItLf3HOe5IjqEbXJ+BoJWSj5Cj8O4wXR6Tdzyrm6nZonZ91eoOZMRa
eFhmR+ygFku2xqeI3bbO2Qq2AD5ROijd2/P4G7MljTCAbyYNV27YRtNjYexD7yIhPMa1nZVUNfJq
/ZONUnBk4kMQ0pHGIQnZz+kKKciLTF6mUyAUfOshiAxx0TsXxYV7KIOt1sC3525pmEapVwtb1rgt
FPG57BHS7uHXx5CjiEAaeMck0bh/aFN3dN3TUMQsgTz/u0Nm1oM9oyududbMWSihwl5rKZ5I/RqG
evMo0nGqdCcTutVaw/aTnQJFo7ZT2zHMJ0LsHC9mOLdRwRdrMUEfZuI0uPO+t0W9UaQUsNG+bXsl
cfY7ivRI/Nevsbh5qUftuWdxmNiiUNxVlm5wUfA95ihlSZmKZn7tBhbHbW5ZcRuxjsCOg7H359KL
qBPtaaqrh6vEipdAxMLYQqPBCOL2ZiDtwfHLDN41XAjA7mz2fCJM/R9ur9u0Qj7CrWTrHT/YNz0B
5QvnCTxjycV0BPQ0lBSCTPaPF+Vlres2aLllB5HK4xz2V7PZKCV/aIKNjzAqEpP/r3RjZwAWrUNt
l7Z/g04r90I73cDbI883kJ6LWQLPewz5eAcaH59TvaleuSCnkU+EwDO+ZEKUec87aY/IrPjDo5IC
cSsANE9rgpVSOMWRb9kUPq1jEEmpPpMtneXYYl20DqOHXdlVnHufU/3+PQGE0X9FSA+KX6w1eG8E
+Lf+6MKdA/RMXcJArsk1hhfUFtST7VloKCoaxwlxDa1Otbb/NcF6/SeLcW8P04pqZV7ger2RSFf4
50f/gYDSBKvW/dLCrEb2Mei72ugUKRSwXHv/1W3PBuiBjk1JeY/3Ju8538LqgQ/LF5qQBS5Z+Q7/
YCc9IGUZtYMY3EO9AFwpfpcTmSRBrIEiP/wQuTe7RPUA0msEFsiFcbNM7h0S9KqF5qow2t5hPdcp
aKrpHa1HHtIFyXBymBlrxrC5wXqgf/G/yK7jChJJkTDq2k6v05v91pFRSYx19q1eOElgev3Sa8VO
wx+FGrJOkeR+Bg+FGndVRd+qLVJx/X1NxAXWDdMlAnJRy7hHRzDBFCIgkYzQDGRCGNsX0TDNh6p4
fBMgYGGxc1YlNuak0RG1rwJhGC2hfJEQ/M00YOOCKq7LrpTtB1cuChECeQq/RMVF3uhZSwiMGRpM
/fc/lHtqTjaBejdVLjHps0WoEGb86uUut2rjmb4ODGGR0REmnJPvt2fpwJQGTkElhpZGjanvYAmQ
rLSNBJYisWTj1kkkqdZprjOwM52cLIZ6HEEnqaW/nc3lxUNa1Hu1X+5raMWIavWmdnfLZSxS00gh
11GGnUbFUv7A84cnMTDTBChBilCHOsGhosHZ2RgU7Fsl3ecDQe3CCC0idOz0b6zb+/ve226mgcpL
zFVtnnisYRcqMrCJE74Xi9lz9o8qayJDdmeEexDKtvUYY84ydH3INCy3v4jFbPNaz2mYA7LRuS7k
/KwuBjMCO2ZIgzgx/44pGuJfcWMuBWcBwg61xLnWZuWHwzqHsW+qx100pmNJFkmFih+MzKsG8xVQ
MzxaX6YepDJn4zyd/ZwtGvnH2qbDqxp+me1dowrTQcwSrgGF/+fBqkcqNQ++zFh8DxCjVK+xnKen
33k5L0el0IwUkg2uyQXtSbWCjhutdDonMimSEOl3FiOOv1wBk7JtaYS7cxCGepsnTcKFCdtdn4gU
uaUUuYvPW2j2NRMMpX+B5mp4xFROP72hxrVHvAsoRU1c7W+rDLtRkDKFmmKNcTEbEpb8j7Tcbg2M
rZA3z0w+NCh5bJw3zxbA2lkTsyTSYmOIfHCwwMiaKMTYBNp4VSvXx5H6LKpMSYP+6pPXEHrPDQIh
NjwgukAYT7wOTQZrV5wC4UNZzRsPVzHKqClmw9MSXiO2Yo63T4550wlKkUZqnZ5LqId/VQkouSzA
vJ/N5hnuzuttJ6ip28yvpDdquZ6UXc8bfWSVOhVTXbs1xxct97x/YImKLNNg0xfcRgP3qOQ5PAkc
aIGuuOGe3I6GlR4863J3B0DDbwKgJqgCryNfgefdscgbSjNnh/e33VO7pWnx7Lcj7pUo1cbAb/P2
vv2ZZEkQbETdw2y2kmbAaHOwRX5Z4CTazaELU7RlfxZidGO2tyL/VHDfqkmR6KRkKTe4h25zZpzT
/qakOOXhrTVjdEeem3G8QJm1C5FDsaMOS2QTd6M0GGGTWgkxMpbtOZrcmTNS1OjQvRkol6tKRTFZ
pwgWmPYaFCQD4PDipBL52PsmDPslBSHShdYzTxvG3x7qBpO0nAcTLBwFo+Aj+mE2LSW3S/jp5i1U
cqohCJc+eY4PZrpOUTJAgL2NA3Sqizt9PQS5x9WtkpOo/Y3XZwspEQbGy2jSQx4o2cDL7NeyMJxf
HIlAHMHWtVhPzpUI1EO9BRkXmCfPTXVDty4grSUU1Jr/jJS4AmSTyGaX/Tyw8xc5M07sbrOAlyU/
oQYVVCpNB37d7Nm8PFDib5ZSM+I5UdvOycNqBKomg3BVAiXBkAOij/nJiyg+xFFseI6YYPNyAKZy
FdwMihwANRR5pZxXiqo7auuI5HL9nncUlBS06M7mCoZ4zObsubZvTRajlAoqEmocXgBEkuzSTW1V
IPIGpaNBynSdpjnlYPj9FC3XKJ0IP6lJblXTYw/Zt/4HDbzd1XVfbppuyCYauZg3jHi60459amCH
MzXjgioMLis/7juIIsrhJL/bwlEM+YEcgJbyq2xWE2Lnk5rj6OU5lNm03qdbouidhYT8K7sZx/hy
LVz8uVQ34FLLMA1a4+x2K5MbIKXl86fQNz6jElXGHhwUhQOC3+lMnQMdTdd1wpPahfcTMfuheui2
38uNHr5kRw7zTb6pB0VbGivqcE4EjygPtPZCL7/mwjZ8R+RDNMz2bx56YEKB8hMjBJXsrpw6wKzj
aJq2MtL4v06BGryaaEbuCxCFCSjg1U8+1H/+1ykg8jmq1l7eyJGr+MFE8pihWp97+OEZu/84K9IK
+bDVnvJniRrnogYlP6TOAXg0RAdsenuR/OlO+JbNW6WVObJKmYpZvrPeXlpV1StIW2uR5MTzD56e
UKY9tSFhIOXblcc+pG+04lEBrZIoGmH2yrLbNxlqCExegRzt/X7KfYGz4O0C7eZuDq7OO7YJRNcc
Jg0C9S+kkkhh7r8mW/HiRXUmIGB9rwuVnmjs/WurBsgDeI9wUnoFGTQluZow+r+27y46hZSjtq10
THvomgFuUSvEbyOeVgHZqrmXBAmfKJ1uwUZsC369o5eqomuCxIFS1rICiV6qy4Nvu1sHWRATRWFQ
bWXVda7vSxS66OJESlR8Y5blEv1Z0QGuWXkryuukK9qy/rA+PRaRB6Vcv2C8wXVPN2l6HYUgo9N1
YWIBXMKzzkzyobExQ+HUdh60BksFb2tfPK3siXtFsI9hroQhKMZk/isBtnfLBL/gF9xwImSeYcCI
ziWIk61XJ2j8eclgG26/Bwx7pLG0ajzbccneXkvhphgRJ/7sr4m4D9nDqSYcUImCnle7L0BcALe7
V4+yJjyfRYgJDsOrucK/PKAjCSSKqbFYDxOQsOa7SFC3WVpdbZ2Ethd9g8dTo7jUBLyX4TximajX
9jIlggjvd/brUOg2X5JRx1CPyEufzgHU5Wtc7+2+HmHC3Ki8QFmFJ4TtbJRymz3id/DU8brc979T
eCJfiTOaNI4NnKv6z9UzD6OVbUxuCe+7QjSR6IjENQ+e7gKHovDADP8hSaM1omIOPJCNHEPbObhV
0bMPPRgrFfkUK3CIhGkq56Dwufrz2x3qSp6mdS5Rar9L80nqRrTa83coeXkhxHdirZQGoU0mDzdF
ZhycErA7sVKl586gNv+1xauADdpTslrDSrHbX5GA/dizMdNSn/FhKGCXlx6Z7vPqja68NBvtbm5Q
AGGh3boNB5DZ+YZ2kZaEZbpLEtLOTOVP1XitFH4DdsbUgzQpzQgXbpTM5jn/D8J/FIh7lLgQW87D
f82U1ChbDr+JbvrqS+L0FQVLtY2Qr4GSH/4fY0vvJ3QjnxmaCiWlJuy04KgpNCu5OzgAEDrscfRt
JEtatiu0pu+dk36Fnyym8AzwrB40vraQ0/UTfByshyKxfhKOJKeifvh8ahIcbnq3WdzAWiaCEOqX
nH3I7FgEl8wRm4x347xB6CBR9lDGrj7FxKOmqzcjqdHJta7k1xHy5/15DxSh17i3eRZdpzZi7NZX
4IvXVcmYiwjHgUabzURn+PJDaPVo/Uxxw7fgJ+T+cNq3c+rOgj2TD8wexKub99R8wVp1p+Bq1L//
5SyrzkuyIzkO78b9j/5qi0457yFCD4OBujSWuF8ZMJAI9EfroYkCQL120xq67GosE3bDrPCoVI7Z
flbB33tC2n3oU+s9Gu4xIVJmlKDMCUgqAPJ7I1PgzH1OfIS8yAD4hBfG4lgER6t3DOQMcY5Y0bLE
boz9RtMEPHEO051uMBt7Zno9StjcCmFsWh85pQ03QjygsDDytIrkax6YUU4akiQIj41SMYkb8Is9
1Dp1x/sxuLpxw/tNZoKaA4nblkzbA1hNXTRh06qMQBWuNNuWbvDQ5MLSYeKzSi5nu134zGXl2s9u
sLrvh/6CvwlaIFclxt2u/mqqIgvfiKeB+r9HV+//Bw8S+z1QcmPmhXqM1bsyNpkpj9IP4F24NIHB
ZaQN9AVpRfWA+/Xv6NUdUOjeG7/Fhfhcw2svKE4gryY94XBJ9mFLXybrWIuFAXwW0jUnDd7w63Au
/LS4F1y4iFWKoRuxI7kpsi05fmNJw+SuhL2VouCjw4TAtkPNe1K8MRZmjXnAWCIqYBK3Cp/ZkB3v
fpxwKVeuG6DbQGmLJkGoJVOTdLT8BxQ4/fmMKFp9JLJnnIQT7hOqxUJRSZI5YCfGmfCn/h+UvQNG
HmurcgPNUvHu9UYV3/wDNYHrJUfrBErM9+OnhgsbTAT4Wf2EaXZ8k8CQ1QrPrVBHV6KY/h5wazKd
CXlVXjbu8zT17shSRUo5PGO0A+jC+2WgvWr70pZCB52MB+9TMmrh/MlohHdZHfThuGPxqzFxxoxa
XBMovWLsnqRoJB+4s2KXHGJqvn0ZZ5Xfod+H9AE98s6RgJq6r2cS9Lc3c3yl/xHJo8EpOJdZAeld
bCTBjdSB8nQzie58Q4LvhyWqlvuC6O4Z0VvEmrwKAY4IdONKD6DTpxenJKBpBYwX5DM1m8WPxTWu
0sFsk6NxzTkNp1XRs0BNXQEHjTpX//+KwW3+bNZdEEsjbXd52Oxb9cbLRDl81zJeWs2NVRkMI/bc
FVI1GO2NMA9b46//htYX+5UGh/HApNoM1zvPhDM8vhXTwcjGXH/tk2ZRw5qKVep8P8XZzUY8EI6z
AF5qVP/9wWWxGvF1ZODPZKFkmOuNpG3vgJjpGq8EZ4xGBdShtdkIFwkFZAZI5VzvFydp5h+iHZ6O
FmxV5TuNMKxYiJwm+C7nPunkLJBJF7XIn2ApidUgeaMBPfT1R7WB84a0WN1iMq62n2w3nTVPB1hf
3l4xQHAmlczKOunIzfFMUv7qy7SD0xfyrFIrvUPgV18KEBwLOu10yVQJoaIMZvxOFMJADdS53jXk
BXely2bn5onkDSV4fUJ2iGnUNz3E4uAhLDexVCi6r1sT/axI5nhRpKQksN8aITPjNYZXQi0QLeOk
/u+0KF1sQX1OhJLJwCezgL1T3X1hW4JuDubmWybOZedpKj8KzV07YwIVDfhub6fMrjed0Tlbw5cj
KdgUQFBlmKmAsbI+VqD/rSHhueXa/5HiMCZHRyheINVwAj6R0xf2BafvBj00JtwrRjyw5ujBLzuW
/TnbhygfFGTPyegI56MTaTExUuf7Thxt24T1/4RD1KiqCffx6EO4PfZLpopVzIOR16wEtCtKCkrf
9KeicgO05Lk/KoVy+GVtHjyKNnH6ROQ0NNenc2ifA5cklhLzvRPCW65Tu0h2NMFugkdQFLz4gD7W
2lIHzClKW59RxSVQ6MWSMA2tGRpp2/HzDEXTiv3GPxG1LvuI4IncclKd6zuBKJgCY+isp6ChlpCY
JX7r4dhRpL6AqO9qtY1bU+6FCM3GglU6EnTwXkGbLsf/vIOL5sAyZ9G67MrO/SgDNfXuUu4DUeYV
c9JMhGK8WIG4xWjyRkisMgbol9t0JRjpLls6FLvVKIId0+44No5hJk5O2lydBxttQYUYHvNTNDIi
osTCFToCfKmSYF0d6zhxgmzBNqbHx1xq8BLwUKT+vNRfPkr5rYxCYBPqz4HRBRx/FE98IrkiKV2m
1HDSjK/EGRKFARf4VUTrUQQZlMPFknizvKZOhQuMltraHw6Vj/C/WjTjPw0IJ9Lgw3GwFBcdxbPu
40uCw9ugIN/LTBONrC9cTA4f8IjLLWBRg3W3GOIoGB7mVLooyhKc9BetPJteiTlLV9C61xAOycu2
evuzT3G0Dd49W2TiujlX1659UHGTd02yGYsF7YIMt8I7Xp3KcmsAdUqxx9Dl/Cp0Ot1Ptl4UWjmS
xJpJtr7Ua+I3jiAtnr9+dnbL7m/K6uQ0bic99oasrr2tKOeMXCwjxUkZ7Jqo4EpOkN1cKU85BDl4
UJGZsUCuE1vQ03AMnDRA8wiZxjfk9286l4qOFKNNUu97RNgbw9/Rm4ZP7IeqMDlxf1q0dcBtQMv/
2Op0SkoH3DtWRLKQ/15MqxzsjKuuzSdi13WGj0C6m3DpiRu6kjWK6ScHiJy3SYTwTGXovLUpqUsT
7uYFV4S9JSjoI8ubXNUTDU14CJFB4oFsb/S+nPcywoMTpdADySQqU4bT1/aeW2bO13rNeEDW4AdJ
13syXLIfxHb4g4/iKScnOOWvtlABM2qAlU4cXS+YCXlnNY2maxgh6iAwftBB3dnCO1Pqxddtb/hf
32ZfZHm3u67DBb136XCLcg2HmWzixt9O+ItnWrHxV4KASxY/8xpeGQceb9mRkXvDJWdygyVgSJr1
nEHr/yk446dKSY2cGYbK1llgOlQM40L8SmVF/Q06aBOTJmMdcXYPhslGdKnJe/pZpnZwhr8kM6QA
yJru+KKHJQTZyha+SHJxRDHRYKP0SEvPyXNTQ3FUalJ2Jn7KF1aWi2sDXP5+JZKEd2Z5FS6mDtlo
/yzmo7cBgXn9/VD+zTGzDq1Dnyjj9da1Q8m+suYQKqHyQm1cIWuY/R7cfnh9jXXOi0ifMjJ7oBG+
0lpPDQCFFwqfspIJZnMy2BzQqdhc7c837KD/DaZ3Win12y8lw6Y3rOcrCAMOUwRHbciRzA89czZd
zkiWcnzVgkkdWJ+asaseuZ6+TfKIFoZ5QCge6RMD1RPTzzhvuh87ZLKWPDVOGTlLQqryZzUy5bfn
RzLSS1XrKp1Oau/E/u1QhPNGj95bHaQQlOjrfURSLu/zrvilFW30coxe5U3d1R6SnWqkFIKuGTmP
533j+TXE5UxNffnWqe7A7u7KD/8AAktqAV7JMn7a+VDH5aeXkPn1ZODE/Q53qD5w6IJFMjipbLp2
R3D26Hm+3ENNkN8GlhYBZRM61w671uO6KtUe9gb1/RnWB/aj5E4KnwW3Bf89bBi9EKpJiSx0NLeu
i7t105aGd17j5//V7Pj+hfYcHQKIilRi0o4GcsJir4qN6ufCFVEpkDlALVSIzpz2gLtrk0CZ/o+J
S4NHug9LQkpJPGwp4bVuZXG/cJTkz0a5ImlgRwch6ISdipamVJk3oFwJYBZ677jvQ7cW6p5n2Oci
7bNrD24sqzWKeIXTok2rd0TdV4XiYeoxHlssybDcjAxCXicpaFz1uCCkKyEBtQBp8etO1HewVWWr
vk6BuZKm3xwuEfpbQOvRqTiULt7prkXIw+LXTi9UsEIoPn1sxe5zQcYjeYnyFxFsS2XiK+pVK87Y
N8axhSnGpd671n+0h15GKxZM0rMlNRrypYTOoBRtw6v6uM1lobVE0+ybC/LrhohryPVy48Y2b23I
/ISbW91QskVH20rGCqjN2ABVNl2s9TxbnnU4znRmRnByNZA3s7gHDEBxLngBJaOwgg8yI4dqvAMF
2sP0bgJQZNBtN6cH6L5Koy9U5OjPpu7Ov1M7aZjpQxpQrmMuGNbI3kx8eEyIjkdg9qrMghaK9vzW
Gtw/+cJVmRsQ7evSBJtydgNu02ZUfqULIzw6SG9YyCBWfBgP41U9lUpX4BQGRM89P6BcdCCSL2Wz
rTY8FD6i4Gc5whJrhyW2owe/qgA5C/xj69AhWRbJVaLquuEDVJf0O6+IA32l5o7F9oCMbIDsMOR2
dNtJ1icx3RyAOZAtmrK3T+A18ThEuJ/pSs0LB0v7cUot6pCdLMijDZWEmgHIHH00kMirB53nFUmA
uY1ro1UYC3jnfaQvxKWEY8KGZiOoG6GomK13aPHBg0eIWvHc/wfm9R0oOGtmPRD1cjduUzTuvp+M
uGG1jDp+8WBva6QJBzro45LI4hB+35+fcpI7jV76Bzy702Ozm4lROKoR0RS+QVUPVN6WVWoBowyD
Omll9GoWfnLOYO5067MGkDG1AuNQoZSO+UbaI3/nzbJz3b3vPAVZN1er6jBHVpvIUvLBU2PFtQ+T
TNSllZkD81Igy9QHBc+vXvIj7wjIeJNKhXjQMCRXeVvawvVVLPN845JL4+TD7Wi+aV6ZKth1XzD9
98wmLl6xtMOmFKaNy6G20BEDQGaUfuxnDhW3jwIHgsTuU/Jz3wTsvIcB5UC1/qOMViTkCI14+0EV
0LhaTkDsDbmKSSnmc7pa5wCCLyidtiohLZqhf+KfeiRzMIzOH6ZJZ8LzxiKnWFt+Ka/5Ndw/7SLd
uqGzvEJMRr+vkCvlRr7yxwT2rwHriczKqQOrSfaX/kjxpAJLOd+Mz0GYe/57xczUjC3+ey6dtinr
Bta7zcG7ILT98hKWX3vYRwzmZ8RZN8uKF1ZK/ML64FZFDv+L7bsxcvobPg3dFFjh6OAheuNlsXJF
Tzm+j4XAXWVdP7rzXS3QLCZmI7P6u728aNiNp/xKdmBkIFsA3ANk4NR0H4kqBJmVWOjiVOTjvNR4
YasSgLHH3TErtisPZgDikDn+05iCLOzv4QR2AFJrZIcrttS/Da+tNLehVn6nKT4TQ9aGQq9U3z+9
/RvFCp1v7yDXSuZ05GOP0i1oBGJum+fRbZQmV5FQjM7f+anRaNkaaJ8WeHIEyfHsYR5ZQABMBiY5
ZaaNRNzCYoFOeAUEbkfelaD8fXk8J4J5yee/gqn9l26RXY0G6vLQ/s1i1QBN/O9/4K+P1a8ryYXh
vrpvsjcz6udW50udcTbZX6LlUvJFs5JRhCAVOWt4EMi0XTog0aUe5f4+4qATj5uyS5ZlhL4TOhNJ
KAC45NL3zpiZ4g0cVXVQkJUcfGgaXUqh912w6KKy4xRLbOWsGAOdRuGFB0YFX3h9af6U/U7KeJh7
o6MRKHML5jrfJBtEa+cd2bIe/km+tcE0XizkuX0nlni7L3FF/vX4wSU0bDr3zNnLXUrCL/KrVJ67
vlVLwEZpgz6hd8jnEw8eoioE2lDIgh8vJPhxcP1QFIgDyj4ZsEyDFTdt9QGZ7RxvIGgNooHUcuRl
z23H2Pu15RE/bGvIuj+K9NHvyhJfjhVXHHtLOmOuaUMySCRiprmOmhWDa+1clhrraWh6GOVxfRmg
WmVX0WFDNo3Gned6QbgDDZ0G3OLUZjXq/qzfvKs+YyrKM6mEEuxP5Ry1H01J8SkFOcXAn96FkQzA
fe5liBTK+z8tCsJ3ZhqTAGJz1uxc1tq+KrLuTKjj0OaVf2ziOiX1ibMjqUrWfwa+1bJP0k10gKgu
zkhyfBeWNGsSAWBSVrV0iWcMh19DWca012bQQetE3kifPkktAlyRJuUQPu9v2B7v+X0bozWjSYdm
5g+LE0mk2rOWjl2UKtcW9MeqKXgZSxuI8E5qqj5jmigDkORkpuDRSwIESeXOeuh+CnGHU0LvxYj3
zTk+9zmQynx5HT7FJd+mkdA2zaeDbkRx7du3MviLy3XjUHdAzC33wFfBkKXYL7rEOzB/hTyT/+Fl
tiEGd/zSfKW+HtHmSDWtfHqp/UoCZcvhWGQ703f7C9jT3kEUalVQ9FZhSgv7XFTHlhSKDHS33YGg
rXgWu37Yh6TcQsEM5DM+S4+GPT4ByGIFPI58TSYQhXlNh6GUrCzS1v+eRNiVytd7gTWFYAdmx12z
fAPVB+Lti4Mazr4IKzFlihkJvs1D/140vEmHwjLPzv44SgTXyeY9MUbIZx1UFe+cEzvwpHIKMy+p
Ld1ZRx9OnzqochbK2JY2ildaqa/Rk06aM/4lGCPTHQhF7RCOWY/iRo8cq8QiuO4pZGCCl1rhkMvm
+938fLNzcz8L2nFD8Q0+domD+l5ERDoteKidTJx5czdPdwsJiJpRVy9yfvjyiKiPPCZa/ihQ1Fnw
wTguIOkByxGHEPyUOna1HQNdF5CJiy0JozCpaOQ+dUnUHCkujKu302ctGKsOL9HMB3vQQX32crS4
V/OWy9oS8BCRg86uBtOTNIM6aKMJRNlmhUhvSBu4ze6+OFn0EZcs0Oi155scNgcpONS6bDHW12SL
yDVxnxKQabpHbKLRNg2SfrIwMuQseiIls4aHsVceBxPPCq54kUygXY9cXCVL3f9LGwMJwE55Rrpw
SCmXxWqdyUdJOjQMYvPUylxErCzmf5hyl04UX2bvmjT3326pYIQ93kSfQxgQG5LCYOyx810xMxfH
FcXvdmfu9clby5uTPlzNX8ny7jt+ByOX7M/W0yO/LoDjxL18fP2++ToUANArhwPXILQkmPvFSlDX
tlpbxKtJWbrA+ERUugvw7HTygW8Ezl1O2Us+8AYgmV/q7reZfAyJW4GSXxs5cSHe2oIDzjhY0fES
vGObdhbBoG7qVnTbtE8aE3SSGFGDkr/cGHK+micCcUy3l8w119J4sV4DXS4WhYV3besHIngGHqe+
gtQ6V5y800theG3HbKFxs3UFblvn8MH4eAOCapIbF7LybOJU8I8g1hjiniYOYpKIL8/N89ouUQVT
XI1wL45sZuZ3VASc5CXALcTXMCtSYzVsz1CNpeEpqF7Z8SYgw5VZWMHVo+G6stxtYe2tP4Dq9nPs
xOrVo+EXUHfFWXDKwKPXpU58GBrfWPQnOjRHpEZes+zEcUrloE+juTje9Oz+BPWLm3pIMz5gth8u
xhLE0p3tHmMjtdaXti5tmuxG9rN0+s41PoY7FGaSSVbg3y/hFQwerk5mIJEuy8JVVTKVPSP+JVMS
fVlGqvbP5DuBAFH4qZ6Jf8KMM2XguzocYK+ITXsIBDQvZvDFNSew+qoh4N8RRY67gFcRaBcvOAaZ
rKL5lN+mDiCQZ74RTZaI8RLyyifoEtjabkNLGa+MxF0lLHW7ilV/pBycsX+EDQ8i590D9eN+gXsd
ig8lI44I+TuBliFtW9Stxc42n6k4R9Mb/2aLloFywIRKjI2/vHsp8u//GafIYMmhv0cMOMztNjAJ
vFxmQxgMSynceX9+stF2VVTfjTBhcl9Bfa2i9mwMocSSwkrvv5aWFMlldlh0lciEm/UnU4iUy9sO
VzM/XSdGAkUQ3vZPbYWPhNcNL0cg+HssUmmEW7ileZmPUZCZwgrqUkW7ZLmxPD5WVohLvQ6KjsOw
FHpkcjAcdcORB95jR31gCHsdfm6Lumo7fGEUb2YNWbM3dSZ/syrwwXsp6Q+sDUb3wqv6Jrv4SObJ
n+i+lpzEc4EPrdnewzOYxZdr6J6FiOgYfP071K5vnSSliP4aJoNInOMqWU5A0bxrfMNZdveuQ+9J
QlXmt+OMysOpUpse7i2+hH7sLvHBS42awNvZDgT2WUaTU2e8ZfET/+XeRMNHfZWGEHQNBtI4ydEI
diCcsVnyAGbED030vHHc+gDZQMBYJKCAB9ucsaUyPsIlg21JVLbOBpnTSUHBFW9LppWglHwr/k2v
PA12EHXzODIau4PErxnNcIoRc3NVyGTVPRoWmsv+qWcgqpu8oQMlBtZBqCk5qpAR7QsmygI84xyO
3rB7uXFqIPRvdWfbWf+kQx1ZzxwTi2vOv2QlaTQp8BZyTdqBBLvcbVUecKjJdr302Rd/pl0bOYiU
DKcyIZueqXisRycwcl6ITEFhOBG20ja+PRrNqLlD8vsWtmsap5ID28Yhq8e1Jo8FrSRZCJOV664H
bp42UXTb9OUczvndVZBHgKiJuiylgTmZyPk8aJMzvubMXBHo9v1l7SIp4yDMtvryx9+EI7rTzYow
zii+xX8iFXsQnJ0znfD71orRaREE8+TceaAUEF/u5XxFzUgWWlk8NAhXa63VINTAr7Xr89tMD3tE
LyyPdfdN04eBRSOk02EK5BaLupmZIeWk24WvCcboWEmTA16NAh3jAjnvpFYoEbS340KgpzYyPnpr
jdW7C/5W0x2N1pBKObhhw82fBONcaqn9vIlsI+jg2RZKwQSH3MSzibPyuZug+a9+SYHngUIQNcsX
McNYRC0k+yXhwc1sO7/gEyy2gJU52hpis/89Lc3pqQhK+jAfKiuBQ8Mifk/NUbfTdTkBd5rcNrI8
5WHhQcnele4SMYfftbqaJa+Tq+OxutB8r/Ru3THvn7UKLiynt667HZt9N1Ur3ZCunsm1MNXVuzLT
5qiPKgeOkJBNNrBtP/ttu4a2Xa3ySUq9hZ/IYQx0Uy2xEhs7ZsKWfZAKF2F4eGELb4EfGUkRS3FM
+eWgufIaj4yaLMnKf84wOhhMfPTZZ92MFmVvlH8h3H0+DEIlwNpV4jPlRXKegpt5+i9W+E6qLc0V
ziBds5VPhB/W2k9Tl3STAL+KBK4KJKI1YPx/THl/xA+3jHvxe5RipGAJli4CveeHh3pzhJIsbwgi
MCnn4nqZP/G/V4UYFoqai/hnKIaq+YmPSAyoKDp75aiFX0jukQVaY2B6BYqsM4hyKKxW4S8Qhe7M
THGJ2dsYLlHH2mQYZhDh/NpA+WGn9uKwureGEh7HffSop35aL3TXQqXdM3OFid9isJY+p54LWKwj
eNOGw8L4DtQzaNHqMuXgDqCcHf1X6uMkMZLDtMNyTQxURx9LB2Xa5ww9FC6kNZxlr6YY83B59iAJ
+DNsUYFF0Tbq6DOdl8QxWy8lEhfD3u9zgNm6zu7Ip/TLjufvIxMSG0/nQQZ7ZsueVS0Da1f6r7B8
1qEA+8DXg59Zt5HYF/NXKUmMMB3Iicgm29twT5FHHknTlMgGD6YyGfcjPx5OLHHleUiVc38Omeuo
buIyW5oOuGmuksBUIyatlFXD91LlPeCyxqfLu0LnUjn7mwLo4yJX/Q+rMEb6E8ZxgtSL5O4yDur4
dBOmhJUqSsUT3q44Urzp+PCoIpKhwB0HCEPnwCN73HwpCtFvg2fMz8CpA9rgle+tNLzOMghSG8q8
bzE/dlpfqDZkNdLY9iymrrCFQeWze0TYthO+esRqBXUXeLEkoDr3cEON+IVjp+RcJDn3nwtpS0NQ
cCQWHGu+JBkCasG3P7G6Mu4ich/nouJm6xNRSF9NhNiRyGGnD5EzqzwNWSaPPdn3gvmmh4nbd27p
LmLdoiZfVw4o2sQC/zwpNiR3bdv/Oy3IazIBGaN0MFMZLfPm1cYnqJbMhhP3NcvsttF33qa5HBtV
Fd4tAczI3yhGFKL9YalWOhjnTkPQO2cr0iXRHnQbSv/TrivgpRZcjiXuGHcnhh+BVOtx8oz1mNXh
+qr9Z5GwaMbKloG02ywKfQwuUUJpBX4q9wISw1EoyU9ceIPUQ8DobDUoTve1JodDeQ/Cev629ija
ZW61GFN1KGO1/NyCHKe1MiuROEaqBKPEaabhj5HLWm/Ne5W3PFq9/dBUklykbtIO2ghxSuIGuXF/
VgXFzt15sbCDE29bxq/ORmBk3coc3YWr0wadt7GF7sv2WnagjoqmX1n3NRcU1sYG2ylMrg4+xIr1
j4iMGefwt8A8m8xL5amLJId5RUj/FFtndf/Mq+aWQQm41fJYJiHBuPFzDuc9MkmzwxbqnBeS7BHB
tJOAiwkYAWkbw6qJH4wED/TqOX30hJmBC3R9VFIEJ7iSg/Qo2VWGObCZCKlkOxp7APhqJed2afQH
ybBNTpqX8cMgQe2osT8ydpFu3RkCrtSXnjmu4Is+NKXvA8VTjGhP+9cs2k3UsuY40v1bxmuckePT
hWOJ/R1B74jmi0n8yAq0fC8qRrk5JZSx3RvN2wgz3UXaIMTa72tI0OrIPfcRJO/4UxFSCNKqaT0t
bX3QWveTgKt9ZDmEX7CJmdAYnzuL2169iaQrQXjjkcYDIBcIWjDNlJG7fDD35anWalcFpsVYi/jP
sqanEsG01H5lMeXdXIRkjvKnhAEGKa1ATNqshc4NDYEhZM18pQagvPpEq7Lk01x6CzhFK+byZ3ua
rvcFixfTeaQPUO/ikt8p1lWc6U/+TAX9ckuAo9g7z/YAv9Ya7NBKhKzHcBbElE+Vt9zuwxSMhYoG
CDbU9klcKeIZxxNvE4CEVqHE8XSPAwy2tHkV39q8sG4aPE9GsgEo8Tof8RGia8R2ivbudQdWhXPU
8ezQj0sdqg5dmZYWHWQe6p+Mi8K/kTFpW3M5BE09OtAY5y0vOfe6v0OKLA5LTEl1CV+ls/OTGEea
3npjJ2iSpSqHt+01ls9/yRebx2DFDmbLDFZLCjf6s6yqr/0Qo9a4Bl23XVh981uVNs0l4HknQjqA
XAfonizEyHCXf7ujNtis9R9AGwcEmaiGLoqUUoBaHfqyepTmRM0xd2N2sbXy8a1C6mv6escKDbbv
+5Hp5vm1lVsGkpV1nPnBx3DT2r47SOcbu3Jflb2u2wD9SEj1kmVLY29OFAlPuxSr7h6wKkBke7sX
FD3K4YxjepjwUVfzcVSZsRWZBwd+O2aPQkXZSuzIdsG1lrl4xUy4QQRFRF6Mi5cvxl/JCTmP8vw/
0w606KPk84TBiEDA9GQ8cdeN05swW0QSZ7eZNrXEFdUDIQO50Q0pnmR9yaZPGySVs2G+DrgLb+Ai
Rqfv7YOFtvZYUip0E6Dwmj13/IjOepCst9OSxUcyr7e6BwbM27z3IIh7a7JMw2Kh82NJaM7mwC9O
HVujg2nqCE2V237zYKNEyFrXqkc8+EWiFXq6AjjuToF2vM6YGvfbyV9UATAYoLI1SHga/uL6bog+
bxml9uVX7kWerJGZgln/Bkrcf+ioeaO6ZZnw9vvOe61KGSlK3/UYCV1/XpG0UwX6OlMLEFCC9Clc
OcdNBRAQY0S0+R8toHp+tRiKKKUHElSSvv0fVCVQBv8l6ZaSzPUOh2mZFkDYE94XNchI6mCwYMkK
+osZIy74s3Me4t97d6YxKnh8sz1NInnw4KkEyDFX3U+iH2CI+Ej/d4LIYfLpsQudzvZtdQoS1Cvk
Mftnq0b0D1JEP6uBW1gXcCODMIgxHp/njNA46uLoGVCWNG/Oiqp/mi6fctUzfzhhbSTmrF+j2beD
gWS76sgRmi+ZgjLd0jIKM5PV017ZqJ3k4PwwdOJdFDI2CfpQ6lQd5gmJasXYM4W/HecoGwi0Ux+2
KJj3jaX+JgpcxGQW84hDrYWcP5PeL2n+i8I+8b/Ha6wrhEZeoUIEB4a7njuiq0sE8+zvoGFqOJSz
81iKY23L6lP8nKyLH5oYUTXGkY6XMRwbzpOPIlkr9b58J3HoQdfxA69e75g5NnW1SKg4v8aGjPkF
4KQ/APYqu2xl3CDWw0xTxSFL+dbN3FzC8HZUTy/OE0jPn9QdilmSxGctadm8nxAuwygSikB4M+J3
dybC8QfHll7xFsagzoTpRvOyolbMOYvvHmP87W2DddnisKlWMI+oA2ZAi95SmgrukcFOwFGjfOxx
/nD6XF/QYYBF6Qp2PhsuIsys3TWqMcB1LRfx+1F9fN31XvicOeThryMuGSgSEYrvThe+ywhv82Wy
qDu7APq1ETBq8d/7+4BauI+bQQCNdMmUZtMhw5xDKxVvJoW95jTw7JHKRCR1ji21ecJGjp2dy84Y
Dge2/c4I9lLTWkB9dUqeswcQEkLm6KkC6JdiwtvN26+7Ri+5urhs3queQ+U8uBa8BddvlfBO8w12
YRUclM+nNA6mpRU4uoatwW0HYLf8i6WVY5rMQZpVEl7UIsErYc1NEBMiBor1rGUOVTwmTmJJEz0k
iF1lSFaySrWO4V0YNdwk5U8skPc7wB12HP3YrJvUk89sy6TA8hF3FKRHT/n2LknCv/OnFrOR1Foj
ZdtMiJT24FoKglLNeISxMUdUQQ7wTkz8qokCgWmsWGmRo5bCzu7H1YifxIRRphXl7JCi6AivpLie
Y7Zyh86oGb8/LVOHK5uLZ5pAwEV+i4b0v7Zif+KWuR/gfTRhubjrch8zmN+iKHe6D6j8xoGlhNCM
L3HMnFOZ2/87Tc2UZNVcbY4EUoQdIV0TxdnzYGpV4JVBxyCLeQMGzczRvB3jI5Ndt2DDcZfrcKgM
M3uoatlF5nvcN1xZOxttXh4t7kVegCm/Y+z+mJ1OKq0aLKb/A+qExX9TvxancmRCda+CzYTvdAhS
Nz2DXWjFG3MZOBZtJT/GaruKQl2fePFkmPbDHbrmf2qtixaCvTP7IFc4FqPaff7z189sYubJtwnS
Iznkp+E3GbDLekqjKTSVDlvj9O48pi3iBumfzflp8Ex0Yx/+ryJNj7IWSBh2SaxcPEw1TQE3cSr5
hKO4SCneeXJk4mmxCYQk6A0OXLwpdUqiyii9Z4lvBjCiK0HPsOzbtahGo9MrJ/ZAwG7r0c1oHqfC
ZEpp7xhZHMrfHLGxjDfDlbvpQD2Xv9Aavlv21ty8kI2Q4kfmI32cGpcu4f8bZxPTtKwY+YjYMGC4
UB6FJWBui0nQbRjt11PUgmu1uqcnp1D8PO5dVeVRxIapNHJscT86omlNnYiabulTI9WKEiDIqX50
OewXGRk2dL5+aFQEjIicY4FoJ6RWzAHOo2DvYSr5f7TY76N7zvtssXhZkJWrFXThs4xMfMFIZPES
M6s5SK2ZMwnKKDY+jg77yOTyulBGrWNQ47GI3x1TwZf76PgmybgFizmizC002J0Hv5dcRfOVtYQ/
wE2k4kNWJGKp1mS0obrTjTFocxPVj55IFwkpjJ5k99BijzxG3GLSe9RE84dNse9NQDc/8gDx1/7b
DWxLyZ5jGO93l63PeIVfipVNMuBOWipCnsy9UFPGL35ICgVQd+3nzF1nwIuLcLAqa357njRMgB4f
B8pCJmz+dqMzyC2vcW5YDL70TXxGuo1gII7nAOCuzKEH9HH2ktSDWXTACcUyMAXnjWIxr8tajf1A
B/RvbkaYs0MLJgXkFms0/Ea6j5xSD8qj7HoIYXQ2ADZrEuofBb/CF7Sq5230u6gA2oYIZgyv9YHa
FJ819oQLypc2lot8LULaQNS3inxm6zvEH06EktP4wj6ahEpaE9879INHD1+CI9QKsz7FyWvIrPF2
mNgawTG47q7GamrhBtz+Aw+0Ze+1iT2aEJubL1ILWKbuJqX5Xn/Z+89JMDiuBvsVg7RJxXN7t7Dz
DE6VAiNILiOk7t6VmW82jrYz/i978sZBhr0YxTU4Dkz99ylcwFNpgv4Ij8VBXJi7dCSSNnr8m2Vi
Kdvdxxmu1+Ujvs46rUCwdX3TRutiq5BYvcVlEr9j12VDSgWiaMdqmYAZDhSMZAgfHku7nfH5s14W
wC0yCBWmymGhJaZulsCUD5bcP+7nR+vkxDEmN4X3PMjpG9sW02b9LJcy7NL47Zqs+xzVwNdLH5Do
ByIkI4bfBmuC0n7NnPVRHI4caTHjtKMq9Pz6GOJjBjIQCo4qEPztAvKdvfiu8GOd/qwHmMSZyAQe
Pg1KprUzlTIvZhvv9kGOACubNL80E2XTuD9LlvoRa9kpRl3uMwqh464TKwozj7lzFyoqoW0ZDURx
5jSkD23ytKgOWdVLE89O8D9JynFhoDPv2Ake5qWwUX2FqNYNY0w/T1C99YSeSwszsz3XK583G4Ed
irqHzq98eCs87a6eKXa57C2GIzGZjfhDwTmCpwuSSTCPddkWTWwNDX7U05UEIxmM5MnE7mYPRyRX
RvXBe64XX8MtfFnrdoj3tCs1roE9pEiMW7/NwWcpC3BReo9g7Dl4pjgfNsG9vgwu/PoN9jXM80gp
Bdw1Vzf1aPXzucvhc2vLRKAVZ19MCHoWARwn4fJJ1AldUbuDZus7jqYd5zXH0QJ4Oa2PEFCQ0X8i
PBfGlEDZjHPhHA+QUiEEGKQRiD30jgkCeSmlT8Lf94w7xSEs6i76Bu99JCnbIf3d+E7Pjigwf67R
CKneB//Me+mORVhNN45oyywaK0HppDII18XezSX5R5ro0KLJpMCzCkcqSz1HIR6TGQhRPWl0Axt/
FXySiy0QNUYw+SnKksRJ3yJrd8sirNYMPDSYwBmU/33/u8xAsGavF2gbQKgFjvGe21bD4JL52EKA
vrkD+PUrJC8BvyyH0+/ZLU2/slq8CNrwc1T0WTM8/4TNzFumIhBwxG/GM25vAwImCF1cuEx9g8yN
udDucmwyq7lFns1R4oxo7pDrdIviMeMTU7e/SMwagvyWD1O+sxgFrIcLGEMRJDzxEqPBu5iNZSEp
5iFftuEl532C2CNEtD2qSgZc+uZO0HPEMqK8WzafK64YKBmVAOx/HK8ajoS/uMA4PgHnm0k0FjVL
GZiAmwtF33d4EnWFvaTLBuoaPCrxgOKwR11I3tFHiybndpbOjeRi3J7fvRZU/ciYCC090PTjPIqy
m70HzTL9xGcjWEpmhSY8+TOPEKTyva9TKEfKraUrCsbsG7e+TvnsNTBCaNexkba1aUoG+rSeHJmX
kPPGVNsv+aK4vNrZPAkA14c/FKKaFYGCOygC2r+oPzF+j+aqM7XFB5kh7MLHZzewPDKZnTz4yRCE
80iygG4GlhQEgehlVUO4Pagwn/9REhNE9e59gpdVjJOQHFwIKirvak6wp5zhNTxw1ia0ALThHlGA
fy+HEo2jASVvghmFjPr2ViNdaA4Es4g2lSZMauvAPCQee0ebGFvVpkxw8SO2KVBoPEpcX7P1nxmE
Ryr3teZu18dSVT69uglRHxOWqz/EJYBJiyasylALH1t7/IsdFF8YbmdrrTJUlZrJyDnraBVfYONb
6YU5V+2VWNmdKz+Ls5nhd02FU17XUzaqYLB/XO/GBKir+xmFRvu97JO8bRy4MJJ75P5Gszibz13I
Ex3V5dJqIv8I/pto+/xRa7s+v5OT9qz8ww5Y4Di+o+vQABzr0BNUbD3nWVruGjhlhOOwdw5GXZf4
6co3NUxrxYe7zDDm9XIaf6hAh+ZFe8gIQlcJClmTOKDa7XVV0fuP3AuhiegzMM4oy43Tb/K4sB5l
avGQ9mZaB9CF7gNqfdAlyL6jG1YVpKxxnIfR12szcMMFQ/Oiqm2m3j0I57ReMBHZOJmfKVKwDnJy
GLkeQBlztQgQk71L3VNrLhowSd5RBmvV5d4y5v3I5nsRr087OaxTCXbG7tl8aBvOVYYxafRq0fwj
i8+9pKiseh7gKYJulTmWDX7vKbiiM+PAfEZdsVT2O3nnTk9SqIniXeCDQEJuPp/cEdeh/Hk/wf29
ckg2LojrCG/gcU+I7C4ecPhLlf/KnTqb7IHIbjeNySFbFRsQAq9/Yf+otA1T7nvO04C/BCFZUlEE
rRoIwAgfVA8dXiH7pMcLvkVvz5IjDMfdaSlbGNCu0a9VPxH5ztjSLwPjB3l4ZGHcJ2aqQZalQyj3
wQC2cmVwlTrFJFqJG8dW9tUL1Kl4CAemfr9ZGZjdat/0DOWhuHoSZLcosJFVOL0jG+ToCxnagKMT
8B0UDiJQkCbuBR6pspS1Wm2pTdCR8Yyk7v59fWb+s+AiKM3Tk/8J/umgm2lXtrAd3x0mH5L2NrNu
gUa5sitRHZKGzGHP9KJ7R6/kuAnNYI3WXbaFc+zfDUGVyEtxzzFYSPdWF75Ykld9qFxvvfLE+gW1
lrxnJqF2gXeJkgAXSOH5bwsYx+Q6KBkzJtujxXu3P0g7O9m8vnnqoMoLyjgu5rxT3K6gD2SXb8nT
nDarpovO1UYKTaSEVaXHJWVgPEfPtTBbdkiQ9JUxTV5PgIqiOi8mh0SH5JM2uZQmovH1bz2d95Qx
O4WLZIsTzGEPFIUMjVO66+NBM+fIvnPcD86RA4MQ3p4o9AQnx554lrPdO+wDGlWtxv8Ix6+Bgn5d
gaMmVnGmjbgLU5kbXmUatoQpx3p2MjfyXK3BJe42w2KjUDRUiZuDz9sr+vWU6r044G2OGFB+yz0d
mctyx8tD9CxMgycJmQOgcjW/ER61zsC3ECdX+h8rl33wBWogFHx8w3V9FaDy5ss5hYjbgKfWkXsa
x4WO5TR42FXQprdg+MkVqEfaYiRKgmHHXfYTZFj85Gk3g4hl2PiJa9u5iDGtVTDBq0ndpiqdGW8u
H+c2TnABq5xElPQuFFzqd0/OBQtU1f2yuhMPi8dWKjPY6FHQs2dyOvhbjEwEBOO3iAPNkwk3JUzn
oYFiBFyUuLH7ZGxFDwpDYdrIYCBGyo9Ev+y5JYsVm6PF2TBJ8CRDjcIrlTYGFQuy8bFStE6fj0Ks
3jpw/9Wcqu8e7jdrQhi+MO3xPO3thMsY0Y8PKHGVDIDHZuQbv25bkM64+ok0NkoA7BHmJB7MkeXG
axAENW/kppGyRVpKTUpwOqcuNT4MnaCwA35S1cpX+McRLj3/iG0EvU7YEU1uzPhXqGEVk1PY9xZ3
IHkagRAaZ3/s7MtaUgDkR6SOr3/SySNXTAhqvIokV/3PdbXQnVKWdVvKthZ0uh838TC4hGfFUHGT
ypzq+OZRXuVDcKxZ69LpY45o0dbmARLglW3yUDeClyUUSASspDSnUCuG21e8FfBEUdL+Nu/bzebZ
FYpojakKdLdZ8dcToOdJ04v0DIBvzw6fD57t44A293JiPlUp2YjG+GtzOaqqsNwICUJSjKy4q/mx
xtwOGIZxy/bp1ClHuMZsxnQ2yjK4nuO8Nj1U6j3b4oafHCT2hEjwuK6OYmq1Sl94HZ0RGi9JiTKY
Mnz/k5mGe5xr1EtjmaVYgKgmZ/yVNyliT+TPcoUGyV13+VhEKr25p+UOLHB4WW5ilqThwFJGqPBk
OZUL8/jBoY3ryaed8kbIge4PnsJd9zDuBtqF1yUostxEovP/ufv8vnAjwadBSdCrtbJuIALEySDT
+S8No/caoptTuiYVEPnBQEt/8OsaOt/7LGPp7XTpnNJ8EAZ7wqBQEaFma60aBN9tkw8UomiXJPzT
rPVXYiLhcgw8LT+6cjfhZRaJm6tC3eRhwGgdthdADwys/YEnZoJonqSn8wi8kO/QhTmfqv7BmaXU
/VDfz6BXab/YyPQAvI2F/+szyvwhJRMPFNeOZdlDi72qnlKv044l2Xrx9/iq7Pg0PcnCugJCbM36
abzTo8tGstI1GkFKIioSJsezTr3NzooKYdlUxNrJZ4BogMJ1YXG7UlW7YHn0ktN3HLwT928kupps
fb4IdeQWNyMOGgkdVw6Ebn82uvAlJgncM+QvcUdaacHxdrup7zTwbKXx1yYNmFJ1Uyb5ukQt7Czl
RnAIEymsKNGls5kREzd7W2iz9lSIG0F4Rb3ZKtg5vwHXcDCuSpEerpoApkNpHyVAQBdr68TROdtX
sUivkW/su4pdJ6qPq/sYw2DQbQuPfn9MtM4+4Y68XYLeVo1IZSx2Vfxlx6THyPOx9B32sRUi+3/u
ymFBqNjZUrlSjrdNGKxK1dSzdqaWxshZW2WylooQHqT5/r1vupW1DuvDs9Z/PDNWj8MczkmffI8T
jQt2/WbeNMuCMSBDahTB83sF8TC7FudtBGOgC/DOn1TVWtZ8lhTkbH7Qgo8UZQDd/2wGxMlNF76s
2B/T1+61X5t6NNEpteX3bWPAQgx5kLVgPCx8SEWlQ4UdR+2VQQIWGrEioicq5P+A08U5fodkJVGS
u8p1Xcq2R1+bxWi5639qVbxV18Vyb0gqkvWu0BFteCNUgTPfTFwJeamDLR/PgKdCga9/PLBpBFk8
nsBxSuNoPXGH7FzIs0RIWzUGff+5FXfB0COlv3WWRVBD3dAN2zF2P5zdP9+3RhkelWRgyA5fQ5YP
vXAXIo867YBkaqXwTC0OkLruwjpoUF+iYqWt8qJRVj6yLy5MhujHZyQXG24Fc02ONtgmZB9iBEMA
2faLkhWOCbRz/33U6JmHCNs9acxjoGO9QVcsSaDnkInmZFJ32LYRDmxGYHH0qJqolYxQ4DMg6oFA
K3JcwgPTeClKq9sGWsZPGCS0hIiVFauu+gaJXaUNpKPr3IT5h7+f4MpxjUjFMoeqtAfjZSjDM3oX
I5zWRV9fjodrVHw1p45tSgYk58GopmFsFvk96nvWdU6VYreQwFhk5obte+UscFJ/JhE/oehLRLLg
BKIQYvbkJYPrn8aDiFeenrYzUmkEypLCU5Ybs7dJCWzLC2fAyv+MftzWEkQSuQqkWZ3kFmtra9JP
2zEwwJAB0EtZnjHxA4L4NuxLZa4I7xTL/gGtdm9JbOKoAVmMGhI3NipjC7fpPbCDIMUaSbaNsy7z
s8ixTftQhpwCdr0naxfU8zZ1+4KAoqN8Gt82YgXGcagBmMKcVBwFNq5Wy+7nm/GbKU0ESEu1a4u0
Ulv69PJY7T3i568AIWvj4+WU05NDLg48XtpubZIycs8sybBVj+w7ppCaFg8J/qecY/HjAffTPUgq
0EGM7OTEfaaZ2cILkHMiLs0jxtE219yXv0v+fCHfI3hy6V6fuR4R4ONUossjoY+6Aax9RcXiUQMM
6Ehc3aiY522K1tIBwek9lJMT9AjUKKafsW4cN+kgxN2yLS47vPpVtLYDmaAxS22g5KyJbRJ1evmO
V3igKW7vHenvZSUp8K3lc9XFJpSU08PhY8UXb52SFAplS39MP+kiprD2Sjdgt4LaChmZjZpyEZB9
mMaACyNtizvM5T9Dpm5ubXLG9cEAcoSr7LJw3I/kYibSnwQQz0sYSg9T63l8mN6CFE6jWHS00FBT
/PWF+EpZoqei62y/VB923Cf4io5CLEURyhBOixfEXjow0omoV4WJJcVqT60LhO4HuuKGxFmacfK5
n/Jc2ZUOgCQXB4SspA5mtMBDDomTPs4z35a5Y13DJazJgN3BOoVVcCJWRPi1jYfYFrHKBdSpNI/t
jc5i2iCzpscDW+bur11RcTJTxU0v/w06tA5em2rpLPeUQOdKIOxpldryJKUnhOkRsnVgKiIsgN2A
TbVAIXOj0PpbzXjsCDv8MAr3uq857QYvAiNICoh8fUsfL5YWnX4N+SCdnKOVbgOZz2oZaBzqfIQ6
1UMHDmZsQq5yO6juY7pfxg2SWaU03BkuL+zbpfieq80JK8rKs2RpYcPFVFI41P8mwydx8LZi/NFl
3oyjUz0z7nyNunjeV5PeNEdSK4PTpneY+56ZnEJCgCmCwfeiLI5Yl7/B435c2YHKKUo8YbzH0QAh
98rSZ9pHR+XTLp5t5aOaBBPtBSzNANwWd+Bczlj8wYd3CTZ9geUroyillHAGgU8G/A/IuiByV5Yu
Bd4WRwxF7c6G+DGeaTc1INwixBTvK47hJRzAoqzMVUCneT9xqub4IVJiXhjd2QHSdz4FkLhBh6WU
hIqWebhR2jc9JxrN022w6ZO+FnfIZwKCQrYO/XGnOnG19XlDEJEhsFa6gJno1W5gyQoWxaQTJ6yC
qO5kqU+fxR8SdmH936S6taT64GBs0IRkvM5JYKw3xPjkg5NZJxBO9zB5Qr2BGQaRRK2U8mzzR87l
vXavAoDDM/8lAbZ3BiGfTOv6bnLHtz0KF/sPlwpKlpws9CXH5igi6plJBUKcwziPTbI4Gvj9Ky3+
tEAeTkc3PsEmWB9en8eibqJkg4wl2BNzStDLIMQo8WRJGlk4eChuqngeMQnknrT+2vz24TtZQ86q
dsSpZl6StrvA72R8TWR3rPlJsPo1SZoVoc6BDxDt5ae1qERJV2UIqKe+iGNIVbHUbLrh/wQBAZYn
ecHpJkQx5F3oYFVSJLRVog8xJgDuAM4GeXQgwWlUuCu1xmMGVGmcIjBcrQeNKtehdCa8xgReKNdQ
+yjqYkMe3dA9xcSx1UPNnX+GVTVEIekxo2jwPxQq1yIqXAIJT2s7gYtw4cSk0WlHpIvaR7HTodCk
aPtUnV6K/xMaQxcFz62+0BTixS5xAUlVMGAOS3pvgjz13aTLPKBrdHEfr5Nbg/w/07+Q5Ds5eChd
6BODsDmyBR3VAvxuCsEVdzmDbsvcEY0es92OxflHr5H7vPvYchxUgnescf/Jr7KhoZJKkmDd/5PY
gDIGxwtBBX9bq8ffmxkRJyIRyh2XJV5G9AbMR0ulzfd5JivSyZrCg25rlp2xy7w36Klic8xoGuBt
pSvd0IzzIJJbDo4WiXjd4Xg89ySChdReAgh2ikfQsElY99qKBNVrBP9KupwSPWO78HOg8HPjA4ql
y8RmTKRKdcOh+zw61N9vCpJL1KzjVOoOs410kt0ucy15xuH8ng+3182pvzbi0AlREcjqFK9fjNRU
rCba2nP8QWkGqMAUlNLY70d5QSlhCqs+T1cDc7GepNzXUIOnVqSlpbXWhSi2S0/GNSw4vzWbZG9N
Hqx6aPPY82mfL/u8X20NlvHDtqg8qY8ZhrViOvqzAiGHkbsIDAw8WjPvEIg34hEDA65DArNzVBNK
2CXrn650hsRir3k9YFv7BW4jXzXsMnWjBPNQL8GlH3F+fZ76f4KqYOaxB1zU7N4g8G4GI3dG0EfQ
+FdhYFFak+RsoHYQ8JXdZXjqeVRSIJ2ovUWikV7o67zXpXnJupPVYPnAGSx8ggCzoPb4R+UqrHUo
hrpW1b0k7uOIKr/s+mPFbfo5DiTIstQeiFS7Ra0K3+EnNlCuPNxU1C6QwatMEcxUgrdqhCt/H+2n
dDH7tTSSOh3jYn+l8YWsi2i05GNRMtlecgx0/jiRex9ZTyNO34UNsXrFWZQT/v50xElDcoEGK+fJ
o5Hyd+p7OWHzwZpkg8NkM5gl4+ci1jGFbSINR1WUI71ObvAHRBNfkgXwZIp9HIKUJ1EmLp5+DjkD
xm3ugXeA4jLldUEv4SyR64KIrEbdT6dujstGYIQ2fGReMs9Pih0o4eoPSKqaXtNCazAAoNCHYgKQ
POxDmtQW8deuKSRVL+R+m6KiolFNFUqz+ZXUHOMvyXpKFvQ5TFfqIpxGBlHZqiZ9VePqPVBGemU3
kehEus4EIfEsvDfSGak0398vx7BeDHYGAT0T2HuPnemgmA+OUYCvFDEX/KrhoLEsf3hmb4/oeVOe
xza47AuS+w17H5gf4ZxkPQ+uGgKXEqc3PfSStfwYtk5LzunxkUilsgCrBBXIgch1YFZ2moiXY8h/
26PsxM/W6n8zR8rNAs/WalIIeKBHqFuF8tKvJesbdGVchNy9OIMGv0BO6gYAuEHiFpWfodtRLN3R
Lj5kLGUPNtTuLiY0hj1/TsBzE6Kix8WtZmyd1+AimGJvofzlofAzAop9R37AXuqrFofT+hajqNXT
zskbNfZj6XSqLeInxnNMozXFV2vRHtqJNsE93wf++4+tOJPR3EPS6eMmkvpLKKHH59RcLsEqx2zS
UjgB/lFP5bs3Pn+kREHxckXOLDutSU4sHNAlgLE2eUyaNyt6gO5/+1txbAWOxTPt3+tdlf739yJ0
Dz4mXMiwT1l8lMV3TvTyh7Ppor4qXo32SLME+hSsxJTrNUVIHQJZhzYv6DQXe8dxEJ5J6tKQNhAw
xSkLRPhFjRSdB/miL9QnydWY3u1NEDJdD5I/ax9oegE1o8A2b7gCP2wqBlWmhfjAfXbBmQaiPTAb
RfI0ILJhXRvqYuwUxe/glT8+EyzvVnMBRLhDZLS2zbnoKzBa6CFfCfU81l5Afb21uTgvRO/4/MHa
nFugmmvih5oVOz8pXLK+EF5r6BN/qgIDDqOT2H7XKREwXbvGuTm+URDooOLVHKcYfNoJAAuKBHIb
S41CJVjl8o+FfYAfZOGZWlm4/EyFqP7jCQTR8lbDlKBQCfdp86MfLN6tXF2wCu3wo4sPHCqLRVva
j6loVuny+CtC9Llqqnr7buO5WmJdts2716Ddy9tGmMpm0d0VGbpm8VoDnM1RRXgqlbaN98Q+KW1R
rJM4LNrrHDGwNwbOthWaTQrhSbXNUfFD0+wLN9UexVdmQ2fE9CHdyuLA21I6h7llI1c72AweLYdy
PUmnktUjTEMzRXvTIoQYa16D0huxwgr7ifhgQ7a9scifOD343ZcnBTe3D+9ZWeqSWaHLVEztqreY
uifJDnXcMxBft6K5P6IGOIEbKE5ZQVXXUEv0SK63KmB1/H9hL9tQ/KhwMAvs7e+/nlbOm5477KFO
qNXU7E0GIFr1NtdB7xj2+BDpO+OCOpLTN1wr4oSowsMMEJsEAKl2oQG5A7nGfe4nnHsrJ1QHzdWb
dhAQk6dgKVXaXyp+7GiZqxbwOAhR9m+Ba4DmxIIVA76SevnHJdRqMY9HbZlQ4EN/R2GHW2bQZ/BF
WSedzrLMLfimxAn058tAz9ShoHBN1Mlo4X/kjwxdiUhM3Jz2ZFV7YC1ovax+dm52wmIos7IBIB7M
aj1fQbVIuOllHrWjkILOoS96WNm16U9Juz9OZlowrmZZfUeOq44mO1IyOMvMeyw0edgvysJiA9AE
EAtyihy8E++SrUriPZjd5+U79f8/v1sQAjnLts9sFkeSEQPITydc3RvXBbXmlwcSTpCvBCf+/ppT
Kqg8BL29s4VWOGtraqKfeNcYWv0Zr1ba70+OWW3iDMlfVlI7DqTbUy9vNWWJTt0TUXbzx8BTY2Qm
bocTf9/3uBss505uHd4YINCIv9KVOytCPlxJ8z4Z/krT0px9PwSuNw6iimegiJTwhRK6AOfyvg8F
uZgFDyDlbzaEIxsmZq79AHfWFNa4VHMalmKfRkEO2Sgk/c1oWFKmRpxpJHVK7mCzmmOBsvuZW3s8
9LKE2XpA7eZAV7kb2OvXfgdicGNzcVs+sfFAUZsYl6EcTr7SvLCyLVKd23jvdewymfM+mbHwuu/D
Q76fRHod5X0gtQGc27wM64KOFm1hhoBulXjtXarv/tRssOz6bFxFaai4JhPGCi5+DlIxOVbgd4Bd
JpekifPvxttm21Y7OxyxqgzVjVCrBSwTNviiw4bfxUSjjF+1VQXDnGIBHfXCVmb+J7q+wGi2w0YO
mJ+YvgqcIQ3LWahNVygIil6tZ8oN2meiV/e7Jgj7TVXEhNOA0ycVPXJ3ihx+wNMyLO8ssPt+8rUF
MnwuzWadKL57l0u9p8knYGZT5r85lkHog5A1/WOEaOhHkPC0uLw99vvRcYOQgpxsRJasyZs525ZT
LlkHQmzbqNOAueRWuM91mEhJoszq0bwO1uNTkzqCwOZQiMCZD3Yrd9owuR74iTJb0f+vsr0Dvnsq
xKrgCfWOeFj4GxayoabhfQMmVbwevVkPpDlfK3gQtiYg5ocnePBAtCNgqS8ivv3nebzjRGbl3Ipj
mTimvEpv9re6On8/1m5nwfJVY9yVCjjQCjubWOeVfMPBafxxExDerXSStnZvule5KVYxoGrthQM8
x11w2gI2Km0kAzfD5loeWALuFc3kLttBLLE3DnAzO4VD+d4LthGQvXBN7BeWPC8ekFGBb6/vywOt
8FUhu5NE0sOTTCUtxFMB8N6YmDn2lS+V2R77LVkkXXSZ6gal2vOiBbFKA8cx+MopLoh1p/JLle1e
MZewRfo4m8g6SnO3Iu4Tll2CXW7Emak2HESDYNNT2oo5YLe+zV9IjZCMJFvX9YDwjKS45ADG/tTo
yDW5powhUvP9GTWHU1YNhdtyIe2oZd1J1gb4LIB89+anXotrvJYU+ZMD2+cNeiZDPpBEYo/c6oio
w2bW7cY/vRo9XR3AwijWlQgLJP2o4rgtlygLrz8JtMv+vqJxhmq5U35NcOXpCPDvnnuDHujOTsyC
cWOQnykdEvC8UOG42schKqbSBD6Lk1eaFVdLgZzZquNpmsIHvdoUgiD88UUCPm5B/8IB903ASV3Q
BgaOIPHzJqBoFQ8MTGnNryaSJxfKlb+SHpzMBBhbMCQG8EsXCaF9GT80MkX86gTdLuPX96F2yo93
Vcx+Vz0Y6YHLmPzms+sSrpUjIMUQqwYrHBdLMY8G1qIywfJFDmIgPf/loFNC17OQpK1zrjYEchIi
LtD4+wSoJ4hlcgGoWkXoMWQ8NHdgTvyK9aIOiR6GA2twzMs87WW+Nj9O1hZDTIHUHq7OsjQhFxv0
xcOo8maHPW906IwZ2z4PpRMJ//dg7mjKw8jsBM2v6lN3RNvgv9DJyz2J1q29DP65Jr/jh1+cijGL
U0vTsDHHMC0OW7Au0KZOM/W2i34idU3Iwei/RYUIFz80rQuvfv/++ozvyvpR123WEmrB/jcKr9wh
xerA/oXvKI2bHCnAY8yWhye70rq0tyHiueTf3UgXviSK67BJRfn4j5iFHo0+SCpycHvr7e/hZk/F
4GgnO7JGO1ug6TSgArtDQAttMqNr12Puyk+sXInGsyQVyOOW5bNE17Nzl2bZ8yKuKv1/MF+gWsaR
l7KyU5K7IHiW/VO6CeBMI5CVKNRUNGpdSOddnyrtVc+txH0abbDeip71DzCWOohNWJgxT3iGENne
T+fcICxtFPJmREOmTWyA0E235/CBf2ATXpSvt4tpuXTwqwOxaga1fM//mPCfBc+CsP5QEAuhwXn6
WR/7PAJbrd857fOWbK6xLMLpnTrA2nP04YAVWLwmCrV4aWA64OgGIsbpIPo0hVDWcogozcYnDGL3
7Qz5epNqZb+pbtTyLtBbx7zcLZOwwhXX3TGL1P0a6NLv+R+gqpdoT+9tlgngcXr+HPWI5+2qAntR
oCtkp6Y6b4V0eiiXZ3egWyqL5LqiEOg9pejHZ49C3X1d7bqyQnrfSm1m+w9rudyIpghvr5YnKN9d
4I9TX0Cf85vOrRMIqN/DZ07zVEFwUAdgrFe0TIKintGWlGfTNdyQdyoje1BlWunHb8wCQvUwl1V3
9P/B3NlwWID23mQxfGej/nxUYRsuclQsFvjubrdmgdR7AgPhJdDrSDDVDPV1il2NI87zO0GAE2S6
oOKTBzeUQK3+I8r1wCZavW8vRPDnr1Tj3qvv+p2YOHgQV/2NLoGCAyxkyyIAwS7ba7OcsiiOJzGo
BMgyb8eK9TJtRc47g3NUwUKvpbwVvYfSAIl2uvzvW3fQ+HcI75rRejN18RchAe+YQggIFvKCdbKe
JXsK/KP18wmQ/imFqhkEsNLW2rEa5lOwKPjduzhgEOObqJ3JNwQp3B1b3DFVCZsWw0oq/9DH6tB2
+FiuhZlZPE+MKryI1wQY5W5AEkNoRve3zk9q9NJT6WSOlqCcpJuUuoM+IFIGRkyZd4QBTr8s9PJG
pEC7OxzuPTj0MAqMt/lBmV//tx98HP7Dda6wyRP2GIa2ZPE7ZKnNIzb2N3UGxYAds+sovSEU8b5Z
OOIMt1fjxiRFczff0zuatApfzcBTwqbjG8Pxxr9ipo0omqPx+ZqxhUpi7eeRH0o4xrIRInp5R/BN
VyB4LDDRkLK8fYj7nJMRnRHHp5vLFa2SxlBUSVbdNFMFLFqEIdQvq38+DHavOHz5XkrnntKS1m77
jJkoPrWg2YFSo5fpS1pJoM4vLWdYcnOMu0e1t8hxEabCNBHW9sNhqIPwfJcYBj6vuDC8Xeq1xcY9
saYG0N9guhFcV1G4PVhC9rTtY4a0PI+HdzRSgbZcL9XwJ3zqPN4NnHV6c1qa5yDzj9RQKbubcyXJ
qzfRZG+nW8kuqSg5b1CkwTe2irEMB+WdhFS/04fYRkh9s82nFZ1LqpFJlNs4rErhncCrmodJgMkf
iNhMyfEF38Uqyse2vBIMITHVDNCV2tZM5+ru1RU24SGztuXVl6ULRmqmGNIjLF1U56ImWTpNIoWo
/qSXpfX9SSdwq8HYUu+FX14O4LllpqdTuY0wztSI80ed1TcO5lvYcDxukFxBd5jjf4HR6iouyw2O
bwgTOaTX/0YucI9XKKYuwSn84DJ/cgN3kPY+by4PTs++suarKWah7JXDusCdAQLtPuD0ByfdXBx3
HWNwxu9uMvTc4NupqgoaNaaTx+H4gA/Dm3yzhGDCC0WaNFPNHkidf8D6XU4ZEuXaO4auI+7M8zo8
m3i4FEGEd7S4tiJkcorlZ37KYqDNDlWCmlKTshEol31SdjUewsZR/ugKrLaNKOF6c2g8x7FI9Psg
CsgxH/bHDEYPgotQj8QqhTH7slww2DajlEwFtPm515+019808LbKKS+zTFXG++7S54trzUspV5f9
h7t0kyeFzWFnxVQ9mhnSVu1dPNsq7KiQm9dYhX09Uj/dVhuVAvoioxvsMXl5ibNubiRbrrkLR2vH
8CCXsebLaRbsOv/lE4ZfiTUtKV+DZVZ8uHz+0SPg4kuKZjCc95sL0/o3uXNc5nikrJ74XZM8kpA8
tcbno46asKxFl120Xq38FAuDPT2e2cKpHk/ZEQ3j/C0D6/AVOgKvy/DjEaf/JA9pyUEL8MZkK8bZ
jjNvGWybQjw4LKJ6Sv6S1vadQkIS06MJPWAtQFDvOsD1i12UZcp8fyB3I8VQMO2xBNl3LsSx/20X
y17hnnFdVpWxm1hB/MYnFf1/FUCBICOs4nNnlBdovWViBzk0nuAcYCT7hXXeSgMvUQPRhjmjRSSS
Sv58yyH6W56JClZO6MyfO6H0ykjiT0TvE+m1W9oxOcUs9Mp3WLCnWk7o2hZiFt81qIniJdsjswCM
pcwcnT8p9d4RyZc/+MjZTv3JzaGmjIuZRmksaqgSbXvgLYRa26LUJnNxm40BH4WVl5xt/whdtXIM
rzOo87AYuMIEDu56m6dHj0E4nhUy8nqlGpotLwJ6OE8IDArM8dizlvtZB2Z9Qh3zq9o20QahiR1V
q0QfjzOphqwmMfrn03b4nomkBBtLgw1xHagz8/tyOVUjRTPztU1aJOaHWiS8u4Z2sO9tbkM92PUl
vyvJH74dXU7CxpDulddqgchibo68Pj5zA6JUAvlVceNLQuZuBdYm27MyU8/uIaEisyX69REPxq/S
wpLAFDl6+cMGdyoiTEkV+oUqp/ak2xiAvpbXsqfNTG5ReaztGxcg9eJdZBNmvZj16VooYZhEfEF9
If/EHAfo83cP6cGLdh1CvPGpJK0pZJsBZlRSMR5kzcv5qCCeB4+2iXqSfqFv5j+xMYFI5j/1IZVP
qe/ShcAyVH9yduttt9FUIIahyLfj50HiEDDScCChUMc4qQtTI/BMUISM6AwBDoMvqQXEEYzKvpZv
12zBVf05uHn3xlCY7pi+6pyFfa6+lXeXyvdNviCGRSin/YQxYixlUah4FkgdNL72AWsgJKFALZW5
Rdbkccui58z7layFUj9aw0zb9DiGXiNdVgGYk8gIQZSEyYNAcM1pPZDC59nccr90LNfIVGArwVHs
+18Bgfo9NmawMRk7KYF5glZjryCCa7Jg30LBVsMAJJzQm+i+1cKi4a55WRywhHYTcEr5DjhVwQu4
ZmerdL6Lk/LsBkZG1W1alhUO3KH9QqZvB0Fh4AADrHOP3UVnd/1sK7SpFu4YTR7tA6pfSaCjaWMR
Ynak7AP+h6k8oe+ctw/k39encT161XuWTm9Xg7dz6a5LwedOC7s7znG9L3r388pGCu468fm9S8jS
icJJjjQlaoKsHCQcpROnbFSuPCW9NnQXR/pLerq5LpHw9QBaZOhls9m16rUgFQW3D2sSCMWu5Xkg
zsiRQfgTi9R85yt2tJ0xQsAL3bEwe7OKytNCe5DuuILyLDhGKE1FK/vL2TboInLnSu6mdfzJj206
T5AogxPY3+drxF+LSK2BE7XDPIHqmwlCIGHIEgItFFVejuRY7cfDgDkJBckyokH04lbrsumeBfh6
3O5+8h3qNuWMCdTWtnMpF33dU38QDwj7bWM42n5jMSAhxz4ny/de0NCVVoPl/GDWe364g+fWoWiP
U3pTqoSDvllyUe9BsWd+25XFdSCvbNaU7+b2OHjvay3VA8+i083PjGv81vepGeUtIQ0+QS/gHKmQ
jO3iH5H8vWPYI/SE5Mwnc2UanOQJov528xkWnVqndjo/jctFP4xNLqOCl3Ul8fe8TVQ0Ad4vwr5B
L2S70PpiQKB25HKagSLHDweVSrgeN19531dcLVXb3RUywOlrqsf6rRrAfFdq9QBrFkgrSlKC9zDN
g/3fNBq9pNpv+moMwCPEtZlMidnVOrN3nUbbeEK52VcBYs5r/87Ue8kXSznsntt8140M4zgxoevj
uncot8N7DOq2ZhjKRbWf+9TvCNWSEvw3Tx7MHJr3PotYu+9m+01vcnsDKqgvDiACO9DEy2z79ZBM
bek9zCMoNMMf3Y6d71noRIloByNR2xtofmMPjZSMRP8qYwvWiKwoRTyaB+lurDctan/DD7LnSCTm
ul1IGDJIR4cEFa12PuQ8Wh4RmZtRhSd1hjOb+PTBL0CKnRv+XtvhkTv3pAPTU46UHP3ofTrmhUmr
ka0oPstN9Cq/1v0mVaVt2gS0rYiQVR0fxI6+ZOsPVzEbPCdGE2r+Kz5xiPxW6nhvi3AnAAfJb7sY
rigOwyGU0KMF0b6+910ZOxMs73OFtzYqh2LbXh4jKoeJb//jknvlGbMiblqeHcVkQHDQUkzI0HHQ
u7GbkTvmeT4JPEVGDQRrMpG3F4zLLm2bUr7a7UZL7ZWa7WDIH49m1rUR0Kc70A8D0xyOFJlZbuc4
N0irsgHlDT6wWvST5ZPQgt6QjigsWSc2GSaiX82UK0vZBAVlQDbj/lWw8zPR40tL3FjrVz09je2S
KlvXFkU2Kor4IchLKvEBPqjfNAg+8o7r1U4BFuhQArrF2YAJegySiAZJjJC8oU9jDSlW01aae+1O
ppl4+VAq9xarTKI1eCGZ163orED6ZzuKAW05gQiLdc7ixLjovQfXsTZuB4ezG0vRL0W4vhdm9Tmb
59vd54thWiERbLE17YtMIND2h44QlMyFx4L7vJAGXzrr7yQbSlFVrtv/rh8cpl2E0Z9zAt1VBU2r
PPXQc0+yb6gVWM4nbqgd1t2i1Ja3k+M/koJHGZg/Lv2+kim0nN6Ogjiy0CdEaOIyT/0x6HoKmLQl
acJ/obCIW4ZuxWddLzWj5LHkPDM3B3zfdgD8Fh/Xme5kpidGAYrAl9UTADjwz+0QvXugTZw89yoN
+Lw19z/QhT5ElqEMc866fdjVsXSic2br93tGvV7ChwSsfdoMLQRFpEN1z3khjOimZFlBL/59/yo9
6klF0ZBkmtNZWzN3V46xced+XlKoloUoqFkHMRe1HakAi3H1xYkhppdXQx9fObrrhAHCjbDXRy9W
u8N6VCDyhMUvqNRNqgUAsFZqaciIgqpAaymrc+icfWvDl+BGhts8F63H0Dmxhw+0BtNUvlmX/0aA
sSWjrTUJ7cafQTAk+YeXy++WqO7Hh/C8YOl5B+A4XKf4NsVUPsCmNASI/mQ16Dr2V9Zu4IewWc73
EpXn/BV2jwkKO6k8bFGEsMRDn7qc6a9tSmlvy1RB8/U4qEKSnPvHfzWQUSgBkC3hKIoyn20dWbGz
O+MFPtOLXJ0jPVUcq1EZBrrnlMipQydaExKfXn6h3nTv8cZA8NHR16bD9vUgVlxx84Rgg/Eg40I2
yoyz24Cr9oFxMeTY+OSQY6dNKMGoxBfI/xYI4hzm9i2ezI0+aDVhe9uFG5Sw1Tjh3RwrFzGsVuk/
S7Pqjt4T5VnhlRta9oSa/cxIZPTxF2QDgATu8m9Gznh7DDMHmYD1cWAXISsZaOgQBzpHw+/+xcQq
P7F5VinjQJnT5B6JOhrTN6skuKsb1rlJTI6ZPjUKfPZugu1F5foioyor8TJKeOKONUwpSqx/dswM
nP9htoIAehLa8PzUzD0ze6NTiCff9uLd1zn+dZGs+7LmL9PI5QMVkgcPgXAugQd/22pBsxtsxWv1
LwvKioV2P8lvjJra1IEC1sBmBq2NkLIQhQmFHf10BLsp/0GQzRscEydFO7qXvvl+TsIMN0rwyxLL
GrQ0bZJiOYtMrWYzK1G+p726XeDQxAJY/KGGE2tHknYbRByMbIEVI8Elb7au7Pv7FGb8mrQ1SC2t
0xikTFxF2pLrhG8h/3yQxH/5XGmCYUp+uSia98mC/tT80Mf/ndfSMfNgr6QWyuIhG2OuqfdkopBD
KMoaSYs2jbChCj0xvkGOYhHGoKeacTV/iTLrCcZuCaDYj43uKA73pjWlJHbM/8lW2627+lcGSyUW
uB8kFTLxI7whTtJssOr9ou4YSLOdARCe5MuxtjvDeztjZo2dSwZDf+EL6eIYu0N7Y6SzdCxetqAK
9VjgpwT+5cZ7V20M8En8WZFLqg/eWt+C0mtMaxDbc3pxuJBlB1JtLcFdnwBo3nEHJtDoM0DczSTb
W2mf4XQAoPyGTvtfK9W8hhOaA2pzVjwIcJqqzx+4WxB/Sepjg+O9xAOn0ZKUq1HoTxsYEJ4721vr
UWM6dN8QbkocZ3qIyFALc6wv5RoLF1JBJ9unpQDH06Cyf1mRK3O3hv1n5eK2U/7owoFBr+cVLXyZ
6unr/+DRjvoZ2tVr8Fw9btTWwh3qhkNqvddrtHBgGeCwNLQS5FkGfPfYz6JrpXw/9qN8f8xux9Gp
pV7KqifzV7l8lXFnIYnlDufKu9EkbBVpgMfUKHPpQuMXXlK8F1Vfi6OOwVy9FF+rNKtZkG8xUuzh
g8HPmSZLtlEvDimPqIEzimDvOmSAEne0QnnPmzKGUF8DIIpGXFn5Xn6EnjAbnNy5HSwEeX7MCAtf
CRCAaPFQONH/ra6zFsEAS7jSYaEOPKFYPAFJY7/kxDOtUD/YCwWlggMSvAmr0AzvakwGXzgyWy4e
H7AzxD20eozpBDf+qblhm+q3PG8zFmhEslGlLydFb5aZyYWGErP2/9M00a+lBBIsApAgxXvJo3KB
yeQ4dsmJnWdopdvciCPjsaFobcWxnrT0/wgUz3Oc//jO2kbzUO8bWFfTGnCBth3As//xacK7SDq3
kpwuXbRuxFtnH7XyUfgG8v7U+BiQyycLnzdDxf+hLmnnvU+pUgCxYr6hTtBUV5m3rYq+1V42meoC
SzuSnbsg6hWZ4o09nwzbQb0STjftZR4TVNafrycLTiLTAH57sZkpWySukXzK0aL3WKAkQZrUa/e9
ENzFcKcLrsYWwmLy4F4FEi1ZvvFijK/SJTwVUbagtLBcumzIvqSBToHO2xd45uo6xTIand80ktgr
RGa3KnG1goqspbYjfgE+EWEeitgeq/AhCMzgQNjeLn1MCYU6t2Q1M9FqF7IseFenr3O7TRAfs4qh
U+Br3W7QHtcprpSmyC3i2D4O1mCxOA5w/yu53V3JS8CW8/ltUw6mOakKa4jh/7TADPg8YnNOF/0g
WU1vz8YDrQuSxJ1nRmNsQwr+KlA1uyzD7OdrXlJugZnf6E0qiJbLLq2JEFusGlHL9QOkC8bRRNhN
3shQiY5GBai88WLNK71XQRFYjZDk+TXfC7TFI0lKRf3Az/7uznc21ruzJ6MwMivvtgF5Qgm0o8xE
VFQYufwUSJaGXY5Fb7QVJ4MC0JHbU5g/MI3W8VKnTWrFQj4//IOHCbQYNK14ToTbuYYTOufRi6B1
NE44kXPZiXZ7bVsPx6XR6lbJpRglGBmWisRc2MRY56Etsofxtf5FhqYpddGmMhtAzJZn0aceUZ4w
8yDi1A/rc8FmEgh+xn7XaHftaBwSd8A4nQUCj7fScw7BLHJkRsREDcx848M3bXKyOliEEWeL6DiE
H7INwyc/QCUh9TEprVkxznEiyrRQgBWkW8coH0JF3r2+2P0cAp5LccryHX0m/+NzrC9hCLpdNTEW
AuT1HUHGln06W+bGuF4LAf6ABuq+2jjz953/g0JTBzi9dfZuFZmf7XfgzwF0lPV+1gqQzo89SFiw
HDtlM7jBBPFnm6zXzchyfOdEoqidNU7yB6lEiC1SuTYN+9VAltoGfLGR3H28ta8sHTCUgP3XB3OY
mEmp0IwmROOMGD8c97+1mdfyRfnbG5b1w9/a062Vi1HOuMb9eyAmEPYcB/9svC5StXL/5cF+7Ljb
uZD2uiYotHMzW7QfCEBBqJ6NBD0ExPXbTpA9T2MURJoo47/tpoOxGzjMOHXfwr4CAJMvuCkAJZcg
nO5hKjZNSqNzgBTIB8cUnm/VhziWxp07qlv9V/WC9iGD1hzj+jDOiZFfGxttMHVyf25utd3DzseE
SQokhLxZryXdqSVmgxbhlY1Gs7EnLIawpoZSG048nYsns8l40aSA6HsGHd2Y4jEGm2lgNhSOU31v
u4NX8Z2urXi+5X05C1XlYwpJiCxeUaC/17bXxFCXbhry9VcBN5k+L3E8B6EmwgtFZK/7ltVOOXYl
6BcxVnPN/CNW3evbIm/8kTKL2SqOMQtiXCTy87fhG+tU+uRWU5A8BU+d9oBPOKeK2M583YkPM9kY
xP1yuu2G7jZ6z+Kyq4Rn/oM2Gf0Pl5Hmu0+UtsYMDuaZNte2WMuYPT5lh2wwZ1AhHlkhqtG8ULjH
jyoGrnEsXl917A6iFmqqUpLhLi5yHFaZoO3LorI0c+FbXojzIx3a8Fi6cVrQVHV6c4qzyHPi1Ybz
HEoxk6ZhMvx416biwax1W61ihU2+YKsKJbnwwaZ+bGk7XPt3u+VCrVEvI/ISrTTZ4XEpgxharvwm
yV1+u00CHUWwqtLVCQjAkpYv1aQHAAEfoL7ijVUAdGBJqce4wvqZWFH2p73IgElgB+jtEWzU69Ex
jkDgfHmVLS3VkI6k9lhxzT93XuzQ2DzTzH6bKU/IvGs+Y5pnRZVAWOBEjQYExiMlk5Yfr29j1Vn+
4T7ZezRLCKeBTVq/zfw7OD/zlocki4IGTzYq89D1JBnnmAxiSzHn+r6gAtFITrxez8j0mykT3UVp
5PM0L6sNzwG6RSvfn3m0SSNN/oOzNkdbnBT1TUjT7ZmhMVxB8ZDTLhOQzQSJY2NZat5ycanncBLv
rUBTlXOpZeGx6NTZn4WCGQAzr76+BYZ9LTcK4GdREHfs6QYbpZVMiPnBN0k9dlyc+pSmdxXGe4s4
tMio8VxdvCbUjPHNmb0Mh9HJgTfIMxf41DLBwpmFZlfmR7jqO8jpmQE02lJGT8aTLyIIlpXBO0zz
Q5tuTP6v24HvnJcfNbb+4Yna58x4MYTlp2zUukuKPxO4SSgNYXQ3Xy2E6nsVxhu8TQRgxbupEZ1j
9unHtzRRtyAO0uc50JUu0KCcSui0ELlcKjB9JNQdap8A+dBllI08Msq30Cn1gv8rOIEJwmPdjZ3s
YGOi3pImH81lzzVNlPYb/wXMhL1mcfgIREm/SL30sb0NecY+mt186yUxSFzt87oCkAtdLqxBE6eP
xCi2eGN96on2ZQyhVmuxa5OocESGFuclfqigarmrQsLZeIPAR2YomusWH4Me2ZlxQmTmS5ZrxIv8
skmoftojC3Oet6DZwYBHsY9We8XuY2pB1iRovHk7FQg2M93Qk9lDbNDjmnCLJtJCWaVmzi4jBJs0
6ssVJsuC1E7QaYIBokEEENsSaf/iNdRQttGetyDWLlhmss8QDmDZb7saykA+9aEYTCGATk8mwyMT
cn76qRvteIagXHZwtNuhubcnzEbE+ie73BsqRFpZGjFhso28D7LLZKgO4Aj+WouiYjcZijZoqu1/
08hwHZntGjL62MFa1aTgHKX8Pq6dARzla5lBG6pjCnGVGHiTHtLeYvnqkINqWd6uIE0vY5tMC0vA
xcDLkC6KzF32Nj6bv+chUYao3R1cjL5hhyh7mht6kbHjGRYO/Ug67w40g5hNEfr0vd/vN+o3mWS5
uH3UtN0pCSXSrOecswoKXf3X8P6M+tEur7NFwoEpXrBDjgTIdUqL8386iEI9GFoGKCGRtf0Y8on9
lp1Pi/H28cNo3gjr3WvYVGMDT6uGASCWNnsGsW0BOz/xkGCIvo57sDAe2P292EApOVeVzp9Kowj7
61iWafP9JuJcw6P9Dw/WMZ5PQKpbwSMUdGnAAf0oZnfR96F/RDNEws0K3+8kcJvHtGH3UBVni/Pg
cJbrVsoISF4j1g8wKfQ5e6UZhBeRFu2awQoB3wkxFH2IDw5OQ6CE0Gf5nE0ISHh9tlyUSEaiaVhX
gC87tNTe33vIv8kzPgp/piK9joOGubUv3UI0tVB7np5aXrtqpIKYLJxEGPEyXEB/ft4jGJUeijE3
ZYraKOYoUh57SLRxZdznRg4IIcVF0w76tkUdTLf9U5BxHhPWtTVES1Z3g1hKX3OSZ229TJZqujRC
TtTC/da+Shx+tfBw6OGpG6H2azEFQw+rweakIq4XhAMvZDukgVsjna5Ojjj0T1i7w6kXwiDvnwM3
dm6dLLfSgB93OXmhhGcc7I+MYaZMxVhZp3RpuvVXhvGQ+GphdLLkONFl8QdnOlrmCItGrrp8qEXb
bZfCxRxfd1J/pQSXCIZh8Xl8+zr5U5TUHq96MjcOKlJwivMW9m42p3hPZ7UeeOVPrWG8dTMNpCq1
BHDnpgpa23iRbK8XGiUEAtWf1DbwcIbbBJ3Nesxc22Kz+ROSMBrRC6FI/Pyxjg3dfdgE5RZgb4er
PE7PeIemzSQbG1KJk+EmoLC/ngHtaxZq0Qcwzbh3Wqpfi/mEEmduknjGCE/jCmUrur95WuPraGh9
1yxYP5j4IFY3cEDrAz1QEjYvhddivVvVykAL2weCUjzi+9VGDO9CWpiBt8L1xOyOgB4qYzv9uIaV
+7R3bGQHeKtj8s/u/KCCxE1LqQnqAyFHED250Z9n0srgH/IxydG7hbnoj9f7luARYgL34awkyQFt
tltY4EiFy13ytZ1PMlFMIXV5/B3thpl0OpvBRPAL+UHd+JGC1Ari1gk1ocbi8xYSOYkGXd4rF5G8
UZI5Wn3eZhgzaV7iWGOO8mtci+iR/laNZC1oia4CoO6O2LgRd3KoQLK9ZvWc13lGxL65sQDMKbX5
in3fwaduVlnbnAnDr+DNOemMAlrgM9rNzi3DKmhugEi9Au4oi8sedV7zYJ0zV929siUBGTcUEJ9J
a8Gtx6+u+LKu5xtDTci8u++j7s0QbqUSFwSlaQxJBojJb3xW3nWpwPdgHt3+bXgm/bmTVojomw2h
7k3J89fl4v+Sv9fXnilVARmfGWdj52/v+5FWOESc1JkYDfH1L4MPf7EyW1rbfFgtwfB5ckocxRRG
l0xP8yxBMqhIkgDKTw9BLC2bspBGdkvsC+4duGK3nAyk63po/OVgA+A7GYl8brjyDA7777n2+NPd
ROypCJpYwSM8tbIE6DFpuB+9ojR+crCWk0tgWEAYlkDnzu0X1R5C8lDaljk9Ik5VAH/qUdBxaCXb
mkOipd9MRI9mi1mK+h8EKsb/I7KonP9Czhlp+9BmS3Vdk0BDNtSiA/fsrJIOfPSJrAKzd8JPOgxM
0Pk1VplW7x1Y2MM4qQXZJxYMi4cbavV7NiqxgjXEjEo6HynZe38/DZiGP7efFaQhtzLkFvipMwfA
qyyc+ml3+PIm3DEiNqQojKmQmkmPJwuQ7HrGuq0h+ViQ6O4bcFxiP1Tl2QBmedNA6jxwAtpO/J50
eMgRNjmgXm4yaHBGQTmSeK9Glx7lBvo4YIigfUlCVkDllaH/NMGwfe6E+JrxZNPe8oVWBRy/r8wU
OnxF6wJHBgpGrcE5e+iSibMbH64ei9x8xHT8ha4DPfrOlbokZEpIdNpW6mGFWmHiR5hWaGreCkqu
z3e/msRko88WYKSN/wV64GKM6jYGXAZvii4H4V+FeEYpnBrmDJl3LwV8vGicUJsLG9EaCFcGTjTi
oEZ885+QBCfoJeDLO7MvltfLXAZ+iUwnI0kPEvQCqFEY4x8gvJHEyOEOB36Fxip4W0OEhOkahC8a
0KC5Ud5A1UgaAHAf3PUgP4pxo6Cr6s7y6I7uU/jsTcIwZ7J5wz8IJTPROwsNMhNMJ2XoYHfTUkM+
Tq1hmZhZdQRM3qlb77ey09oyuV4r7nyEsjh1g9DEoADp50C86nziwD9Vq8BwRum4AMeJMSXB5+m7
QciD1G2OPrS1rzGPrNcEXNEkd6PD/UfGuMA/LBQf4DUX3ttyk0iuLPKHCxaRj/8VRSF3h0vdnNND
6GSgR0sPdqZrfjuQfcxfc3KdKj7P6BWqD1Fy8UC4KdcajqNpJVdtQPb3tYeUnzOoPCkfJBsg/agt
baWDFO+lTPWmmoiMCFXG22pOLWVjSawIrybbO8kACPADkptSHyatwDARNp5XefFiJfdwxpuP1THc
Iw/7IlytuAuWpHWN8qoqRjVw2Xq1o5r3I64jJdrEV2e6d1f0TSkevRdq0b2IzDeOw0M/8+3MS/Ke
OCPU0UN9IaKb+/0KFihe0JSyuZtukIc6VOmsPjjB8aDF7SoS36ZHfZTtXRHXVzhNrWHVk69U3i3o
vr3yfzfwKk9xwgCQPxlTrVL04QmT2IyvuSaOHsI5+h8wfnE+0TNXR9RwDLVMj0Jjqh55yqBdsdCa
rTNpmsb8XZcAlK1Uiw4E7uG+CWhOsTRdrqS1gmo5xeFVfey+YdFEGLRcyGL26skKQrIRZZxgfNsg
5DPygCO34UiCyy1gsvgI/kbkvEimVmqDA+pKlD5VGiF0WrZ2lHCS1iRlX93V+BQ+/YbiXN++ZFA6
ymY/aN9o3MIXvqzW7+UDetneGVMrT8yz975c8wBeIUDO7JBmYKBlgjC4f8/HD38JOfTic6bCUTAb
+W86PSOxWGXirYZl59aGN5t4QCmRNnMzUdU73CQ8R5UhqDb5PHz3YxjHYryT6IuqDLNJfmPjLEb4
c+t524fMr9+1cehJSWUdjIDdvLJTTGcsNd4PpwGY8223ZkgoOPQHSXwhdZS7KcPEIVTfC5MCx1Zj
VpdoY/NeaGw7doXcYlQ0NFwaZCF5B29oObeuD64sQhTdUUgvdT7V+uj627SIX3HtpcJXnKsHMHCh
ua+aH1UEp5OQUscuxECouUmP8LKgkmQn4bGXP3HIK6xX6sDYNV5pcTsezKiNC88CseGKPy/w4/P6
DuN0qshHlQ705OrE3CNi6p0NV7c6cE/MVwWRwhReZxnTrU7upOjYuTW0EsjA17sfH9v5wfDRxYYP
syXWZkWrArAAy91hgCPNxyMQ6TNOAA1UweR39fZt3+Aw20+vxr/wZopFF/76N/uZdbOGJaAV2If9
VQkL1Nqgjs4nOJ6PdGi2eoLd5DfDwn2B3eROjBmkMSeBEYhxSEzLL4nKXknYYHdR7e4SP1JVcSNn
o3OkdVtPseQypl3SUXiDs/Qaq8gIS87krH9jKRR+exLHjcCTP/j18yYNjNbwP6AkEiFiLZiB9nWA
jSpM1qPUBpML825hpdTh40OJq7G7Re/JpStitCA2NJK9zdiKw3VRrHG3AbNlwQGvLgrUFf3FNUhR
yBZwrL9duJGzVUkXjiZ9vTHkrpJFxPHBvWKo3M2VkajUvQfzyeGX7FFfiVZJ/I/YMuz0q+f+sn14
mf4/wHVNlW5+4Ncle0++7jDZttmLnDNBaBRo32FH9Jt/mZmKaLLHRmQ9Azit2hvxIPCBXkYXKuJd
FhPUYrHGUiwgTgOBlJVF3phuVjlt04NDHFBlzv7A5UfFQanjsJV56SjvkZc3R3x3jEc7uf3OG9fk
JOX4sbPZ/H1x0H9HRM7Bz6PYMVcg4ZjCe8E1Q9TZ8WM4PeWo2iURnrNM80OcyLNYnkURqco22zXq
3W1n13bV11T1ODGPiGn1qZeoqP1TPFMI+kYnfzc9Bzifc9MkyGDRV0GPTz5vDX996HHpcf4V/h8Y
gENCAvQmY2RRzxpiIsn+eY7KarH5c8t9QiqRO2DddRsCdPl0kN9vOzh0EvWDhEzrVr9uhQw9YdGp
PO0qfnZIzBkqBCmgHCWIwNTyj4fsstgunWWcoYQDaXW/F4PGcoxUsHKhZ2vvZGiaGG4gAvZEsPe0
ftUmqSYKZvUPQFqY1gFQzjV4up66ItxOdDZqnfhcE3/iMA9EomygukXw9kPSHp08ppBnPf8UqV+z
To6NbTmBk6UcjAOzSXqeDCTs8ePobR8Pb6eByVQ9Nf5NfFoq9x/OvGmZXR9sPkkUKIOopoe97GEx
NeXssjGXT3vq21/pBqTlv6oZfR1Eqtj+e/yOLKx0t/nRb4jBEMxyXDu8mut1AxxUaZZWKm0zzRcl
oaMtR9ZOOEU3uiAVqFkPfiVRwmfly3bzJJbU/zlw85Ah/upOJqpisWg0bNTk8RWdRILU5QBF9v4M
XVZmm7dpxl/z5K+DflcEqfXBc3uW7r4rcIXHOM/ZPQewhGc+/yZjEjXP3zlTRl4C0+JiQQE5wM07
EyUD9OXe50YHd8pllCdAck8U1K8c+upvS8fh0V72xoUiyzLKjk+LNH7m9QGOLgF+NejuDcExYRTR
TjSpl4N38A6qdQAJLcuMpBWHxScTbMUc/0RXMmg7u+PSgzEIy3jTKH1CRwUzLM5E9FjolxPGfBuq
PP56O3Ralkd3RC4tpMP+8TPMXdUkhPzzcJMT6s3NLXT3oLc9D3IvYyF7SXVQHJKQAnx91Wyj462R
eHhYDjL8T8aI05W9ggL3Pbo2Yyx+zbadBMoQ+zuc2wRzjdM/aE7gE7HGo/T3UKXJC6X4PrRMqIH8
cF4/LzaFEXpjj0pzDXS1itOJkFUT2KU/QOQavLbgIaZsP1tLZGENRdC6k/NdpVv9c9d6lrEKN+gE
tLRPWKlMoP8hj+PHvZ4ka6PwdMEI/O/Fb5Z0MrO03Uc5W+T2tVHRaOu9kYUjd5JthWuQaIJcDoxc
PzKzmDkKzqaZN+6s+2DWuFl18lX6lhf0D9Rf9eevgu48vYwI+5b0+cNYv64uLql4/8pHDhlRyNV+
pjsHDQ4myh0keeoIlZbpoMw6+rfo/ei6ur5MDaDm44BrtDcUK1ZvnFekHG/EJjBfYNNAnCu0qbHE
64ctfItwf6MjgN6b/QaT79tbyWvaQtBebHWEpDHaBfwVQxHpUxkWJ03ymw4mT+H+FG6Sx6XfX85c
LC79uD82jR7LqNaxjt/OFsYmEgyyJNcVTffp2xHwyeBG1L/ATrDzX3pA9rxz4AV7v+LrUmNY50/F
CCEyd3ee1p5Pj+8JHfInKX86jEOlRkejdH+AXVGXtDGDssAh711T4Es7UA+8B1eRaXW/J90Y/Uxz
eKxq6Mvgrb4C+HAEO6VSYMQG/klVFLtX80W3ycAG7leG+sV2hJ4wBi+H9CwgSbe7YQEnNZNi0T9K
UGiw903fg5f38xy02un5jqR5UR5hZ+h7T/HcvZ7wZP0l7hFqOEqq2UwWc0qsRFBBFC8cNDDLj40w
wlEyfFVKzIO69yiEdy5NCbTcBlfRgOJWhJJv2PSz+M0bBoKSNa1ETym8Vm61mzx8dB6T371YBN7J
GDWvgOv336l/F1MKa75tLeItIK8gnS+ymA3PXgfNhPjZMIjEmCnUhQr27IJsPr/g9Y5FGyHr5Cfy
Otw0NtWnR4UYylYv+O63hlXraZyTsmZmea9dCNeQraOAO9xMrgeqAA3ZvVgUlZWdxdu74sJm+Qu5
HHUdt0I7Fm84yH3kEK3cuA9YQgqqw/bZ8PkdyrL/tF8MEDXxwwggTr6BDTx2Lwgc6bFOB/OibGkV
wzLpH+C4mlO1EQ3DXe1LkhxOnvQeNqeobfePn7rlYz0HGFX9sZvWRqkAsb/FuRXnEY5D/EL5m1yg
B2QpHBdW9cJWu4Mrupi9zndMcMOtWl7HAMY/vDqe9dSNq5s+oxLAlBE2GQlWwpwQI55yPbhCdwsw
7hc7H188H64QvLFizkuQ7YGDf8/pHp/H8gYiLzqCACLxk3dcU+LmR0B7lL9aNd2yLauMNEvrZfD3
sjjerLDTbpp24y1HCyCT/2icMR54kJHARWM1g09CGUtANUYk7Ugeq+WcyXkkA7Bb0O4fuQrH10tO
fccAjmwbQCDh/Y0XAxTC2PgB2L7UFvdgkLMujG3zPI637wxv1Wt6rTZxiVJb+w5kjVJgMhWGTT8U
JrcUMmuAcR7creVZRGtgN54xqj1aGW9m0tJRPR4P0kYNdFYZLny/C2qu5mRwt6uz2Xxtr8FQp7AI
/FVwoDhlhgSsqyAPjGmM8oLbyW7Et6pOO+flFaBTWp/BOsgy7mFGIk6cO5KyXTI2XSR70XNmhyHV
Tkt9oVFZ8u1oTCHsq9i8VyL/hR+GmxR4GBB3RInWPcWEodpf/cblH0tWDfnocjZ1P/oYZ8F6Szem
+h6to6gAJgy6QGTd1JN6T6+vAs1LaFQNSAFNSwYeL54X6MKYUPL319H/cGTfzq4E7g794FdRcn8O
tr9OHH08RdMsT3zrH3llJ3f5u/Jy4MMwaLVd4LLFKE1xLbXL5l48Ljo2oMk+TEDSij7Q3WeOE6oK
GdfmK6Vkwa3j8bcLpnkdrcLdqFAA49Lu6ij1tQX2IUri0irmgMiimlWTHafVwNvyIhPR7EXxX1VE
wwv8oKyIBXGjoDU+vMrSd7It+fJ205uGj76N0HiokZGis4OBt9c1A168LWU/1Im8h7CQKPPyL5ca
yT7/av0DROvzV69+rT7EmhhSLbWE3WeHh/GmYQWdL0/IoQJ4dXXtHDwTQeYicp3YlniM6CDIgEro
GJhBkgfvWyznqmIfFthhRm4Zw2g0jBcdSs9cHtqdRHYRn9Rg7cS63Ovtk+35S5s6G8VL4D4Ub4Bg
J7CVgRiC+37HdOkMvh51SKeJ4SHbD1R77fhqkInJR5PB2zeaRQxhE7Sby+rtM/CvQU8tTqAuht5L
P5L+QcuZamf1VhinB55PvyhHLhBNlG0SqdxOk4UajahO0y2UAGvDpjpe2fD42X1ME4w3nis2+PGF
DGCupz3czMOX4Tk2TpelKdBgWV9hPncla3D/Z4AZrSwFTGS6hCdq8fcnSYyz2dn8olcMIm3J8Q3B
5K0IHWDH/ZgsIJLnY4hX1XLrJW+wKLeDVgKSVXkhyq26nVp5f4ATJ6jsVgimC2AJhP9CPTp8PJjC
BkCcQUL0QTjil0suPLsS7KbquOucfHDiP9yC3mOpzSIQVG/J5U+Tg87zbPHcE5oxmL6msL1JCVut
RYjY7GIuyP/O3+hv6uSAfO3f7lSDoDPrtWKBTvbKbresrCNRv9x2SgEmelcYd4I1/c4EFLRz2Bol
+KSsNMpuv8R4OeLoJuKczsMCkZ8ZFhH7M6w+uCf/cHcZjroMwVltof+0O/pmzqw9wJ3WJ6Mxcb5B
yfj8WfDHOkZ5wNL8zuQQ09H0XmfPk6seKfYviL0a0Yb+8+/kCddo8QwIgWn+IT1MBMX8xzmrILvB
OcHmQyJ04AeLbIcqKdSubiZcttJBoMRB8Q4HnZRhuLlBz+ef6DThtgxZtAu2AefSpkkxc9cb8cnz
CmRWtT442UOP9tc2XinDY77vISPIzviORv3zPc/ymBEg6HCjr/zc+k2vTV6NN6cHbzD6/LITXyOc
buTkn66yJRa88cNrCTpX8yD/S4KI5gGg+VP/IbeZYwfhPRQHJKcN9eMS56xDA/8CCkjxuoxuoxn0
GzmoEh0sFhphlaqg2wrZBbt8a732ucXysb6e8ohFBOHfZ+3VyIrhHDRhHNCMOayxbUt1Y5bvIaak
lwgHb9/3oMcfyiJ2om0Pwr9JYegVXUv4mq/b88m8+x9W3jPORJ9PJFFIC1uMZj9BwfOACMxGjU+4
4JSUrvytUZaN1lFXmy+59vAqkHZHV3jKEQlaezvaBKlAFqBZf/0iWHtZaDWJUrB0YPb0D5e2KKGU
6d6Hiq5VsuCZ20HusYqJZGHvqauZYr4Ak1vffIDSTOUMfibyXBicYRNyTxqZI+vzF8v0tFADV46V
YodsA3DJk4IAuBWQ3Itc3o9QJ4r6Pwhm3noIQ2XFtUzm/Ym+0KTP4Q6RZSpCknAPgDPbFq32bYqI
jfryQMPYbL68NVXRlWhtCZFTjbxqw6oZNmZXGOLP8R+KH/NcbG36C5zxlCs95hk+f2K4mQNCAPTB
U+1szpkVdMZhgkSZ5rFFChLuTVFgO9yjDBuf98og6lecTQi6CfbMkAmbe2KYbuPlZ4MEnsIhX/Bu
SgFs5frh5jfAyohhUW1JkR0E/w1rz014jgYlToJGT9w6OGtKuiaUdgoPNzzuiISSoD63oY24WKjs
NaFnnZZ/hobvMnlBXmL9AOJVvWcmGyGfQ1tClaERY943skADDQYykg3g9zHiz4YKeVcO8XDyoeGJ
8P+rT3wN+eeURpF8tFErqAKEtteclbMtwFXO2dWj1T4QVYwqs7ZkGy3KdJHiOkhZCvKVkAjT+jpF
vqpB14YMwJCAbyJiC9IunYHmv1lPC8iE/siL9Og+H6+TokoNd2Ep/YTeJ+fJSOJosPP94hkoLgXn
DrL8Zju8yzPFleqnjkFC4W/1IYaOeFqUfKWzAf4Bo8HiNiw5gnGt8IgIjB8PSQecN85Gf2VY2iG5
Mpr3v8d/VaLV4xiS9SqG8wipAOW80d0dLvhdMNECDDwJ5OuCmI/mNT+vvnxnGOPQp9lBMXHpu6cz
FJ08PRjU5XuXRaxBh+gnTmt4leYhrF1yMMyiOiDTxRw/cqyIvddBcKDaM2MMxY3YCjJR7N6ju+Zv
cptUNske5idDtegvWjWAk77NfuGtzoHm7gNM5m3YamfYZCnR1iLoRzOsg2yMCgbpJdpnbUzGftp+
Pfc8z6YL7j4J0pz6rO5fCt35IW/ol65LtmBBGBX57ZLW4UoK3YXBLYH1gY6eSbelmBqN4ibWydXI
N3+cJq5zBL9Txc9vbH+AOJv6FM5KbTCC4sR6AN6MRRXOMqCKH1nDosEvP4DSzjSceCqd6z6vU2Qq
bgP8UC2tgQBz+6wuOw2+wJwRpDjVetZRuIt/Q2rf+seey7dl7t1n3lve5L/Z6FGkeFbrqqxeHYfD
ovbXd37y3bjVA+4vmSrDgdafcUXlso2WoXHImau3eflHlI1G8gW4q90Xzx7qDZn2zDHD7S2OTrfH
L3cJacYQiSlszcirZiEmXGKvE6ZNWnvq9Af4+XFkEEfef7Rn/MDVLXaPRpoRKvTaGwbiWQeyaX3a
goONxAiSGP4Ii9N6HdPdDR8vPDqXJgBsI4M6o7za8dxToapeBxSbrhh4EIznuVX74pn4cWPCjQhE
tMncuKYgk6r6OABeqCrWnvFwX8gIcpNZtTzEH6YhqV2JHh5kezIt8HmvCETUsoH3nX7/0f+4uyoN
OJ68q+ZIwnWeZQMJGjdfS///o/ZDGOb2NZB/x60BfdWKiD6VXOq5L9giklBy/zvHSdmI1zB2jvdd
/a6v/TuANsJ+bDRc9X0FMFtkdXxrQCrp91HtlP/AIx/x80H9N3cQoZBo4BKRfLYzwb7zRwgLZ+yE
PbsReYkHERaoFIhiy3aPPOeR7HGUlf1xtYxoz86mDJpiddWqeQEgX/teWDsTbqh6ner4MV5Us0/p
IECUKu5afMBbugjDKFQg9RE7PoO1jDkp9ra987NVWAxDa0j1cAVBCpGtJybOeV/c2E3hGLr++rCR
5hBX0+zJ2yfxkUxzFDgWKqKBhAtuB+ankQDqBm8Eii8UAZ5QQtTBz/RlzFsRZsWVYE67/LBQTtrV
DS25wbP0H6sPvtqT4yMKwUJu7ddwnJlSPaw6ntrkX0SCYMW/IQLm+ePuqESFO5vzZ4axhMTacUjA
3sTnhUpQWR8q5sEgKb7QJsE+7PQkV5xcHTMjQXmT6zp/mLUJ90Zej6m5mE9xenrJH8oCqYFJtvkJ
YcggpVgaopo0cyDgUiGv7AALRtimbrINbc3E/yVr7fZ/DQvJGUIkAbtLebC1V5vb3oRuFNsrrz9y
FHvbYDOLZWbMwbVmo7v8kcbesMO0FTPgrkjaWlfhta0zXQFat3PEdy7G+sw7QLrqHJzw1pEleeTl
kM/0stRwfzAbdkLxUcE0lTd/1CFPyruC3iI5O1Ap0pqOf5rgIIYp/vTc4up71JIEEzy/xyvFdVp3
w9yxp2574GYS/m+uN5zejKqlU8P2E0OWOrGRZUBVpTFLaB4iGmjEOMGTDt+ML5xDsCnQyapZWlAt
8LYPqqqYtxCKoRwUFI7dNaiY0iAkUwru2Jxyh+9k/SGJh7rVGbGmZSGAZbUGeXjjGdw2fRGXn2Fw
PcUVYYfHEP4NsbAVFBz4SqqEyy/UhxMgFBQE2goghHWTlzH3udnXILyRyf3+56XInxNJ5Fqizb7d
OQp+oFstvxBM5yfMp4StxewFYe7tMGFTmtBluvZhkeWddq+otC0vDIBxsKLX3nwgfBY9rEKmZ1Rg
CbzgONYYg1ziylcnfkNLeozTVTGteIOQLT6jWxugV/NQ+rqllr9ggXtfUZBoCyJbyZvlZxcaFEtv
68IhaoGTLoOEoFvkik/tRzSDgPcpJatjpprRVjvAq9y/xje5QF4yi3NxCO6iZHMmHLVf44mEcw3D
bISsQJFzC0ZOZZplLHFXV8wbBaS4d+4TK2dg0c0n1vJ29/Z8D2nz2ND/iWVNoV1sWHViQPnK/9/0
635XocVMHiNInktfzKYUrMcsxYdfNFJxfDz3lWlmX/kDWcqGIbIjmklXivwiP0Y/Yn1V80mBa774
63QnxMovkDCda3q9ay3MHils241p2Ai8V5FuhxmnhpK80ULukCK5RkmT7ZZtg4XSn5KupXQLblb9
kDUhXbT85i6J3B2U4OBqeXgnOvhksyMOwPNPtGd6UTarD9+D4MHAh7iDsHYFVEfZza9donBAkRSm
P8+UWnZiKzjPySoZMefrZSgve6JyQGn8eTOGwjv+bNlfSw69uiP9KDqFpbXD36If3OgVhQRpfubF
GGn/KR5mNpwH6/Toy4BKmRGmRkjCEnchp7RK9yXd/CBunkirHH+Oe2j+zbzRbbnbjD99T775O+Wg
nftlul/DHRnKZ+4ePyEdWnDBWYaT339MMuTFojyw3jpniaBqArOa+WM832YbEKhud6xnPZNDIh+q
vqmX+iwgmZ3etwyh8eVwGM7RGZG9A7LBgsyasFiIcObcZ1FH9Qt3FdAO70avXFpJdhiIQzFZBUyn
+/vAdDLKLU3FGSQlDvhsV9SnqMBpMXo68fUq+tP2KYRuYVoB1oXTADs2Wkxg13K5kEyw9mX8pDb5
3vHCK77SdRI2U4xTEPT+O/CWt0vYmFaO5PWMNE4yLjK5wG60yNOHsi6YKkPS8Z64+n4ijo7qeYZl
ODNvB6KvhC2ptZqHNGhAjwv2z3Y1LVg2l0y2TdYnFjlrsr2R5FOp+DGs0m0glwszkAB07XnrEm+H
DCoKUkAWfzGZJU9nfL36yRQAHAF+zRgnGcam/9ivQk9kxYJxWr5KQvJIWggAE8v0GwNixQRAeJoz
ysOSj4idQh5Hsydf4Vp2WrC5Q7CzTbOS7xqXVWWT5JGdyHHU/S+/MtLc4eTSsDVp/9Rf3lkCjb+J
4W/C4EaO48E71aCd4arHWgc6z9hyZNz3k9CpG0C3ZxoF+jl5AxqEFiYFPc15t3hpw0d7LZ9Om2jA
y+zN5Cphyil7G+GKkG0iNsYeaDKAnaJ160oUKw3FsiG1oIu3WwkrL/QxlNq5WUbpLZHSkM2Xwc4h
jucVbyVsB5CcVl7RuCqZ7H6MlJOVB/rHcBolXcWQYxL1YLHDPpX8vRVqvJXGsRTfqO1pMrYhJe86
y9itQOq44/aXlddJUatZb6aSrFcy3qhrPCQRJ+wjRLmQkdmfiIXGIJa0D2q77hP+m/ppN669m0WD
neYWwX1YZ8JvdUC5Yp5JYSJ+oM3TGP+hsl70D1NJaOsAIO64SUcjw5qV1xQOp1cZXz1XbJ+/Velc
ZZRPvckD25joqK7yhb+afAAuorhcOeO3W+hOzxcpHC4ilnSym5qLY5RO5LmI5vxVvGmbNMuSlTil
iJU9nEESMw+zR243qHqK5j4lNoJcqgvbElYWeheLq0kD7Hdf9dMXiKmMuYg710Cg/H83CwY+b/uC
AsaCgI4OngZN6pquKO7wAkYOHg56AyN0ANXMgtrGKCWFsJwg+bjX3bE/SOf9Tr5B+Xb6wC37MOSE
mKon3sybGS0J9inMkPV5TfVKQFnq4Y6B8E1aEd7rkkpBarlvNiTcciLDUuntXorqpeSfI49lPkX6
GhrlJmUo43vzlf1BAXdDLAGS+ZuEvxxppoWZu4eSNJRxLHWUpaM/NWDHL0ZmZ5ry/croXWeILYkC
c3KjiRnrZ1VdvOdKeBh/FAsqkyjzxULpfep3VmvLoqHDBgRRiQuUHbQYgwgjnI4JrUDr6c5vKajN
7arjnwvE9SrE8tz8hTfCdpoYljKZkpUpqrb89jhiSnJru8wBnPOx3eb2vttyxJpamjc9ZNBT2oRZ
sraYaZIvPKAxElG84GkwledwLOoFUgIg0jLv7oNEG4oYaMPOYY4jCDXPAnkivtY5Q8q33XVej0Cj
Hg9pS8LjBEpzPSTdCItnKnKKEl67ZeUm9tMtOL8HooaGUue+Yz0dW047qKQ/95Vf9awRDEqD5Lr2
EpquWzhsWbeIV3dwu6tb1lAdWCvyUivwCmnlps3GMO6jAygl9+bCVALULa/fiiVSmtdMusUjSRN3
3mf1VFVK0ra2HnWdfz6oCCmvXgKPnzlUT1uQyYo5Rh+iykJEkBy9IGa3YLhh4FMRaGGysLobDwcr
/UvjIyk1z6QrM3D5rfQa6jsoFCsOO/hmd2NaNdp3ZigQaNIWdKIJWPEQUgHUNdd6SBIK5fUcSK0G
HOTCRZCCD07gwbuBjRpmFXrpBqm1ZdTDlv27DIhICEZBcf6ePu89Fzyx9DzG+RC5delOQrOdNdI7
7O1y+pl/neUKgnfpYTUsQlejGyqFHxi1QbTozmIeXWnoOEh0ym9CMkcFPbclneMSk3FrfjJ/6UeR
hfnL9QGdAK+ABGCWwNFyguOLzPb/CzOkIpUu6rLVnxiZSFcnTgxIK+acj4I73J4i7r23hulVSjgJ
cKZTSX/K03GH2i5pVkDp5uzVyTDGt5UpEQDN0OEE4wYQmkHYSD00CvVNwbRbxUUv6NyWnR55xPma
ImNLx0FYq3C4Jd0b3B5mdimgqoR86hVyxDqhr+dUw6KVDwwTp+v5rIEDq87eBRIWlG7iorfJg2wB
JkcFrGaEPxcP2MB1RTJYQa2pR9iMdiPLvTSdl2PX5ZXMesnyIyeeZJ3asP81BHBLSau6O4b8fm6D
zz2CLI+FIE5yAK2BoA5kQxqII5INkC4yNf01KAOTia5VB00fFBcCesCRQlMWC0sVaV/gciyKG2lA
WpJXTG1nCNAowraCwt3piZVQRhD0mft3O76HWno6CMix0O7cCGUPmGWRsVuS1Eg85vJiUhH96qWo
8NIwvTiIc+PYGVcywjPxIdnOKiG1GJ56Dv1/k9n5fgWAsBlUUyD5aNfnD8OQI+UebBxu+vXWcm89
fB9E/4vbwrQ/aAC3sCHmcXyWOxya54tGVVH9mhp+f0SRo+PL0p+sEHE34BVUzz2MuXfcAHxgx0/w
qLqmRL0sRRtP9k0ikOm7SsUfOaRTbRkD75twVmI/SuId8nfz7xHkj7KpjM+Vsvk/zew3rDNZSq7J
D5e16MULX0mm5+q3TxbRpdjH1tioSvAMKUEz2yZeR5oLZNy4HLv/gG+3+L8xWMxnnepjY7q+5FPg
nczjkc//O88+OVoeSW2MJkOiGHVvoEv4lI82AQmyzq4NNIHgj8ly/AOrbFqsv5irp6TnlIRWPzuW
AmCbWL+1SU7daUUAwKa7U9CYHJIkBWc5ofpixThMycSOIWfU445Bxzsyvrtza0jkbu5GJ4fvPnzk
GhHW7zZDZhdX+tsA7sCiIYk1JtLnvNtnddmNpM9dPm0nYk6O0TZpKLygHcZ9MfG7OwF+yRvQTglH
p5YV8sJN1e4nKAh0bY2k58MAKINHAi9pzpH1Ne0vCGWA6/uKlx706mAU/DH2N4+KacoduVgwZOUU
40gpOUGacKSLszG46GsVsiX9lPcxLIYwJDfcOClbSyPuTsKt56zv2hF3WVuqbMwEREGhpTZXr9Id
YaS27yAERAqaIgFWnntuMPoFuVZCEIc6SfrffVQ2JZqlS23UqC7jxSgGmt2PzdSe8yCvtpyx4Bhx
NNEOxLdDET6yzdMRubCOsGJLcs3HfuVgrGcJa/JP+VnwbtCQ2IKGiDOw2u5OMQc8m/f4uDi0t19Z
C7r8fMuM2uo4O8qdiNQDdQ4xBpdsU7qapcuJRhR1hAjLGa1jrngtJRVwKWnqCLNd+wML3Cymil8T
Xlkg5MtDEya2b5Ou8CswLTC/a+Chmab2aX/53losNAwUwlCkiv9TGLjotcs8adsE6JJykwXCXxzR
6ZKRHP3JCHFMhycAviEp66tCBZeFG2EiZWp4PkDv9CDjCW/iV3gE83wtXsPlUtRiAvNPImUX9rea
9QWPqa0+mwMkHk9EBNtmhG4VtoGWmXW/7m3RaPjBryLfaBI1KHTD1qgTPWpI/vBrTTfXDj8EeT0z
kcCSck8JxkPQ6EvHjd0SS4U4PU1myrk2tA9ofJ4LSCXYFc3G6ZB17vOGwy66EArWw02/xoEmLb0W
k+wpNOxg7YkM8Dne/NOSdVV7EZnolrNTiUs/GUoW0gtmiq/xCfGfPsmJyVjdq7Z4OhZt5+7ezO0h
W5xP+VfJRvjDBVXmaNGYN7miOQP61OMJqc2wDnMJPCeGpGEUJuuMQPNmiWL/Ucq9drS7PV+VH1kV
drqVr29O6P4yEGvCcNeP8kKnHRFv3+781sqzHCpw7xKao8H/XYYxhXvFRNf7uxeD9vIB3a/s/CQz
6mhuVWlv8TsSE90MJDqIRR77VnuLVKTFjqoL9/zbNsoip0BQpwhzSd+vT+FUubdGOt0VhBwTVY5L
fzE5aExJXfTJTaj+t0OHgIRmL1tfWuR4N+ywphoNgaOhxiif8eli3sYX12VD9+pWKF+SXNE6O4bK
oKGMQyroQWbX5tv4KaysoVtrMwrh/wFDAiiMpNqvfRo2n3cllTWpyVcoquKO5C6CMRdIzOVCUQjV
75G0kw531BD4zpecQAr6ZSWcXLIyX7YqUL6FYi9tj24uqwEBl3a9eRrKdnvudNzGFVPmw5UXbSHK
6sjNnnyNuoeSjoGR9ZZEuEtLvD/hXIDOvfuZLKwojn2cXod0+iREWKzqObrQfQFhmQ056FB9US4v
twDRnXQrSy7Rh3+WqFsfIOhcO9FdGUcGE0M2mj78ySCh9xfgnOs8jps1EPYmSXxANgsO9gREyAAQ
nTGT1J37aCNs+rjzG6/vbkNnT/rQuwCoQftBrpJVPuhabUYy2ygi08jn9J0l8PQSMDja9bcGZLd4
AlprwR6iO2q9VlVdTgsUvRL+OhKWQithT1KMylbXlurlkO6gt5Bt8483b9WNEPAHx+2n5E/9XxHz
dolCL6tjkgDrr5egdpjVSYpHrHLSie6aU27pZ4i6t+ewfCpWjrYKmexH84+iGUgJYI0I8EqyJYTM
EYpuepOtEfYfCOMmiLt6VeGUnOUIU3efoWs9jHeW4qGbCqIAmANvOI2E7wKesRuXVTdFmChkbA4a
WF92wsn8N5w6XOzmHYVDBb09q/syROzydo1B7qx2UdHdT4HvGTQ7Xsq6YE660aGFMr3OVqyZPFZz
yuCo9s/zNb2w4a+GQsTGs1KS6uMfgFtBduxGzgVy/vTJbRCg1BLcHDC+J8su6xowuL+lxwD4PDP6
ICky/54tGRO6hC/UOzhgDarPCnayMn2D+RfOfCzKzGfPB5ke4Ds5Z7/dpkpC2eggG9a9ZDofutTT
js6qjhnfnM0IGLNyBb+/cds2xxOBe5D1433hrUq6EpCisoVyaAx/8FIyyovel4gn1u5FvZOLm2iO
peuO00qSJeW4OFM2AVko2MlqdcOuJiiP8FyMgx5863sez5CmxZR7QurJHp2b/LS9/CUCVfdoqTz/
nsAWTeSD79OOLWhtwIIFs+dizwjCBzd48I5mWMEviDqkyF2l5/1Pi0UaHHjtIisV8QAuX7OfoKJ8
HFAEeMA2vOD1xejvjiXbwcuGiFNzUqmtQmVuzoj26s15VKbqLoz7JlqA7G9X0S7YKvyLnHLpuRIv
t83Lw8g+q4Br0vC8KsFDD5RnxgHfgP/4BRQ+sRbe/ZnOOjk0FFFDc0WaXP9eGr2HuZmBvhPewmdJ
+H9ER9e5BG1buHwN/i70tGvOaMZa+fDq2HC1rKXgovOapQwdNUgKdjCptEiRBciYlb9NhuYgBH3E
ENlu9kZCjbbufeUM/FAfMtV6lIFG4I9ZS0yBYC4sjp7w42xTHLLcHZ6gevdOI0WT16S290dpL4Cd
Oe7XnVsagIUtl7mEURpGDVd+RhCHTuslmDjEn60nP1uLmMcQtErtfJrwkY2fm2ZqONDzKy1MhuV3
oAzsEu4t9LdRlv76pm2CtrJNpVHE1ZJ2sSCFxCg1fN5TGpN58xYfUHasUyoPuGWYbDnyON/Z7qa7
y34+sAQaIa31xTRN7ZWNKCMpb6yGYg/o9lHvC7ylPnr3oMD4Y84KHeVXtnbUMbkr1nsmDI4VBSs7
ciPvOcbHAtzBgoYTqn1BUYcUhbFEaBd6FV/1tY+GM0MpuAZr/7WWjCmrxeD4vUwCHWydOi+0Ltdy
6V2EKEdIbv16gFU53gt3Hzrf1cKBb3HN2YsQYtBtYQbNdy7LbeLWmFVk5oWKQMfPzLuxRR3QQdg+
iKZVaws/bq9qYGtS88VbsD2K6MmjRfhXis4u+M7Tty6Dau013w0HMbM2uGoy9XCYMYQmjvRXzpuM
P3gehQdeOcGwDfJES2tA2uZpw7i6yBZcD8p7fJeXee6UuKqCrnJnWw5EzHIcQ9kH8ZJYivGi3rha
MTRPgJ+QPDGHx+oFp0qgDvk502JHfgkc1K2dqBVj8rpF+5qHLBKiG1bWKRcvWVGwjRvvxxO92dsY
I1GKpNlmxOjF0H4eU+FoKej0SX52LkNBlRoqc92W/wT7kZE+/F9+oWBqTBUje3x6G7K00MvmgLNh
40bCIFERIFJgjVshpxNjMps2pCi022FyjDktE/NCSfQutf69E3fPAClkHYj6sb9Mwj3mQBLmLblK
bKLLus5mC8t5UXDo8h6HZ71fzMKUPFqkeAsXt6s622fCaiHXQsxhiIaJGfgqJfgkMWdZ1Mi3u5cG
b2j16xBRCI6ZYBZSXoJsRAbx8O7TQmRNME0UbBeJWoZHTgQ6Oumt2itVs5hOt/DTel0Eba5G8sj/
cHuMgI9Go4reYGJIhaypWcI6Ctvf97RbflyqnvlLKVIC4h2KiMpUM0Vpt6IhAUSaFLqhWKj30alv
xTtl4Ei1Bb2/lxeBOgClDWWq62iNppfi73De32mjInNCR3hw+kgFfQjdRGL9IpOSEQM3/JWJT3v6
cPsRI0JbliIUeoWTWdiqxJrROaqclIuiWVdhO4y+ZemqEEBS8bpAawQkyCdl7VL4plOdFVumvUR+
norw7WlBJsEfriq8s6JD0v2XbHAsCdeNCrwqc7MpIRpJ0Q7dXhbFGdFBSbYETNiqkCNhlqCWxA6h
zuTtegBioAWA/u8mD64uCllRJGmrQDamuMi4mALJJJ9uKxeaITzdeqsARGYh48rh3/xCAA7yBvz/
u1hdx+2Gjb7jF3NFkhA7TgdJRQTRckRu/L52O3uLIO439QecOvJuYz+Enqk3BSr4RXBNuyUW0RGa
fd9lCdSNoVQWRBepqaR5t+v5Wp5DzDCbqSsyrtnfWsnvSyPiko/26zEUOKPdqA8Yp0mRpT1lqQTj
wGSUKvmu6oMF2otnOtau/2DXlTzsDd5qoMFkQZ5l0sA0IJmlMPaFSj1eGsN6fU2StbURNzki9JyG
AT23oDYMm336oEgjr29rA0M0bPgaaL7KvqSpE5GPvhAIf1eJOymoAj3lnDyHznX3nnjZueyzM2EY
dYulvt86HKBb33E0ejek86+Jr7Rw4XdlU1cTEBAiG68Ot46d9foXXVcBvCD54Qa2JhzsYpIiy65t
4tvnzFUnXdWdz6zs6fXppA/TSLQKmvDsFSaAAHSWhNYQeokoHFvMWd0dpkE18dpQfSOL5InL/4Ea
wmJfhXxR/ZP2/TGGLgYLcjXy3xH4/RqPlXU8vllxpnEzFDumDAlJsANGFgXax6kyS5mRxHpmM9+J
snGDbghNZdPyzk5NUBgVwU/CR3lmeQAz9HGxXdoMOWJ1/yQYIuBYuiYTqjE36oriLwN66/72XXQX
NPzKZ9RZ748xP8vhsKAj+QLajWp2eFcXexWGU8LkZtzz2TCk8ZmC1dLMjyhpGEgY3VEEyuyCc4Wl
/tHso0Y6hYfnskG0VLjvfLK6OSH7dvIF+AzuZi2IC8VNgfsXSRmjaEAhg3oVNPhhoStISv7NPiok
jFpSSqzKS5RsbpxKTyX6B9KKfxGKS0jsk6kYUL/l8bB5/rxEs7MgpUOjALRxpAMvWBuO0wf3WZcN
htMzZ9dR5kR+fpLKVhW7/sw+T8L/pTtOeymJ0Cdw7kh70OlPHfzXhoDb4ZrrTpUueFVsdSbHbsA1
x4fMNOJypQGZX6HjtDyQBzhb5B0fUnxavoIL5bUQCRXBXXTKm+0IUXtTQesij5RuRx4LXtBcELhm
+kATwyGGH4hXoiUyog7xxX7gwpgDeQL/kIFpykTE7Aqpa+Sl+QxaPgSHxmtZi5VJ5WVf34zwy0E5
OcibwLCWIQLOBVa5xKiaj0kA4MrcXBwkmKuNf62j1WtS+VX7BGtlyCC+mHJE+SOxV/NCajhurWtN
1J5I9LKQIcRB/Y+5pineJNYMcXPyk5suL08+o3DwEYYkifezyVS2RwHo4PIvFfzUBHmqgw3GGNKy
spDRiNNE+MwImWsTEqHVoFqkKB+74tcNj7HJzBjoJwfAbIJC//KfAxTb2OXPZKee/SNaJUfjcFh0
Kw7WpctK0sFrTIi25l0JdqymDZSWntlmhyxCztK/wU1kP9XpmJTkTqhXEMoquc4ah0grnWBdcKM9
Ws0d66MUx4KMSbwa1hrKLLTnis7SBwihe1Dw3QOHhfHDPYrY8RImXqAXcdIYY37SvlaeuAYOQmvD
bHRaJhtJxzkey10c/nsxMHUM/hD+N/t8e3aKOTsB5T+KbJ/DpuLEzqFCklf+oMFLPoEg2XnikTNk
3bUPhi4AWey6WnAbQKhewtAUy4idq97C6X6+8oDXikhY8PA83gevyg9qCxIDf0+UcBY16E2NgAHy
VJl7fgxJIHb3WA4W3zWw+kcavt/R7DI6xG2w6hva44gqI5N18Uui+57fAtUnmXlBEzfs7mSCfdCC
7tbNFSeF6N2nr+SudTBzbFlj6KVi/aM6p3jc1te9WXncvgnbKrZmTBfc7D2U8lYW0RJO09x5upCR
pRT9+weNEgs7H7Ipwcu9AP8FYGhMOlp6EKl28bmoLCP2MO7B56g16zNxJza7NhyZAzVM3As8GYuE
j8HoVQh0oDW2qSOtK9m+cbryiS39LmyUGFEEemX5/7kCliHOyNoDqYNNB4/yP1uSGoqv0BGM8JVV
xZoloBZ6SIM6fDNBuPQFUUXZyK6MpPwNqBrsu/sEGrfWC5tNQ2XlR0sBI3Xdi7YEmGepsafUEuZn
UE2ziH4e4r4SQxFk3Q87Q5CZCzKSTdlFpyn1+S+T2P8NyG1z7naLcWtSs5OI++EfVnGGaaYGlkoV
XbvT+yjZgiDgWIbGMgUJg5w3k39IrISo7sR4+Bon5y6fDVyV7SH1SLNbJSCy54hWu3X52lGX6bTj
HjUtbuvtkytuGkiq8D1jaaMMkYn0h8Tfqx71FKJMacixmVSDPt8RaIFgcbZL/4G21OWLnB2ySpxI
Pc0zuJM+efYmSQGenn5+XinRp1+z5yI709wG0xNBic0+OWRm+cgpcmp/smY6tkS/vRNLncoK5JQY
cloWQ/AQGcOFfcTm5HJmNyU/9jaE5NjzA/ZCer+HT7mMw3SSW8uh/UyHQ+qGWEEkb3aJZdiOGSj3
LVVPE2vUvHbB5vFcrCHrvslgajE9DlwNfWVMoarl8pWa8DiO8+Kuk+OBXSEz+W4Kq/MrX0AhRvRg
Bk37FyPzNZVp/X9Cwe9WWJWrkNHwSdG//+eTn354KWgasFU4C0XKaBO1+smrtG/Y0980uTwiEENX
uNnAbMotLIKAllm77fBAU43WV99p17/id50FI++U9KDgMXrJVomr4kBMeNV38zP8U3hHnbfZ2mar
gnMDuoq63obeYP/y2IkWYTJ9W9hFT9UkfqOIDiN7V6L81DakX0YxGvox+CMxI89AutABqmV1Jmac
XjzYq6ERx+6ItEfWtpl2AVcAXvMeSbmfDBi50Ic08P9riuiKFwxxYoPBpspxI7zfSHhtvVgEnvEC
89bSq7BDTVqyWLtwTm6DJC0PfjfiMwpKjhJO95A3oBlBYUkvrAC4EtLpimgWpWTDckUub8XUPnfk
IDbot6X6f91NoYB1wSa2fTKiVTwWyvvbvF1My0WDUlaTYCbne/NgNIMcfuP0jprvgILATOD2ewyJ
9bimaSd4dnZ2EPHY50dYFjr64N1umtqrLeNxSgxYl9dvr23zT1I7BuwU9uaHjfekW3LF/66Izxh1
H4MZlTi+1pp9aBNk9/nKmzvqDA6X4M5gZzCZ19jxwo7CSgl2ps7fYxROPe//T+BpbelNQpJcGONT
4jMr01vahkkSxdW95J4j6y6/s3su1cOTaTJWSdW5SBSdSpLkooT+HQNbuAEFAVpX+MQsWQHwNHjK
yO/kxDgOGRqxLi91F8seTnoT2Qync1IMGEPNQG/otH2PcMYGqyLdGKJ5s4G0tYTy5Hkg/roxUZE1
N0tuFhcLXxJ0WG3rN6j0m1gUeihrMTUypMnluYNRUlOWXHE/yQu68BuIu33LNkvT1rhsul6ee8Ek
0Ud1rfIGDLwTGo6unNlwg/m1EbbhUrL7ukyVIhc2czsJlx2Mq/obQkQdsOdO7qnYekmj82Sjv0Yb
JiboWJcXN7gVk6Rq8noc8K5C1IoLdWLnDrHynRPddzBYQnsBamGlyQsEoFaNvhhXE/VDACkp1IPx
Sqg85yM+28JMeLk5nQgLvz/6eMmRdskY4pudA3q4hybe0KaRUnLMxqUUvvwijMNjqNoovBAZonHv
kgBWkrJ2jIOi/SIdACXqdAIUTfs2Scnd7UDrCdRcP0nvmMuoqgXc/UmzOQb5itfxEl0fGQwJ27cf
Yr5OZrfTBtlCubnNAueMYF5KQBn74ImBk/hvE/MfyVts5CB+v3W9KNV3ECZR6J5r8FmyYJqPjigF
G1JU+aDcTyigIa7Dg1BxxtZ4uZs5tGaD1SuVJx9NX/mBDA7Ds0UxXIqZgoacGy5UvnkFGtuG91nC
AQANHkAl4kAD2QweYbjgGvBHV+rogTcHW7IW+fatJ9Ay9EN7PYsX03Zw2c5zis239evOHUwlDiLy
UvBLpIBkkfujYaGKPueeqyvug7fH3cKxw/fwF9ZH+SADf6nV0IJwDNHAD9W0R+ivlysWZD0kYgp2
+Y3+maSMHJkgJJFoGQEDNmgWaRqEfpKtJQtTXhUxPkpwkqQr0mogm4E624D2lnBtw1yhfbJZVqfQ
lxtALE9vMEHDsEDsPMM50zk0UW/EnomO2J4HFZy9F9nm19apHnvjDgEX+/hh6VcHsYNvkKY/TA9b
YWVQK0wTg5L7PSYfp39d/ullGlHtyRJCUIUwMFaxqQwbm/3MNW0D80AxKzZvN1WjHHs+a37sZV92
NQAEu+g/e8Nrys9U9K9TrlZ/sQUCH+rML5tbLKsce2Lxq3cGsUonqXYd8ABss9a8ZzZ/FqkREwwv
YNSkVUpm0/KLhUaB+M03zj2YMccbesgAwueanr/u9oMhCpCxpNrkcIy5cFV30xaTrp1+/YWgzlVX
2sK7TJvlwRfNlBMFgMpEQJhEBfIXkgZO2JTMjB5LmWj3/EEltNAFs8FN4ED4YwdorjS5wRldlokL
D9EP7XP/eIXWvo3vrzqZAKXK6sRXv6whnHdUsIxuQcRmKXs44gBrNBe/d+J/AYRjE9LVU1nQL8V2
gvBoJm5YLqIyaZme3Q5/G7cRf4YjWdLSloZzLhaceshmptXyds2A4YhotZPHJAl2ik3TC4258pW6
/hp8T/Sw5wFT3fmyhPP6q1NcVQU8xPqc5wbCson49L4cYCkUPyk1/n8sf1OVzu+BFM86eHHH05Lq
H8NB0GesehzOdbQOxOxAjWlPjH2eSllS/duDn1Yw3MWWlKQ7WGyk+f9md3mhYtVib33irr0he7Xc
RCq+/hO6foy5RQ1jqAgblOaQI8aHdNCu0mPWFmAbWWR13RATmjhGktE0ucnHWLC0djuyZzBG5oij
Q5+ABydLcWmof8fB2k1db6iDgX52IcD9kBLyOYtOWHNSGL6a8XFAfZIy+bPFXs5+AVB9MtZACosr
STs0Dp3TWY/oyboTCeov5nJgyxEfdpZghb5yav6pm4zLenpBlyie5rkPg8XwUuuXhznj+66Fa9BQ
8mrVBrO8QpfxQ+Nh3QXqKo4A1MpemIT7JDsZ80tnFIzmVlCueh3S4q0ceSKaxUgKUvsXkSKKDRBk
ilnQ6h1/GH5mVrEhAf5Glg7wluqe+JBsC+Gcv3Rr//1pWFRUKdyDYr/vw7yxrvOAn7XE7lvWcntn
wxMfN4loLnA7zX7TypylF3MzsoaFcgasrFR9yqt33LLELbk2TlOcigyxEFVWm5k2nNmyactLwIwH
tftGt5BtuVzOxdvFgaqUCGyw93YGICwvTLlg148EbOeShRoWqtBVpxlZ5ou3HZs3Joo+5nSExNnJ
btxpxilFTUxR2rNE26gVtUVadGLTfMJzAcxyAsK+E1AVU91IHTwCb88J3ZJjQs083lPcgoC4mcAl
DtwCkKnZb7C6iy80Uy4pJ2FTiW/CWm8ezc/gXrG1SUvWpf3GttNB82qIufK1ArrlXOGetn8AEHOu
wJHGRRyBhCsmGdFWzTHtOiBRSqHwaD3BVc7Dzemvium2gQGb8IR4F3wBvWCxV/xsXPG88X+vq/e6
3+EJTKj3/gshlrCxDw8mMAMMYlmcV4tLfMzsSIV3Fm+M73hhAFfJ6ij8BVbzk9+i1bjImsJ/a8tu
FnkV9Ms6yxmzFYeQmCMJ3A/d9J/XZ+3Bw1/oNlud23y0cYtuakbz1pZFpXM7sa9ztkOOiStsaTyu
vjI1hslIRsyHltf6/hyXG4MrFow93+RvXorDR9Mwg70DNFJKieAYxYA8XRedcUD2fTTMImgJtiGQ
7bUeUkMu91paYEi0Ftf+6lPNLUtc5PD61GW14/PgovH9Cu77874TYXMtmrdxgC4RszwGm+Xw3vcF
EooEZU4DAXVSSJAvR5vRd3aE8Ca8SxPaGP0M2qy9R4/9JkaPAPCwv9nEBKj5w8RDN1DE7v3+lvSN
a63ZhWqOuAanRSm7UgzYwkRcNHPNr/gIfBbAMKLVfxY9q7ipNI7VXUwJSwrsE1+JCVT59pq4FCoz
/XIlNc94rVVVoCQPvvSBl+3XcqB7vOPxSmINfhicyBU1Jm0XNe/KKaaYJkOl3968SBFelG+KR4QE
jpAED04W1tVy07iALPtTmCYA5L+SIbRmdKFUu/jVemyoU9+SYwewu2JoDGE1n4gtCTCX8Ab4piJl
06+SKGE5KPsABcpOoSvLSU2dzSKPu3ONzynbAvt0JjwfZgMjCSvUOFb2UkbW7YmU+g/C8u+gjQkh
hDy13oOTisA/n/V4uOZxe7KpGi7zpPA/PMhI9Mg/lhqI2OHwJwCvCXaUSSDVLWmqX4SrKUt40m5a
6LRNQvkElCQJYOH7yQA9HEv2ztOrzDw0/dZrAUAt3HX0BizSVDUVRKw3Pn6VH49tA0JaUJuJPXRD
i5HQDytH0DKEr5YuIQ9rFUUiz75yinAsg7wB4tQIK78JPkZ/kkKTOiVwn6KdtHN+kn/V0cYxRfz5
OJ9upGj7eW/7fpA8LBmW2KmqXvtH6X8MC9npx0iul7+FBbHpMNf1muTUkx2Lsymuk7BsnhLYCsA3
daLmb0fmQ5AiNwxIQV0xYnceRG4fEcH02IDWoviR/hngu1PyPpF2Jx1vFll1J9BYrTRxijM2WWBj
Cjq6BUjR6Zq+z8ZGeJrNE6Imqc9XcihQpl83ffR/xiIzsMOs17a7tXV3crjYGxXCm8HUiaMfA4BO
46/y1dAoilyUzmjEfnnLeV9NrnwAYbi5OuljZMtBTpkDmCdL20Mr3355oLgXd/8CvQuEuYsBorCq
Wj8y2P0/cVD+uO6XscMf23EZx3HJ9XhHUl4kjnenS4VtJXSP57yKQV32gX62DgkBpHc8vfOxkaAY
8CzLsTbu7ZqRwFeXO3dvYrUDGBnog1D6VzG6Ra2yd91R230QFX+uJXfDyGeMn/9WWw4d3s+/jEFk
Gex9n/qwO74Db/7aoh0tti4o9TXRcSzO08oX39SEV49NjaZ4U07jnK73KK7k4p3ByrRXLa8/6Bwu
xpjaaAlnRavjFSeDSVujNeJiZhc+1ij4gbD9It72B4BcwKsMl98uv+jT5qdDTBPgp/YdF9fkQRYJ
c/jBb84z39gSPDhMXYRhJte8tLBl8SBoopYhTfgJIiF9Jtzq/vw+Z3xkIGgXXxQkyMOOYYG7HTGF
uBwO6D/xnVoJl02Ma3vvENWGdMSvSPCGlxV7e6l1McTUW8ETMHvFwHnGyFeV01yyHSwngaSE9+NU
eVEnzMhhSk8N+nopc+Oc+/3L4W6yrPXmpYZF4oPl250rZOjp1XKkXzV5heqRzY08alnYqozlKKnI
WsvEsPR8gcrSsvmFbM57mOmvAYA2ZmYTkxSM00NE6mEM1BgejY4RLZky60uT9vAALQneEhXmObWr
NkYWv1uh4P3Us4RSVUC3SE5ae1NOBg/yVvduXcGIlH0XTn6O+nPif/eS1MzPN7YdhczlGeDPAgT9
ejdvvDIukVTXTwpw9KhMw9EutemhzAUuJ+iV2a8hUH4S1eUIMXLLN5gqEw4YWvBci15YXc+jijc9
6V4Yul/yNhBPe4NDcU69wR7yccq7A2Jl9F3TJyrat5zQYhbmdL6kuUNABg9/mv1Yw/QXOwgOwXbj
Z8tKBOgi6lsmthrmqVjkmVAgWesso7AfDxPk+zBGo+TN6akMiRI8u3YykjCvMCOQMWxw+SRYrwt/
DLxvgyOVc0IN+Uza0zy0vYfV8v6BLhAa4pr5SQWY9gG/RpvKg64mPr0xM0bCX2XtzhB8S3hKfzfU
kaaHFhS7WHSAWz5FTAwStr2IArp3IkBXAFliYFeS75vjBY5QjDLGIXd9/xm8s3wy9j1ZD+ysKYap
TxPPyX/r8yY+25Ze+6pMqYjelf717gtc3OK3b0Cy1hdtFH2YKsffHEvTXmhUExojNmNQDe92KgqH
D4lOAv0oEKf0FLtAXGah6ZHt7GJ20Z1IlnjxoJN8BE+1grD/5VL7pXo+UejYEqUH8kpfT5hJ4qnd
JihMJOgAmTTjUPHM7Poc7dLvuV3hUS5bHj2zOssFngtCZc26GPXBf63SNELEErVrpqVy/djAks0L
t7V0E39nXFSJ/8EEyKgUsRlTCSkPfj7XeSz6dH/lw1BeGnc3NvloZvlXMPz6lu6j1WzwpAXYZkn0
wWxYnIQnQ3zIzQjAqp85UrcKjhj7DBIQXnjvI8bjfwc5+ys4bHtw369Cb90wKxATTKWFq2OCxnaV
k/eJ0fwjslBpaaP4XHRCXLGk4GYCNItGJAVlZ5wX6cybt7Hv9+EEB8ByMrEUSFn97zkERolPZ+Oo
1cWE2CDadrotAusQ84R2xa3E0N1omIOlsdtgCl9AUjdtxmbZ3kbiogc6nPO/C0bWmMqBwYVOhDmJ
Ir21I3+w6Q6MNMt1tPSKY974Mn5Db94obzAabd92Tbz2E6EEx4KWbwbq/xWs3sWD8gQGBgo977+n
96fAm1feoaG4esZ01MpYLYUeNh4cDtnpBQUQTZIzXKqalLrq9Fnk8lnL+X42nua/YyIY3ISRajYf
alyvvPnJauCukORTFR/9ZA/yH2VuEaBhFy7sBBanGvSL6ONq3JPOsUq+Nbxe9VyOyBFg/GfFyBwR
VysVa1W02+b8x3iQCTew10wfL0obOvYLg8WVTXuNUs5rTE36T6OJQYMdfTu4TuVxWF3Ul3wd6N+4
dCzZPKD+kifnE3zqtodJRgErBzAywdO72KUwgfb+jsAm+sCSpZIhsW9lb74bYO8evwC7CaP+GAL7
sr1qc5J7w53jcgKMWgONn88sFLRT+yyqyj1K3iy3cLx7rEpsjinjvycgkf2rO1ytEDzWqUfVkx5y
B2tnR2hpzh5B5HqIAt56EPJD4xeRraobDhL8jzScPxc8xTLrpxUPr3rT8VKnZ92P8q4gr1INxMgB
nErwpB07jjr/OfDCqH2BtFPBfvOjt3AJD8YWFjDfSo8L2cWCcMmIOqfI4Isx3NtB9M0Qoy1/03Pd
3GnPa15QaFTSIV0fMgXhLxdZd/p39k8PeMQXsuzBZuYLNomwvA4zxWFj8KBtWkdh+hvN7Smu9y0u
anBoSVUZeyIcqJrsoZSCW3D0LIENCue6R/yx1mL790w+vl416ty8zo2/9ICsR5O5IK6f8gOVPR7f
/UwLnoyDJ2Cc2iHs+4NnC2ZJz1OjrjgYDk/fbWt0+CgedMfiqEzILDNg+h58/8nLaiLS9UJtKuU0
RZkJRTX8byLTzjx1HQGb8jDH+KU6d8lNhfI5NNlxDZcv5juGatQt1fqCvQZfX0xzN9Mzsv4pSbRm
O0PEItZmPZUtbsloVIy6t2rvD4ExJdAvqBA1hkaI8JTSdysUac1FbRj1YyQemW0M8zhR9rWdE4eR
O5LZ+qg/YVQWIF98HsoLARS+qrnD2G4FXr4ZAWgLn0I2WGrwJVYWxIn9gIiZdDzlUpcg74SId7OF
V0u7BZ/R/efjuKaNEpxlZnJRTjPD7I6i4CbtladTL+bN03xEVdC5iat94/A7PW9my+B4g5toM390
giNui2N1W7pZV4kxOmceNLIbIzYlETLKXTnSttcWE9V9it8iV4HPIUUPhFcxbDfWWlAxr1yd4fuj
WrkpiEB0y9mWHnJ25Y3GAJob1WenJGQM3Jw7TNAGyJEsrplBUmc7w+JtAVH7DtRLaCKyUOsr4edD
Jn31KX673QnAlstqDFMpll9fHS2kiSl+8f6/KBEqGi7TqItEePs4jCHXU/1QGySOfyf6Wb39D9IS
7Hfc5M/tBF1noFU0a7ftZTMmCqqAsjGoxGrC5CYXbfDsYdkdBVOH1UXkCORtQYtbZ2D3WTD4YLOt
HAz5vd2AVFYDNaS29cYEiGZSzbYHspUerqo0Vfjz9xHIsuqovPrt5Rder48NazYMd4YtWutYBvWf
q7ET9Jjujx4ceUCvtPw2/g5N/cuiY+1/OVr7E/EtvVj7op1RkOVo2jfjBBPkybV9Uftf27r/UIg5
clT5bGZ4vePRjO0Z/XIzkbLEmxDBeJWfQcEDNXmmXtZcGlNU6AKHfUHxlsY8CffmYdR8r6gSrkvc
2zY04yo+U3rRm3UFPBrXnsHk3923HbiAq3DHpZh8Cb6nHZZKDsXXDPVQrJwIlFHC/5TPIHYau1uu
TShrYk8pCohPCjhfKsRgjqvTystd6oydpBjyMQiP48WYFXkGO4YwsDyDXOczDjku8oaVWPueuLJH
WbHFf6IfLh59L1bNXdRYn88GjmVEYdyVnPSQk8PJ4XqVsmVtKMjrwe6Q74Yt0YiGvhWiwIQi9ymz
YYy9GIcZ0WmdpPT7JPcYqqLcpWbAtB5eZiTiwTbdOb2abGuUx5f/VlhX4uqaIzXo/n+wkiU+ZtQS
gbEH2/YAM53bVO/Gd4afMX4qp7Q224mygambHzRhdZ8jGGD1LyYTK8JxuACv1dzKKYPSc0se1cRP
fxSMEHLEYlRJIv7SfYye1/qFxpn/7rqVLxm1ZzNfHdSTLiNHKJTXKtfxjXZaLT5hslX3XGGzgqhR
d7VUKt0vj05ds1bY5uG6p9+vMcMRhl47Ca9xTvGbjf/jOOWIrrFvL6ZEikae2GAKJ6JGbVgYkksK
XOCoBjUk1ppvlqJ+a4m64/KrbEoFNIoIquzmdXCZeZPspfqJ0t/jZdy5jYRTeG3guQ5JxY8lxUI3
eK5erTNeD2c7GxvzEXldTNo6J7z1RD3N/bUbNB8ah6l7LeuEs3xCuKbaQVGj0EcPBDQWEgFhq0UP
b/7G0JMQyN0B2c0qkPQjJDVnw+w3J89qI4t8lSnXVADs7om3o6950nQLiWhNb1hdUM3futOCIFAY
KT7584euRSGhpWXKAZWKJ7pE5+THXjiuyN/yHtDVFrdUML4sAMEkh/MyjKQ7+6yPv9RW6lJ1XS8M
cONWocai2eksgNCX4F102r2sQpLx/qX/OTGhtGKXCSXf7QLi5szShWpv/GbCUNzI7lK2YrumKH2f
jFV4oBUuW+xjRlVoyfNrFMXcVZnKJ0I1O9KdLj/8ZzayDjGrj0udK3ohNO4s8bP/ICKgjgM1fpoH
5ehxPOd/Xzbi8F+s2ESf0DuLyKvJOXu1GturKA7pl5p5tEnUNuCGPyrDPDNwRVavigglUF63xJpC
nxnfTl8Eu0R2PsRJA3UU9QLH4fUwAyhVfS4Enm1TPh1rbV1frB/IES/4G4bGsY+7Uzhir8ZU/tdb
twXIE/aJmpOsNjBZzXxpXUiqrtAtVRkrW9vI66O+TC+YCYwTr9x21Kj8O197hc1qgKRqrD5C4zp4
kjCkNTTgoBDQyWE0497+l9B1ko+xhUlFGlZl+786U0OU3TyKUhRU+doQMgRP6yxulkLJaqMFH77d
SSJNOywfXKJJCo+FRMCZWiFZCYySz/DRO4Oh0s02PxYD2IHidIXh+pC9YpGrxHMgLFdqFYDxiCEN
0MeuHIy3FQ2e2Q19AAkeYcs//3SOePswx6WLhq0jr6oNzqJ4Lyg/5/bWTBrVeAquX+3gRNIuY7SI
82Ue2fz9MrHg0+5TYj2LRGNkW6VAawuyzzIrt95bd3XfrtSpV89533laXSyQBlrd309urf90CRTq
sm9suKJzJgpEsXwtdnv81JGZlR8aQKr4F+ADbgBq5DIYm9Od/nkpc3+yzkzIInt9FIsmkG5+cM00
GoVGxXZE3Qo8/opGdUCd7Z5bvhRpmjW4MA/yyoIgoZUKcGuxVwtg4Fp3zDfoIuL08LMAjeT2QAJY
Y8g/xBPaWkMcHwjm2BgXnJgpKvepYbFoBphi5jZJ23M6dlHpojsw1K7KkR7awGLfPzI2xdnHP5mf
neCnPEfuYP2edAi/WBvASwgsxfp5hS5BcBoxlw7IseUP80qhn4mKsUnm03dsw1bPaQhFFSZWU7ll
fbRkbIioCDkMABQPHkJGReXbFfw59kH3k1v7fwQ2u87DI6pCCptL+5isVZ6w7zmhcpVoTI0h6P3u
QXxOANqSrMQLc4wASpV333jDWrAjQwZ/zwllYpmMNEAAqvId1BRDwmrpF/ScaaQ2WlHiDUKOXQQs
tXxSrb2aU8Ktn7bOnpNFF3xvOcRIjyYQKAjDh+8K2hKCw7ydanQ+uXKvzFXI51F3SuhkHKBzZp2r
6EBjv3qBtouRvHdSOBpg2WvgojZX3bUx0Dj+bJJiwoPX1CqRy9+Fdv9g+Ej45Lfd6KH5OLhIOjK9
Vhyu7mbMwX4Q33AJr1mwVZsvIgxc3fxqH4+SYAWSWSSfCp/Agi13kehhcWFt3kiEfbX9V0bHxbke
zn+SuSzFUZip1sxeobfHGeBGXy65q/9a8DqDyok+DGDG1PnF7O3VBfkyiTtQMhfSwyLMqJwH9V2m
Mh7FOp6hkLvKnQyCTbJJm0dKrmjqTuJsbfgU0ntjoZldSQmPiyhGjauZqCPBTh+MWO9lCsumH2E9
YwSZzbqSxQuaIVWtR2oTQVmA56YKRaYdgsMSp/kg/ntC5U76jS8ZtAsGQ2HYfUhnXpHH3YWWD2BA
j8uLTvYhz7b5uX/oZG/JUP/X5cq2/vW/oSirvL51sT1rv4D0gMYGgoflJ0kOLMGxEVgHJH4swfa1
B2ZUsVL/frn39lqY0X1EQF0QUQGBbtKTZzQD9+XkNHVbW+kEmVMRbEm4Nyq6ZAGflS4Jkwb1uEQ2
0WVdH410tYu50wzUA4/dpCtQiWJATNpkqyXx0E8FHzcskvkTThRMCYUhGgAhVL1aQ9mfDYu9KUCC
6nH8x23GRzm9GOeI4XQBRPa3GWW/fvYKNKpEn7k1LVdkGqDjt126aIQ3urJkHgc276lIQPYOqRi6
6uY/6JMcDmIEEJuQTlGI9x0YNaTfgMDQ7DACKQJ86kywKGdclCXzGr3qIZB8ZitZ+Lh39qwc16X3
3PvVLM+qdCRQpdtwuuCSkZzEnwTD41ZYs5+E98g2EIq10FbAi5dWe+JY1tdgvo3VpIds13Ntq6wm
bESktXTtfSTgaUVrHJ9qEW3MOM3P15g0FvmGrFpkOJM58t7xmixwupjd1KmYm+/RxpqUbwC3EmWA
dBDaRpdKZtwGqPgWlN2PbIgcKn8mPGfKe63aYtMpK4jStNU8L59KivgQ4t8eptmw282MlO2loVJN
84kAUWv+Va+U0IVm32QNFk4xgwlcQbg2MmEQzJoDwx1wV+AWXdBqk9b9K1sTrag+BCLxpAHHScwe
dCNwXVxSx+pG0JHJcbYIBrXOuZ2a5Y4Cq1as1wEyHWimQXlD/TCuI7G6cmNQoEzKAmsT4hAMpCp7
jUMVbI2dprqjHsJd3ScdKUNYEmx9v5NQQh5wB9pv27axBZOnYu219hVs8D+XE76UvgLLEHcYNXBO
+ZUoCPJrd8TGgXn88WETb09y7VJnQLe/lnJh+LEEJjP8pMyTmjfW0qlIuaWx133i9oQmAWc7UKKA
it/EihQXix/UDumu0JJs9qQyqY/NDjV4YtFrAMSfmhYEQJA4vfSuSMWLRYyWRyZCH5fYdeZKD9mp
XhmbqDe+0yZhwrFTnd28GewR6u7YhWcDloN0b5ELwq/plTIJsCNTgs1IZ57BgD2Qf99jiCqVHCNZ
CNxtiMYguIv+lDtKD1464sMsSYrvPiazl/vugzgRS149BAGet4xBivdvmOTsH0hZUgfHXMEY53fm
F7/9cUcGtJixPv5Q9UnECwK8GGa2DQd29tqZ7jhimm4YyT8jePwfCgTMuACWe2EbD706zXVn9R5B
OjApD322LJrO3jFBXz0GvxLSn7/THP2kEgKMvjQ02kcKI6SKAORR24YmIkwgxotmg7dBaMo1kvXs
M2Jjz1Ua/+m0KvkzmPDfIDpilKoxkebE8g4vnFDHmEVDKIIP7Fp5XPt79h/ZVTXP7uKwlGG7+MsK
HBj2c/6RzfkZ3YFII4/I5U05D0XTAY6UWrp9pv9MyGbI1Ur4tbPF479b1wG19UybnhFcd8wt3yJz
GcpDVU6+SIQfRSX6b0he9WEtMF3Z0aDpGfJV71RT8+oKeTBe0DB8qu4XaWWN5oSqfBj5Dj98E+K5
N1110LRqvfoM77Y28TPTZgbRNEYX8G/UPwWaPXAEvHMCPh+PwYnz26Z9Iq9OVpbjFLNAyIFlnIJ9
F685qCHC8qT55Ay5KNNWvGUlGIrMB/2emWYZTTPNBZKv0QdByQ2Uy3elKNt4RJ4BsHcBAqzsV/2k
Ko+JLgGPa7pLpE3sdLPGRIDmDJc/eo4lRw/3ZOqrvcE6TSGmQpbK6IGghiGQvZcsdMpwi3ITPwZZ
bDkaguTawkxbyyBUD9jtTfRU5lWHvzSCP5+KlacuKuFyrbi1RVixhsh/lqhC+bXJ5HZFNSKVE2Jq
mzQ4fI1G6lr/lNQ/Ab1hNcWFVrFOtNvSFRrwe+zbjloh6ZdFqHF3zszzCxPxHx6HhtjZ0vfO/MY2
0t78C4UxfsQAbap9Z3GhJfLlDSiZAC/fPqYtyAI4qIWbIe1d87BWjD8tOUFVwxRsvCxFOC7xngqD
Q9UJX4BuEW3o+76GiZQSlRZP+VjyXjF6QnEq2wqmd4ADDEMyiTLhdCCQwTo5pbWbxJdB/Pq+OJE9
FUK59jBfufX2Sn6o3sajPkPvoPJtwHqZ2QJl86MhEF76V6MTq4I7JkeoTDPTfAEvWu9suRb50/jN
VcK4PR9jba6yn36/XOjI+wih+8bW2rKX+nx58+2dWQB4OQ39PWMvbH8elq6wUkwcXN2esShPjXb5
VH+AhRYE5+Y1WsNKGLD4d1Ne5k7WTZDCBjFtKUdlhxgzWA3bOAx+jX0OsIbrHeLtjghknH2MCCMB
2QbVK2VanfHPywOY/zpDXMfhSGfsbxHAb7NAxQhKAHLUHjFXkr/WMS7Dt7r/OZT6h6ZwncIUc7NQ
PeHA/fr8moTdv6TXqhOyyvaULFp69qEjeiAxHnzwqHRKKCqe63VKz9OZdu13wvXuZdxwXKMpVN6M
Vlkp05vEbuZhu6gbfRLkd589YqkzyLEJhgMJ7rONNCqIexY5MjK1HnNiZ3Fwx2SOmIKhy2DnYPEp
Uu7ZtVAY+/nsBstVRZisIKRu1bARZeJaahIUzeH1vRG8k5+VwM9Um8no9DH0ueOG3oEyO32SRX3E
5t/kQsndwcIbpJoFYIzueiVNvadQ5vOgPeiWEbr/b3zAQbIIUYCoNbm2diSSgYqNKbeRks1L6rs+
+IQfiwfd9uQS3O8ke1b9N5c3nXI3zKEAYyMHP2eNJfOc2YLb9IRvPfE2rhRwP/ocds9u7j+dqcUz
beuzkHnEuqYIQoKm3KXSXj+NPShoSLCSvnTRTnsJRIKwm6KL+exkW5wtqGTJ2PqhRz855CqQMzAJ
S58Yh6IGKUI1WpIAFX9l3SprXQGYH7srQZkr4d97Pzvs57q2hNg+3S3WP0ySs841CbbVh8QHaA5b
20l6QnRhtCQRK1vKCF6Wc5Cu0Jcg1enR7aueT7tGmfllMqG3RwlwOLDAoMor7btggn5/UZCeaaLZ
tOyVsqhc/QHyZw/wv99fv9l5dxirFi8vOnXF7iOqAd0dIE+3xtJjX7jfsaRe8BOgu1fvfnPY1xvU
+/Enpm+EvHQEFdN2cUJLopofbFAuLKCuH3mcIldVtF8Twq8Af67danhakTIm5N54OwlnGeOyy7mf
pSmZ0hdJphdWRd7pgu6nC1EM+0Kn5PVCjl+n4MFsFGuWmo67ah5D7olPWoQ3TdOigqqMWOgQhPGH
VxTzzg2zq3EDzFfI/ucEM/ktjy9f7bENJqVASjvLGbHD0A72GpBRCFoNDyecxMnuc6jsf6XY/6ut
O76TW+gBO2YQKsdJLh2UYB5dP4oA8tJj81PjmjEgINvpGUy1CNThWq4VbyynL1NKql1C/Q3zzeGb
kbXN54CAktZxvaJtuPn38Jpahv4/8/8rriK9eL9Ym7M8UOgyEREn2HaZ/nyiyXACb6IF4WCUz3IO
nivRbDidosGiKFW9wmHmUbd27fZ3akJt7szhu7OM9VtX4spxB89w2RRfWsvMKkgRY/6ffcW6ryb/
dwV83XkSvXYG1xyiBCgdFYPVgJxRz25H4IU9dvTO/vvysdkzjj8ubZR/kl74fdkxbwMoGlE1iM2A
YfaxU7C2FZ5oWsOTGVod6WRX0jF0F9yxsNpfd6bdFzz3o6/znvKlpgm0jSyJrFNYnjVgzIptTsuK
KQ7aFITGVOhauppkF864GVAyO+E7xKUPcp2uHdA3SDBRW/714TdJ4KYsG8kxF988mW0f2kcR1Dmb
pJB6lmfgFk8aVRBY+4nNmNohgz11JuwKhOdLfhWONXqtN6pcRU3Aq3AFdUO1noeW6WwMr/oiuipu
DyL7GcyQxnhPne35scbTJ/l+J5nNyAq1ZH1sW6hfdSdIWf6yWTr9tayOuPntxFjyl2wdvUVZdvni
rPNInrUH6RJQ9AqzoMYJQnizqKOSATf39toKy+UXgo2qbHQrFMuGYPditAQzram+QrMxUBRiAd7a
QPPhhteBDMmxnejw7dTdcZVIDhV0DRd63xd4XYq4OK+ALnHAU1XW7jdVKqhwlvsgj63UMcd0Bnxe
CfNoxjq9DMecTZhYUepZoe4n+XqmKg+w5e5cyn0LwK/ZYW73G3GBb9WxaOxYfhJGN7s8B5xiXDQb
1OBFZL434tqIKEGgl1NQoB9LoPaSk6G2//SgKP0+ztV7DwpG2oAn3n3g6IyMV67KQYmviVm3EHeQ
1Lv+IK5EdhOHeeBBCKuefTRObP0k+/IAXPRWv5ooF+Sk9UKy4bnEfiWR1PTSO5mP/WoMSiuXetIk
+YQES1+gKJKU1XLklkXBqFevjtW8MIJnHOzWIrTx5sbM1CHowLla1q7YznPg5ieDO5ndUx9Q9D+E
QFknrEauYCaKAgv73pwz0FvLRKZszvYjm6+FxtOvbyNsFJvXeCUzXptlULOqE3iicmHqjjVpd1Dr
Vq1rQrip6Uqx/ZCqjLM0RLIeQcivzYMjsU5ULQfIKaYGXkL2F7aPsMwL1cG87rHBjL2rEWAX2hn4
OuzwgrlfI7wnNiG8F3tdPhHYNgc9fOjPy4pci+DUSasok++XZTA87x8Aay+EOPNjPbO9ZtQcHFph
4mL5IrChIwmTnxfsPkSbTjoq0K4ctLJPybfFz4BQZXT+TY4WDdBeAAbzlyashwg8mpTCqyJ9hg/I
tnDFVr9wqvYlpVDwesXvHpKqZ89mOinhhxr/cTkckpt5XH8qlSfkSE2rTqpLOnQeVwMnJA6bbVi+
ypyJAr2RYSz/mRydf0jEYa9xE0fdBYQeQN8b00rZO34T6Ob1Z+e5J3ypqsrq3zPR601IXA2YUseB
JoZmqaPJ6OpTpodsmZgiNmkjy7lxkNYxwa0IR5uagzWKjX3hXIt4QmkZ+oK+bAdgVhXvG8itUk3l
MrpPPKrh69/hSQVEAwcZfibccS6pkQfJfZrPbA1+u+p0oXTmqGv0aJE0ecAyvDmtv6TqmkqRlXsL
vPTT0/kMI3HVSHbGkcizPWjc7sF2WiMnvEaJTQoBmy2c/HOVclSCOp5tiFVRe/pgyb76iP3puw/C
DYO6C6b1x2NebVocjH0OD6YgQ3AiESm+3nUauRwtn+P09zGoPSwsb77i34jKFismqW+19AQbJJ/y
+RS5w8/5McYViSs27n9Q7SQv7HSuM2rmmRDi4l8CQd8+gfIZaao7PPmXWrGFvj9JCAC3ukkOnIyl
t1vL0vBwUF+JkmXgsvoiKznqhvbFEea8aST+L7JSrd9KPYh+OiwbVNnKfEq51cKNcH0ij/Dx5Wdd
VAW8tB4jkunb+VDVtux2ZRkxowcydu0khRFmMIupm3zc5tT+1glAdCsufuyPHoyvJ0Hw9WZmg9x2
1K2LYnOPaxnyZIgH8wri8KPCijdRJOBq42pkHjRPmd1l12Z7zLnTlYjuf5Y0sp1l0LAggAZ38zki
jiOhDwFCgVQOhS5JRQn+KolTcda31qm98HE6Mhwy0YviLRRYvN4gHjCxYjXDJzX+cftTOqyQ5BSV
0rkEP7EPzAm2SE4rUD9qDvFDoifaiB82Wz6GeJhuhEJDmQHwIsPXGmUPVuWJqD/pKCAjA+sHZRwM
Q6Bz4Kd+HC+VAu4Rcnkc/g8O91r4ONFW5jiikNKzbRtJqaZdDqqfUvzoFMXnG7Q8Zaw7pdgxUsJS
VK4Kg4DikD+TW4/1K/vyRQ/OQ5jgolhTHYo9uZOPmEihrDS4/ht9aG8ZBsoEDhfIUisFSPmXyVOI
b2uIniabe4v/ZwRq66UbHttUwNNeQ7AuOwjgsmQwLJ6FMHkgWS7hZqbsfgyeYqHCRPpsU8mVOYtL
s96GMyZb7mO3wjet7pdTTP2VDCerp2SsrJRVT7+Jvu2BVwSCSj4bjIgW0rIJukjHszzVzNAZlAqA
ZBINLVqOPwm67z33ZYiLL+ZlJpTlQ7OY371UiXQMdOWbgKWhhRzgzfGTGo1rBizqLWWd+FfgIpk8
vhlqJTDuWcZ0h/ogDMM3F+ch/qjAN5lSs7b9g5b8rB2qey5KK4i3NJNWC09X5X92+dBTxmIjYBiU
crWxH3tZWbEp6U5PEr4JKJ5yxooxTVFi09mj8JgdIabHRoyP7aR0ucq8R/yj09Ig1pysn6BPg26N
f6lYck3Hmwvrhf3KZ9XJ3lNhAycHKUxvHcspg+kgDHRm4YnjMqQKzg+ieT9FajXQCJzmQcChwdG3
ImtJ82tNWN3zmSRzAXwKwQAO9d8XsicypbPcOM1zSTRJ2sDBieKp+ME1Ne6bSEeVW3FMnNzdof01
PduYyMH8bWN8fur+W7YJHZ6OG1xOVjVBW1bPRszqD40VEJtG3gukSiWE3nDdwyubg7dZG4PtLjAu
QFkcnlEtdw9cA9ImvpVOvKDQsOzI8k6CezqsGJC2Ef32xnoF5fOpq3Pom4pmnEYI42Ns3Sh+BMYl
vzhpSGk/5G4a86dQyiGcW5LsuAZDsTLq3cZrLK1qI3cV/jOPpNtxR2tMz1EIZO/2219lPpiux4K0
7xtBBnySupLxpnaVWzdBpIZX9H+ljoW0RAziR8uO0fxWUKZoRpoMnBDb0NtjyRr4IsAgJ3O0XbM3
mroohsfdjZ1u2MJgpYOMJdIDawl3MzPUdbmoP2gAGjpmKQ32/m445LlslrROctpQTLnPztVHmztC
OTtaD9V7pBnqF7mHk2AozEHHeFKJIEHj5NfV4oN1k534IoOU+Clvp9JNLJ3nX8HLq4fORbY4zVNa
oiL9K/tlv3IYF59gkVsBZ++0uxdPPycQR6e27MACkkU/YGNRHraC/VljlDno8A7QDikLmr2cBoTt
ObwAowmZufiJh5gOACdjsbZrTRjU3jwmw2Hv912VnwV65bcAEze1ieo0k8RI4ts/GyaYEf44iouS
3k2XL/a6Y5qMWSiwIVlNSPmCIGfn+N9RAuWBaA/bFmun7NOT3eMlEC7cxxUpl+9j48m+vbmdqTkb
x1vdr9RAMGI7pW+lJSso3ForQyYdUR8qgXTHySWY/VgeuRHM3H/rLLVDMbNLrTyGKfgvt7R2dkR6
SpHHxBSI62z9ub+HpK02wktmTAOul4bKDdYg7nCgq38e3ghrbwPaUNaeee7xybiKfw4WOYyuViYZ
aUiQvx7S6nb6Nkem2rzurKbKg9SaYrMAHLfFxPpHfiGTiTL+gKwNH+2PhQIX8+gmUcjg65ePuwxD
t9tg0+5FtOT/flB4fq0ryqZ0i0jCKJYRYRiFJX/Aeh0MpD4x9CDUBTjsUVYa0CoV+Rx98X7MBSgC
64sVLgzlnalgiA25nf2wcWzc+GDm6UWsAbPJSx92MVcuf+NW4ShmkRLgqUxO1tEeGNXNf5x5Ns18
7KfREGL/YpFGtc5Pz/vD4r0rkNms1vrEffqK/qFn0izZkii4AooUhbEJa6pxhry0M9mznVD1V1yR
14bQY8kfjYJz3UDA2OJJtvzXc3bB5e95/GNwW2AQtT/SoMEjzpyTmuyqa3RJ6J+0RCgo3t4IWZT9
A9pfk/8t8bBi61AatZkNoCy20k6QENAYi6FYsN3BPDW14tnCY9MmWsY6KbC/3GpoYy2izRxhS+Px
n+yCHupYr5KbkagCsTamNn4KvI8SP4e6kpOhmT5uqa3fBifLFOn5tLNJp4LpAGYeFpPZJNmIqqHg
ykxpcp0fW7wqIK1c3MA1NohJimTW0cX53mUUjfKz6HTkX/GfeAQpPyN9DIgHf8J8+SElMNxKnE2L
9Eu8eUm3Fw9/F/7PUirChVo399bEFqxpUUGTLZFYCLImPJtNnJL8NqC9cp7wQ97p07oTZnBSGR0w
VKJxiLJnDpeQzn0aq8rr4a04OYEavD3i77oD6nm4dc+ON652YZS4QKRQrH6jNpBoB/KoadtHIJvM
KW8aWuxFaxV2EfyLPBhnRxlb6WWnd+eUufJGwB96oDY5KFFB68j/AoeVQ5oi4lPoXEO55M7r3ciZ
ATt35Q8bgjGr7g1NYUS3Nfc7ziz58YhaDMP99RD4fYgTXAMAxuCIItQ2nsW7EqcgWUVZJ0jvN1yY
nhpbAogrwO6cNUU3/NOnAe60Y/vzmg9IIPT/Rb5xgf9oh10lWXAAIPnuxgJpqQ+XN7WuLo96Zg9Z
BqhetwaYf2CI/FZ5S/Tvi3vZhfVI+muwox+2pm7PcyHccb81kxzxZFuSSvPF4EbJEHsabGnRyQOc
6T+tZbem/3rhGwSRom1TIiAEDzKnvjXLggEJW189iAPVD4OV41TjEa8AEm928CvCxHuTXvVUtrru
FF4kNheQ8OPs/SvlSpP6p+bi0HTLhSHWGWMZo+/9bxY0MbmVEoSsM8OiIFNgLq8QHL8ESDCrq8bb
qvO2CKhRpgiqFOx2P+rV6VCw41G9hnJ8k4mRZ35mxxi33rLkjnzW1gA4K39xGMYxVO1XtROQll0i
YqRXLx5adjZJ1M4fa0TpDKnGUCumpswiC4h64/3uzOYdmWrtUTwYQPQQK0EwZ9aLhjXwP81xw6Ix
cMqZMaK7srHpJJ7DHIKBWMtNIuqkfLaxNShCgvZp6BSievFG8QsRaQq/mgAEWRZa/rEvllpWgoG1
/Sm6bNRQRtW47f/Rfj81Ag7p2/TDNKQ+rOVxxIRguh+dNJyHDgBLebvKeZWh0c3FJSWlmJW9DEGf
eELFw4xBAVF/C9L8QDWgoJ7uEo2TrS5lKdMnAsZ8Xinn1x4w5rjYOkEWE1RP/HcOq8hkx8qitSPp
WwXLlUpsQfs9UprrvGHPl6T20jRO+uGr+EBM2pOc5cQHRzCCdEjlvEXIPZj45NUYPcCM9rHostBP
BnpEvBu81r110zFSkGP40BTkxHJUni/hQzyioSAqPbfs+wLEUaSYmRY9gwP2XOG71nm8wmzUBEX2
3fNvKh/rxZtPWLcT+BQ+tayUavg//JWS8Dg81EAh5dTjdu8KK9/LilNyBURXeXFw19JotHR/NCrw
FzKC/Yg5uvVa3JB1aL1YpijksrakGtXVz4Q0gttGLVu01BhJGOlQSqsUZaZAB4iQnuIGQ7ZQ7HVd
JjJ92YosZQuqhpMx2/LxlN0Gk6xG3DGRPoO/o1n0/0T72Z11mba+7KwNCu3Gg8VfT8Du5YHFE/2P
lReEKj4KW29X2hZ9KPAIBEcGfjIGTNwm0bps9zoIGQNtqmpCwOH64/xU1P8cH9BPujF6mElLDsZ7
nfWbgijM9GWfxfd5qyZzgDkG/dawqPBV5ml0+X19dl2RbB/JeEbr0BIyuzLQW90kp3SbuLMsuMC2
THCx4xCtKzF7qc1tB7cqMbN2AoFX88bo07cuUtIpofBxDmLF9YqDqTxLHAR4xe59mNXVZ4HjVIRz
Kz/eIin9UOTmrhbFbmmIHoZjT73mgYIhs71icSN7py1MnSSN3nhgdGJBRCaO2OoTormo6WiRUkeU
0d6CJ6phKqgFoeTcjZx3V1cJRoDjmp5n2lxZ3SgG5i1HIIXdYqPF/TO18Fo5kFcDT3T+PjawhhHG
Gyjt1aZ+rRNplsipN8q2ro3Fq6MdlNLQbBneMAWcUPwA5vrvyyke6woA1MJYRboAY7Zm0FW5+ml4
T6lnZOV5BRlr3JucuhYljBON3MdbCvzlZpJU0kZvUYH+F5vyJB4Mr7zp/KYHtRuqAAQulZbUD98K
AWTtHQQR5jOQRBB8oulvtnj/01+MEqCD5WW+B75YZ2lBj6vENUJAAUvZO6uvfvsM8Bmh7Z7zCEOd
XMXbWxg7XyVOoKylN0kDZ8q12IV4Gpaq+ytwu7pMq4bs9sX/vlSnx+9G+9nREcyjwwMndf7+Hj1F
P+OKkOZCZqaP2OIXS5WyJx9hUQzDYzHDbMwCuxuefUf+ikvQqa23olk2y8SZyp3l1+olyF1+v1S9
6kDQ4mlQqcREer1Sy0izVbP8cMQ8haVGeVKnLOwRYhn0TJ+HclYeS/ZAZ5lrHXS/ckcS+UbsdOPW
l5U1IvTv8lSEXOh9XaSlWq+TAzt3ajE5lo8Sv+QNhBTRP4UbCIcFituWx/5uEpcX/PSfHrTPh91T
Z3ssf65e/+Gymz7YXVWuX/xxTJvaFFsr0AekM3Zq85vhnjZnvUMYO4x3x7pdN6qfFwmANCFbLkDN
Kj2LV7lLvtkbwUNK9e6XFrBga7wFSkOF0YwljXpduozdTyKfIfMxqR9N4mxy7GXMTcl/DlesP8zT
gkCe/oS1i4NUZaDz6fg8wSnv/HEMW448ptzh5FrrqhvPae1WL3lEyxLk9g0G66B9/yekDcAs/dRl
HP9KDW8tnBc7XUI8rgzP5IdGZ7lT4YKjsC++BIxgV2As7OfLD7v9kT7WKzYbx8vE+fY62gGAY2iJ
XEUPuOtrK5dO1wnl6n1JoRkXxQQLYC0dD78kV5vrJKG6CIsyqMcl18tbYwFudcUcXDG/6/t6gkd2
7x55AqdyJhgOaWsIWx4kQSc2zceEcO+/Y61uSyMqDZYAQlxPm7WFxcew/ws3H2T/leMjgImTpCug
/RVMBbx/PjsyDr1hPr8JhgmEAnlGt3bgfDh9RjHM9nR+G6PSJMfVrZub6zSL+r92aXmT7Ny8Xc7Y
kbACutRLG0TcuKdo6d5JIWNso8l8wOVXcp+7Ai1Ceeih9H+BYGG0LZsvKXSVlMTsYB/bCyj0/VmA
QcYY0wJk7dHVuy6x/+W9/0dakrLz7b/glQvMrh2v7I6ZqKROdKHLPQrcwXEkoiKdlUbV5ZAFt3o5
ueuKGSqkaRojCImDTymvqxG15M9ea0jirjkw7KVtXCg8PogMQ3UmrMTbixcLpPFUmc3weqqgFNjd
OLNubmZIu9fDSW0Cu4+n2nmMB7YkGCNyD6orLKe8ai7qLqLIBFbfcuvK89fPX5ngznZINPCKxdaV
5+4dzpisms1AbMc8J6QrfGAlCxdTbYby5vWZx9NoYU0YK6xXI4FmilYs/MUnKrUJfLHbUQFJCNm+
P8z//nfDCkY6kwPYEKj0ep7cnEoETdig7zunJ1jk4fhNsScT8jxWJmraEGe+IXg47R1niaPfz3gM
B0cVnIAK0aELoBnQrih5cDipjO2MauSCm4TAw8WEIP0h8m5/hlJK3wlINy4PnqTyhulSdccpwvLM
uy9PVaGjBX/xjSsXq5SuG7o0lpKsGxPEbYGE0+k4bRo552aCRVL8Mfx6RkRKbOXw4jIrSMtSZ7b4
yUqVpxZjdUWow+ATu4oPj245S/wlqXslc6KHx5IiZpQSygTjlVCVj0sr5hE3hNNJGoiO79r4OuQ7
ov82WBOmfL/dg0PDpQvynrmQ8ZzwIzefTjU6j2nfJK0gMOUGyj2jcPRcRbmOmC5kEE9XGr7iBn/D
w/LyK4OGsADK2CeF5SR3YKPbi+lCRFE1AV6xkR9ZN3DPbaPW8hcRdvke17wQJ4SXIYPkU5/r/R6Q
CzWNfXINOV2tQgpTDlWHtjTSFRLOgw5txo9F6EKLkZSKEsKDFa53Z1Vvg5Yn98Su6F/j/wXHEbOO
TaElv0tQ/W9Z5IevvadAKj9ngHJRVR/7jXqkaxMoUBb0kvO8VQZlplZZXOGci3DDF7eMf+ZBUMaS
7bD4JZrmiAZA687qr0gfpkaPuUN57yUuiscKK+LdZoALW5nztZFW0rruhSrj59rmGzabd4x4dJQd
genI8gvfHizHgpKYJ78tt1ca0H5EW7sJnHW3sDUaHP6nbHruxLr2eMai9mVe+HSxHNcYn+zVlv8Z
l3NnMb1pfeJgv85oi+zfx+3A/UybrseiPVAPynYLerNuNLxsXURZBGgNwvPijZZ5XW7RedwsmGMi
CLZ/t1zqY4sVS7Jc1ftd2Xstl+7BENNXnfxLxoaLuIJ3Qa4bI2DOl9MbzgqiNzX3vDPsbxJ+UUW+
Zq+hfj43EFKdoktHgo1DLuo9GIwGN9YiQVS4QlKoBqSKXH8TDkFp6Z7jo9PG4WcmOG7Oaz7PRSvU
j7hL7E88NtlzRex/CzllRWCS/8J7cYlFTY/GMfw3gsbjsA90FtmKvepbSa23c/pTSCnLgFU/M4NM
9mkzfStWdN80G6dho1cVGUSh5wKO7sg9NA1B2rpvTeLhaWGnKx+fgVntg0sMwlGctQL1YAUFvNck
qXu09a5ftCSeqh1HWJWA3OUQHEMba7Ymq4DRpkifsJNleQHfMuGxkk2ysMDQW60xe+jEUcCS38FN
iOPn3qIq+Gaa7/tmo3AUMsO1d7La5ES0IUD8YJpQ6qFtcrJPTYZ0OV1MxkuiFkO9lu7NgOkBConb
mMyz4nc+wSNxLcxolhIObG5Y4J6WRkYJ2sGII4SRgxafNXtmgxs7oOGI5JXpza+Suz1MtvWsgXzo
bBxTrr49Rp6xz0DSKGTT71FnG30ht9Na9hIIURhRhVbcMQeJqiklgBmFSN8YEemAdGUp9Os3m/L4
3vDVv5DctqjyMdBk73mg/OApKQ7igYndi8RIfYznqIOParkoE0/Ms4CzleMvBujchE3lyh19FebZ
9ah2RyQHZ8Gx13qYLYHB3XtHtLKW010nufhcZRCaUVfz08mivT6U6a924YW5v2+36elC1TOUOBzl
rW7dBfcDi5ECJv7+jYR1XjeJFh2Jm3FsCrC0k4f9wHqk97gKUj9Gft9tWr+05jzczidHfwyYQeQo
y/OpR2mM9kMO9sLjmttQvACZKGa9XBphhmWpEaTE+ZROFpRaQOA/JlRC9RWHvcZZVgzH0kFixGyB
m8/JjfKyA9o7CzMUhTLX54505bg9689WwivnjCntVIXZQLKZOaN6pL1A0AqFORa4Z3t8jS2xew+t
ZBsAQqS/NLluutTXHIdn0VfwdQooophqhHLExRDTCkaTjYVwGzPvSIfa5x9YtU+KFbGvMLQSqk7y
ATz1SLB2gaHa49Ib1w1xYkan1ZCeBes4LmIALf1nHxW+oesPtxXq5ncB2pgZVkUjp2DUUzSzyX5g
7DuThUepYfFuYH8fveJdgcxS8FwrDAtP1m7V0sDwhCAT3NviD49R4aasmd1v0a5oSWVzvbJo+b24
uYfN6rz3C/SXZgXC8g3AgO31SSoB14QT2g28C/8nLg9YLVb4ZKwWSEh6COZRAuIE2DTWwtkRaJI2
avZmqKffBVTnozvW6CsrL+LkJ+zGIKVxZnXeErZ4LhcDRRE4xmNAq7wB/k9PcAeizc3F+aIXCUtU
aIzTNS1LDGcrMzRzCeXM0dyw83gkx80gvbJdhkK/3rraG5EhED8pGHQ8EkzPeK3lUNco73kimWay
AiKpGJMGYcJVxNpPd+ZzIWI9wLuM3/tW12e2IrzPXdSs4lotv46oqB/mkyGVooTa996dp3HNzHyY
JSNsdiDbmFH806/cqYLBtor8jGYn38s055B3CxX1NWk+c8H3PNmzwt6VAUItBsZYeOJo27pIsHUU
O7SO5ouFzs1CsMW65GXhHd8wpRUmGh2KF9OEG6b5rPPsLYBcGKR7T0VwpoYtyHdvdnfoYXPmHr62
SdvmhV/ZeItYhRMc7zhlO++eYDvrOvEDTEwSIMByh9HvFzBy3R6MOyvQ42oVh7CwmH9RbimZqEZj
5FomRRWGuNgRNkkJYS1RU7/rX9+0qbMBtNaj4d3Y8aOebgFPukAobnU2vBIrJlsUgTEOk2KknhjH
guw1tL1mXi6tAI8OGyhcFmnE19h9iPccPFdSj5JEXibFMQgJ3hckwaeD56YZg/Y40PsqeKgr8C44
88OY6Xrvxr1WgGVj5yJ4xMyoDggcsfF9UkisRHpqZD0ES/IXlobYwMsqoJV8hTQeBd96PX5Kqu/g
SFhn4re+EsJrHMT0+h5sEH844jXg4QIomLvmxgWtOcac2WumApsRYAReZU+WeN509qR+6ibTueeY
jlR+PidDOrf3GEpm722a0pA/gJPHxKyCMtBc0hsWtBsoZtIGivyhpql+nHh3PlUuryF3/cCMSuiE
v4qMlCHzMvdTNwC53n2nvMrNPoNrnF+ZCybO7C7POlghXRL7qzZWtvaJTPcw7flOHHobAa7/9Rqs
7KNCeIwR7WxP0/baBKujdBsmXS0OJh65A4yLsqt7xqa1BKXdoCtli8Z027DnSAMW0BzY8hUjR0KQ
w3rPkdNlT4NnFOrQ0AdiNORt8h85z73sQ4gxMecUfcq7B7N9v7hxaDXA02/dzeXGkLRHlfSC/vg+
tlZG1g34/fKJLhlpo9AqlK7WYHFi6xmiSMXCnsJZv2rlV/iJH/wZbmJMuKsDjM+uzW8XglVhoS6P
XJylqc9Wqv95U/7QVpPWCsycBJtEvXAP77vxvR25W2hfM6AROElOWGKE9mQ/Tf8x+xKKIqP9XcvD
0PM3K33J/CaxNqZuIuo5qPaOCIUpx1Vzreajoy++NeMWNcfTAXUDP6qgcfyTI8mfiTXI0cFGqlPw
YJw0ILE1UB0H/dJFhWmRF+LKWi60k4f7iPfFq5BlHxXgR8xUvKEmrgbrTCM5YthZUroMacXYlK6p
AH24kmk06hW/OvDM7Jl/iyIDvBRwKnXgNPea+liAy3c78ApppnnTVDrfjGh6WBs3eSr/Fq9IZahP
uEYKHekcwI6lzK/5BzL+Mx4epoaij9kyBkfvbl+QEmkLlvVKOVRE+yx3I1GUfHaxAV2ZpQP61pWW
MkKORN9hY1HS1hSDDpQnQaoNQFELmGVN6gOFozDeCboQkypIiOij73tryqj//D4gcp4mPbNltJ58
dM6w4sQTiUNRlQPTUbbXEFhJPFRnVkjcqnb02vvZ2jawfenUR+Q9neBsZE7oKS3YRBl8CN4C+FLD
1BLwE53oSwnymbJf91WpqRIyKirL/+rppqpFnDkE/I2mhl69158i8OLPXT+NDUGJ9g3yF9MnK0p/
LxnJoeKeV1yP2nmFDZg/2SkN30APTBRFj+27FJQAYHEsX7V5T2oCa/ZFu1uRwZMFv9romeAz50Q6
hM5iF35RHo+0P9Y6zSi54DmCKbBqObVCtdEU0pDON8riMC8Hf2Z0QLXMKbiM1BEfDvSeWCCv1ct/
h/+5UCUP7KSZRgx9jhYArv18YofA1mXiS4QgKAc0WWaRP8kx+se8EZMFVWdqA7gBwu5GXQq8J/sa
pe8mHzZcxyQtx+Zh8HDpAjSPGsT1OuixUSoYri0QQD3BUfrDwqYGfv9ZTctHUILMul5pvAEvYkuC
g7T0krDv/i9sM1zeueDBlvbImao1Na3byU9+0WCfoChZqIoB3Q2ak/TwRu0m6PC5a5yqqGc5u+cO
ViLX/VlpotA2PPOxvuN7QVhKgh8T/G6hPW4MulD4aFYB+CPhX3p9wvDubitl62zaC1Mi1qIyi3A7
wAeCPsEwdvLnAp0CabKEiz8qM4kfZJkJO14PykzyeR1PWgKcB8Ic2k0TgHYGg+5LhhP7Bg5XB/is
g4W76Nz6fFDki8qNIrl690nXqKToYN1ml3zYeqjlg2BgB1VX4tBhZTAtpAnLdrksCpL9dkfTxTG5
PSSwGEsFhtGgoa9mv/0yJP0l+5JkY3W0+STlFt2b2iziyr03aKZETtEB0SAFmGcBsi2os9VMWg4Y
mTBDEHCEy7JWCPicZ4vUczGkfdsWu2LtxpItqf/zUDI4nM23ACi/GeA439LLq8MqWvZeCAcMt2UT
ku1dfoEaMfMto3RQeor+wFTSTIoP34bOmK+n/VingWP53PNLSaRE03Y7tlt4pHAjXoFccUJgB1cK
+iafm8FZ6FZ5Om77Z+ZgCGOxhphrwnHq2jW/sIapUrmfpun3BP5lUljMqfbXjX612/7JjqqwL1si
0cGSMmn/fDPNqePJcTPgUlWE3NdRgggcIZ8DsCxHVcwkXcdwRC08nypljxUL8ak7MrxySHJPLxyY
Ziwo3HCnbY5swgQJUjZUXGUxt5sJ0BcPKNb/8uy6Z8rOTnAmCNzWY0JBPxIXZW3wxgKto3HEiWFn
LRup1KdkRRcEbltTCZulGEP5dpVmiH8800gTapSedGNjbJpFIIdtjR9leZhau+Q6QilTQwkut0de
syXmF7/mJdFfut+XlwLIHoHA3HQXKCbixQc+SVVvw10zGK2oyKYeLdtjyNiyh5/S47SNTyQKdVjR
RkTyl5C94Pdy1T5Um/yuDvS6HIwooaO2zGQLJ2MTRiDlJMMknv6fsH2RGWrq0uyaQvzVeBmqEVyc
6O57FyyjDYFzzSPJcsBSeN7E+XNWtb6XbhupbAO3PvzgCoP8kZdk7hpcI8NXuIIH7ceFnmekVgSW
UkA9EvtFW5Dl91w9uXU23fGhxmu5oKAhoJXV32+JX6FkUKoqmSerPBEmHmv+9DJGO/Z5hG/OyVOH
wUaBzBou/0Xf2PxwpXbcsC3xV1a5hgn/hA0PRQOHy0T5S7ezNSkwOsBO9zASNhkJnMIjY+2+DZ/g
v4os/cFJ0h+GXzb4gJmWH3Ksw+pcEOp9YbSR28HXUMbqh4UfHsWVPKTuDcwLi3DVYuT4ggy/opHF
QVyQMjVSTsGjG0BfDwW26FiOC3IwyJPuerU/wdahC9LlllWYHFi4MVW4Vl94kVnNFJhyut0FrXq4
qqZsQI37QB5JyEnvimKLCFXCfMEbQu10HclvFpfmoJiDeelP7LwfmmF4rcGK4Oa/AOcyi68LbsT3
kZps37g3mT/67NYOTzx+9TyZg55H3tBlDb50syxLqwFPDEFWdVecxozFXcA2nMoI4BmXiW4SYjip
6We168seEZMufIDHb3UdkaVc2ToaJ7BOPHQ5/zJfJ8P41ZDPn1asd8/eNhwRE5qlWVaCm8adLH2a
IfbIFuK1nCpNDUf/mt+XHgJ6jffynOsHgxO8qX/LLNcgTzgZ2ab220VV9Ss3HZdnSz1bNHs7U2vO
lCv9TMsmWe+4u4yxHYz+mpuvSoAXMk5hc8uwXJGFjdD5DBu/CnXIIVn6FOKVGnoMTFwPlZdL6Eln
D++eyHUL57OlWChEUejNxGn3yx8GuEqvPVoIehEZXlDTg5jqO4xsE/0V8m1ZKpNU9crVNI6lqhz1
togz06nsJahK0UEA0ahcwzzm7oqFLdJzyfFVvP0k0cjgBkDzHPc9hW4pJ8oWU9MOvaavsDxoeL6G
Z15SyOEho4UNjekaKLgLKw/MsYayXnCI1fHY4+Io0Rq6LJBqbyXa+kR2nwTww8T85LaGqjIrXxka
EapjAejr7Ogf/P9WgXAZJLiuE4eyM+GiOL6+OFZ8GbDKrxJr2B184xq+uQUjeTHem/aY3UI0yOfu
zGy/mb7JVExiV02JtsbFgJ4+TzDzDMplyHYiPYkqYazRMoOYbFEqCp5pYsU2ar84BIFn3V1dmvPW
bCHK55UtMXbp1tLQfJ45mHsw9bqcNqLrwm4Eyldu1Rdpa5aQ1Is0CTWxdObfyb2zETTPgkVVwufd
jtMD3W97qhqlsc0bu8aUT297alhMUs4G5QKM4g6/lRiNhypvNPqHNuJtWYfOugpxuT4KhOpns8uD
UDabGAO4PzbhsoCqAR9UC5Y1gi7DG/SfGLz94cM61oU96VT3R9tBGNWBmpX8PS4OpyZtw7U1q1xF
DZ6qAwA9zXtmnc6l7YCiwB57YF2NI2el9wvTb1udVIl2+qjqy5zHv+lPGZPqYFFG9mGTEmXJ/65U
1WZchzzyS08ollW58Mh1GeaMoJLrbvpgAu4cCZ9gg682L+rDokP73VD9FRoON++ab1GJ6vAE4ClN
OoHaDzJXCPgGu+f/zW83LBwI+xjtYoPxLqIRYni7YH37M/OsJNE8c4AtRHM+JRYvsJ5mZdrKfZWY
UGXKRcpUG4F0RApKQpF7IIj3wAWyOQlvJ49lKXXcnc+pXKaJLJJ+b5AfNo7jydbVvG8R6H3FTMQ4
aojHygWahlJF0Z7SaS057fSgBkz6w8jJ51d4m0Sm8TC2IKa5P79GcW7roaMmUpejYHg6aIUob+9a
SlsaW0cg5d/9Xsza+KERK5yILL+PsJ+GN47TW8aqphu2CasvILDKLRlU0Kfzfh2kOYz+qrO+aWDA
9wnf8G3ZNPiAprukY6HTWJTaUkvztCwObeZAB1kPoD3dQ+JurPcH7QgU9ArwCGWonlhEeKz10Oyi
HiapWMwxcV6fiGqhS7XFtm4sMAk0SoahqpkzoNqWW2p1+KZPTEOD6NnKWDmCLdgf0vOvOjpGaJaT
LtRVlQRnXkxGAn+h7aD06t7eGH7QHBokwmuPEvGEznH5my9Y5NO1MNAcUCqMISi0OaOoenyXAxaJ
pAnQIuVZppyl9GbYh1M5TZV1AQaDSguC7r3+5mayZ2vAjRSrpc7BpAOk/G+gNQsdVCyUkTh0oOLA
mvbevQswQBgHm1imk+pcPwMJMzFeTmFYQf4DDxq6xyiUDqEoCKcLJBZj47ZseLHNP5f6peMS6kh4
rZjOY7LIJjK2/YP5Xq+7C+WsqJoaFPEAL20kXSnBPKqtUaw+MKAFxbTDLHE3vZJ2qBJyHQDyleup
g6V8tMJEARccG/tbaWjy5i3Bc7ymBXu2heKCKjhe/85atS+KA2LmFMQ/xrx8rskn3BJaLyIA1TIq
Vfx5qe16htH+yCL0W3aPNni3+XZijjchnp9CoCHhiD/VqPg67l/qvAUJZqBpkPQ8JkYP4gS/MY1a
HWsBGPp2b/HGoPvAkhzQsTO4531OPXAmtzoRbXihupz1EHhd2RvlVEF//4zkyj1L+mbOj5JqQ3l0
swPInNJBmQVISVbYe/7XVHiPVfnY4hVV9Oa9pG1aiZgQdt1llm+q+VV9MkRXaY6SjladBIUZReps
F5O+hZ/p+HjjKdZllfCEuKgcl/Ut4pKVaa4aejg7Y4hhePSSq6KUj4gbSB3pmKLY0tvtDmdSf2IF
WaRYyrx6yYX4QqapQ5jo9TUJWZWOG5RtGdTL90NDyljPftEHrnM1pFrH0CVdxHTPknX0Ig90LOT8
q8U3PUUXWia8L/V8ckEWMkI/FBSO+meDgCnA+ze63VpGxMLuLWKjC+DTJ/SCCDjeIeneRh1h3lQC
WJGz5t8Wk7RNxXQB5A0kum8OBju6uv/6xLHBwR5kpnctFqQPFiJcEElmKeakPRG0jFMtPX6JBUrg
e7QUbzzL8O6SAThbUPEFpjaWMy/CnL5l2kZ60rqpZeUPJIvgbXWIHlyQ675n/ipzEg34fxAZLBaL
/u8kA8FYBSKOGI4/kM7DINeNZ+mhueMO1/ROD/alhlohVduxgs2DnzTr61CH9fLuXuGwTYKSRvhE
NnvRP6KTOX+7ViNJM2ZJavELv98Lxp7H1qNQbylJyca2YMR92cpvFCEd8fPCSXi9LuT8hvsnPhYu
V4iZ5eHC6ix+8LLIGy+rUJgh98OsbO4+MPuQufEPipLy8mVlnrcNRlb3XqUdaSoFUsZEhBYbgE1C
v/EgNZI946sPmfLhPc2zpysDBt9YLVLPxWaa18RyipDHegoxjnjk7xrxtxNVYVl2DhiOhYDOcECV
hzKMyVyBBjv1OEZrpHvo4+P3Hk4IHE3frVWlqTNKDNjqcd/usQ3e/F62h2/0WlmnQ4wACFBgb/7H
tHXQc0tnH2nsro9tDA99+kqiWeatwDh6Byr2NLdLxc3w2yca3+8AqU18vQF1OeI90BWFPPDZJ2Xh
R/hhf1FxGE4on4MMEJqsOgBazvkENFmCN9dNfKutmhbWJ+tC1hvFwKIe9z4631heMuV5mEU1RJJF
fvuzcPMmxofotfq1Oe8uSqi9hC+slVADZbd1zJ+08r8+0sFytL1lLx27bkEvXowlriI8Fn6bKQY1
eJPyBuO/GxSWwJGVzTlSF2E7wY2GP8Pk58T+Qvwq3ABe/ZMVrL80/QDkbqWyRXjqMhA2lD5csE4f
qT1NAxsdXB9NMWSZtf3MLmw39jV+mb//n5whN1lXJGBASPsmFYnRxeENAlbEvrebu1t9UQwejfTo
0wiWg9my/RWipJEP24p+Y6UZYw471/hu4ZqvSr3w77H2TxBWFt0JPNzxGC0TUP/wp+66DyT5u4wS
JEXDyqJPtJGu66Jl0W+LIcnaJiGaxZxbHLVKgGCYwOhv8X2MRht03djO2KHiYXfbUgTz7yivWu+4
S+MbkFMcs5k+oYC5j76NoNDCTuM1FlRgWsAO3Us6yD4QmJoS/LM5izApiojcLpXmR7Ys8rghEjvA
JPcWaXrLyl/gG1MMxBn+FT7bxbPfL8cF2Gtj4pNF1Fhv/vla5h2jUoMwSyP2YAqkKgD9/o2Ob2fy
2CeRiSYNMoi7QL/ml07dDub30EeMtq9+nAPC5qIGahUiG7TYqo5345zWlqXihSkv1RGX/ENPi2FC
636rgRZqma8/qKCeopsKloj9iTvZeGdaeBy4NUkz2EK8S80Hy9UUW0kquzxH6n0UoEB24sVimpDl
VyKLXpsGtBfxgXpTTXClhRsK9N7Nf3Z+Fdbsunjq7SG3Twe7gVv6Hb1FCcVKm2nOish+PWeH3Exp
AtqF8cg1T5s+7jB3UuR0gFpI9zY2OKoyarfhj/k2rS3By7iwjQ+LCazQnb4sJwlT0qx+hECYOBUu
h0wB/Z0A8zLeCwbjlwiKxl7mhKqjW+S0UCj6NVhT6w+dO4u358fyUxT73s75RMZNjabbu62qb3Sg
Ljp9ZbSi0L9SEPsVt3dweEXNn+9Ie1Zi2z+5XO9wxSLs6AMIGYfmaWhMHxWkQ8jiN8euM6NqUmAc
I6J8gIa9SLkF8d9VGwQWviKNG2lLxCiA+5bWUP/zERY6dn5/rLlmwABlSOydwODniJU9RYEX4KVi
HLq8vrk0wyPDk8mbvhxBQh8IbzvxpS+19cGltqmjNLyY4w/AJAY0PkftCiJEcFZ1GGESZq5iVlRc
q+k5R4BDMMDg9ucYrpPyMvSj9TAkSXIEi14vr3F3y5zMLxSHZSvUuDoyDzZowj4EwX1jeEbue/7D
+t4nJmj6IzPm7rH4hDyaMePDHj5G++pchejW4zLNsGuTh2uhnPz9mWCW+pXtDsIkrSX46Kw4+nJM
lDRmGUAInKET7HeQw+g9jvL37JJNXHqnzEndK+yisZfRqanvvCacvyS35h4iMA7ZfiMYsvpy82Hr
PVkCzDVIKus1NFCBCgRoo7VF2pHwMyvAhe1v3uUjOmEd64y7KYP7NOA+CENNkH3IIht2BuBPkzQf
dKIxhl5CaFMRN1caYzPDQ2dXw4nmhPYUcfUz1PyV78u06ZFRCzMPc1RamKGJdMcS7aWqHXbiM5r5
/Jm67XtwsWQDPmGLnm5l2Vf4MWxW+NslE3okvmNq9XBYn1d49P9a7AU6r6armRpiF7XNrmJlAIIL
vnmoqnCH83avA+r8vtpXU8+F2AnMmg3VQJmg2f0F0Gp33TpL5uu6UnqeKmVLeHUrb55IA0c5pKUx
nRL4J51GlCTzTkbJpmgNsN0ljLkrMeoXlHcJC55aaOYh4u4EnSV+9cuI90Fs6rCbRl/tw89gOkHp
xbSpUMrJGUtRieUbCYu1XwskhdIH0buzwr8celCbQcKNeiAo8cO8uuaWBkMNSe/b04Na4qUbBtCY
uK82hYkrODtg5KG62vaAfq9yy8BOnrbaNRlL1z0DSrNWutoFrswxkEQtOkY7T68HqLF8LF/QzD1w
Nxwk3mF6pz1LN+KcV6m1tXMk+1+S5O8qQW02NNLD17sKGv+mWLdD+96JSvF5MdtC3qUxThk9GWTz
mT06EH/A9p8DnGYJvSRfrBlhbGaH256QbZHDd2SdCGCc2nKaBgnnqkD/hpjdv6QWrM8/wfio/p14
hjS0vGHyHAsumo/C1qGq0J2mqx8+I/73xQaln1+D3ALGoy27HGV0PT1zzCkgptry3w8rOQMzUbpY
+PXe2F5MITQC8/Pv/pQh3P4aua2AP9VlRqxGDovmY1X5cvFirmqzccw7b6yW8iUqH7PElfBnjFvv
cwHCvXFQ4Ht81n1I0DkomtjEdNFMsT3AKo78+r7MG6VGSQSu5oZuo9Fam8Zw7p8j0lXv3cbp8mDq
qoQ7WJ05U8fylG2PXCTtu50kIGSSMF1+o/keGxNitgAzJmpt4QyQ0FnxGRvnY9LeHsgVcZKDB77J
bWTCPH8g7UUg1K7u02g+sL5NOT+BXqrWU6BV4a/B2eIZ3SCDYN0lMcn1ngzzq74xh40zahIfRVk1
FZ5jsTr/7EZFJmbwxI7eTqgZB/tDWGidX2UaAuC9A25TNKZI6fFAH4eZjEyzqVwr3eLpi6XOlPOn
Jb7kaerVp5BGsoFxxazdeH2lU5ZzwB9MUBilocCCBdsz0av1LxIN3YJWlRk6mNomi0BDLhO3FwP5
GQpRndZrlBy0lSa4Wr1Fov+Y7igC25Y0nG4QWItR7lEJ/YytCzHxrUEz0btDh+0spxR1Cka3ynfD
A+P7WNewWvx8pqwpob1vjyYP5ZO8wl01hSJ6yAVrSbs4e5LzEJ9p6XliXAEB0NnPnNV8PJieEBkf
o01qoui0MDirpKXZsakYgHCK+gLyev3P1SpOjSgam+QeLUH+2tRK7B5NUpcrBwcwtdSru1dFwCZD
CV7I5VYQtasnUBZYbLsM8ZJRXSsbl8awS8J953UrkZRiK1rPJRQeV60QsC3zwyuorLH0rfRv8qdF
1ZE9tsB1KoK4t4MIcMWWHZveiVuLqq5cXJev0Dc/4jUl1+eanh4sSaRwRly3WHjNIdM/LpXa+M+C
sjRegi8NkwanBqsRBRdWfoN82i7xViVeKABslPjPbvQHX3um+mEOi6MOjgjHjZOy7nyt2q7V19ZI
lzsvuN3vz2ih2Em3wObeChfBE7o/zVvVA6c9kHehjEFhZ+/K2y9dNmX9eexBEBDY5wBXHZYhnPuv
IeRQwUUjNfq1YkWNLIlQPdrYjE7120uYA0/zdyKwUu4bI+JLWCwso/BWbuRNSsWuS8cbiLLFYxcF
yOPLHp79/n/9e79HvW82iRgZ9qek2iKBqNux/HbzPX+DW0c7OqVvissHmyjv74HD/uxJJuT1ulmV
IKEYgxn+oc98qiW3/Rk2S1Z+mwluw5NC9duiXKvVNDY3DkhihLgejO13g7qua4N5FjH56R7lGS6J
Stf9ux/t+A2fPwGHGd2jP44DKHsdS0wJc/ldXUimt/+PWgWdAfenoqH7voSI2jbaiEvDBe1SFqUc
HT1qC7UP/7q2J/ns4Dim2qGHQTk+gew/A2nIRwAM7cM6Z/9zLGmgDCno3WGlZ1zbaZ47UYNlWtGA
MdISUrbuTC3CEGnn8S2xJEAFdtz/t+LtpHkHZB+Rawp49mAwk3acQ1hLmdCpEQf+FozWI9QgGvQt
+vYwzjUH0/Ouh/PXbyrpzGNaM4wuJa/hxaCHJN7VVD3HdjQut8o/8iJw8IpSqpcgbEvfz+ETDE2g
0XGh9QWaU3VAgual9K8xty7rPUvsBuWRIlArJ3Kab4dBbFQwoCpOBFYGxuuANyrMJVfffevsXr3t
KTSxl2VTpJVQ36ha5FUvdlDK6C9nxfruiNhZ6DDf700FStUr/B4qbOpecK5yp/JSxRT2J3gVhKih
kHSdDqXDk6msxYaKr/giVeTw8XprBPTvB2lg6AySOekt2ey8dwblmxvJA8g8pGNdUABscSzPyHU6
pemgr95q7KGpHtqd5x7JZGvwKz6czQq6elnUqxQeNz2Nn03Xvry4s4ge5/M8jtQ+V0B/a8U6vrqE
rv6EOYoBU2gt+smUuiKkwZksaPb1sZmXrz1XNrrZ9jlZaNplqF609TzCmDwGvgi3VpMESMMfNq6Z
9qSDt/IPxQwgOBtLooO1289eGs7D6dsKuTX+JyY4JDPJKQ16nkp9cjbrxQbE/FXG4Ru35UxAGpMT
iQXrteieiyXW+8T6UIy+g+SpA5iu+Br7YN2ZhWygZBdU8nT2IQf61Jo1E5GFMhgnDY+PjwkJphjv
cFs00OiujK4TjW9RqrJP7U1S8aIR77aZeByoq+w67cLJlklaYBoBCMW4E7EFrKnY/L/h6u5RnevM
DbLcVynd4xScKRNrPFZCvjQaTlZDxlsfCjnK/m+OdN7OdgLf6lV2yhFR4PCp+d4mkoQ2vje7j/5p
PAKWvdJozZTSWiRBHryjMDCIhE+6HldhylFKT9cU0ZMRsk+wQ9EDhwDWJBaJo1vqAX72gMZfxvdU
weB+yM21aP9Vp84zMyqOqDsr4anbumxnOwyBELrCbI5PNGf34hHyH58t0cRJTDUCZNlhTgRMRI9V
zMy1Xu1JH8YkWeszurBvOPhrQqiiCETzZUu3ooHeV5lAdzyNolM3lrKOv+6ti5yMLPKNYYkvqm9U
HD8rVxxiiProtrcdoVxN6RSZblYgOjUm3I+2r1E1ByENNQcrPcvPfLm3IfqE1Fv4URHDygh1avh7
19DBX8qXLin9xleWte6vOxb+wnJd3BhF8T+MmacPwUYs68YJK2XRbxDuUiF9gnPXY6252Ui5c+Gw
Yu3QeVOSan34UpRe3tSIj7V+C3EbBE/BqCimBke3q6r+pSaDnrzLefXpupkKKjQg68qwHgPYiIST
GQsDdyZ/8/581gAHQdWxL6Z369qVmJKOyfib0UL7WESqUI6raqX8GOaob+7bJ3PFuChqZbVUlFVC
R/90GpRpjBl5cAiCj6QOIMnrvJz8OQSprE0HexMzMXIWQzfG4zJlO3R5W4gSwXZTEd7EwVt7MktO
ihGLPacOIyeLuZbOEtweLmTlzbzAcaT+2Mm/DuB5yUqLVp7lV8XqTloLVOUQAtYpnyzNPd33xCS1
1kuWCpLowUoBLfAEMlFLhnU1rafgx8l1DgVuvBMRs/u6pvq/yDXNaxgUL8iAh/KiABQ32gmOJ7di
jqmvkGu49TJrD+RGdhBVUJbwaR2aTx83BtXGF1QlY1qeNuLlEi/1U1DeVWGQPsMC19N/mHzeEJzg
UAEV5MLyeLQp7zfNW6vv0x3HDEID+3V0D+gD5c9SUcVYqZbhsxl/SH17iX9zbFbB/AdH3sUm95j+
/IgpftGvehZyhwFJDN7iU6DOU14lTiy0PBCFsL/cZmYVa0GaRKVRsSdy1OaEtPNEY49PkynLeYcu
YHaUlLrqkERDkEfYRH9bk2HRVK8SUVg9ozZjuGczi47DpnzIgBbP0qv92lF+61Pp+ZbetLSr/ue7
0j5glBo1taSIg+TntH1EI0/iYTwohXfSLmWU+LAxApxFLWP2dV7kM66DAhxUEHlmz2L90ocBv31i
PN1hDJG9oVWwb98WeN1LV6CUWfkbyjRUMjxtyBB1UUQP3jkD6uHp8t+Wvgf7NOZLmibqaWU1IS1p
6yVcNQuhJemie+pwVIhnm26SRgZOuI+IxmfwL3N1xyCgqE6RmJlfBSOBEyWsmL4P717yeJnLtxGx
YOxzFPqz9JOHy1bQPwyZf5IYbHinCniq2hA4OCeKAafjKyjns/beYWJA1PxB8vgnfG9HCNikRsHl
OUFB2yerTAR0EF4Rjp2CMNy2qIPazXDDfH0Rk+hQNGcMLRT8Uh4zz73ewcrpemyoZmbhlnQQH/JL
450dpRs7hiWjfBb7Fi6qBBPHvSxkVivKML8wcrV9TUxvPM51P0hsxw1sP4QUIQTv8ZWrBO1jy4hm
lo9CFgVWoyfB4nlV7pphdJQOb8OI0B+Xk/6b1Y9ElaBCVkGujfL2lYREdHZr041HSesLlT3UyjqD
xdozxOOg/P7kx3BSSCFyOwQGlMD5EtGi8y/MBaxB151CeXF7H/5MadQpCbYrC3oS/GnOyVHaInGd
gwITnIxqpE9qfd5dQZgRvrYSB5DCIhc+idcBar/BMEtZ2lO8c9yq4e54gWrbJP7jsg4yQ1qrCPsM
dkKpeBf4Gri/UYnxAD+mnuqjQY5cRHJzG/IcfMD6ggYJkB4qDWzCjvkXrW5rqESsyAicPYwOuWTa
Olsu1DCw7QSp0hkdys4uImPVtyAmNzbU4B6XxwPNZiwiTJquUqyklLIdG0dq8VkArUV6c57eG8Ng
rYoTFpMjI7KOucqMg6Wwk24ZpDXBEXYgPOwiFGVUJdEVpo9++0EK0Rvg7LjFHXA5MutAof7r6MES
AmQXLP9qD5IDYhYtugkvujqjcxB9LwgJ5XuUYd1ZzcmbQU2BebXivOX07yBsNiM0OYCK3on5z1Qn
1SABLXTRzCdMCTM+V6zbZ4mytDqGrMyaGtAmwYecV1k4Jcovoia8HD5B3EKMXvHxZis0G2os8+Py
+FKXiODKBqUsNUwnyDtvuxwcoRTmic1xytxD30BfgtLEZSF8QVw+w7rrfePpjzO0/xePugrnPq03
Ok3NByvAUNzfCZeFCCXNpwgiIZSE25VInLscd3sqqxQLI+kf+XfQkylQCZqMd7/ljAuvXrLoi95o
AQlGXRBCtOUBjt4m5OdqqL6LGMV80hAqfBjmR/Vj9xftlELoo6ECQ3+M8BPZJF8Qiuqveyg1oQ/I
ksbXiubYfAQ6StyETj4bGkdQz6oMnXoF/iM5OtJyYMNELogtQNIAF2A37d/KFmNjqWmtOnyhAuFw
dWAoC9Io7KzIrdRtzoBnI9epys5fy3//ssstsHPvdD94Q1QrMDhR63yxrkOI3rpe8Hcvf+ofKe+6
a4We7Hw5C4DjP7nkjTSq05rDR5PGPuuc40fcHFUmN8Cc0K8vXC4ob8Tnu7PlCc+qNd9uhoo+JFpV
xp/vHKNTMMDwXs8M4eT++nxRCsEnkCD43trpuyUrFx8VIKcvKgEm5vxew5oRIQLf3jGEwzBIgleV
xowYFlNgRACKgQ8QQ+5FGots6U8ekjsD0zNU9maIRBunIur0/er6u1Y13J0FER4W7YQScDHnoPC6
7Gox0mTEydCX8RxnAT/vcvJQltDL/05lsA2N7aMWMGNsJbH9z5IdWxafQ/fdwIYY3qfBKWHEFjk6
i7lnj6kj9VHDV2CdrRKzq7DllrZCKY5WviDoJAog5x+Q04OxTWM9JLOZn04hSOh3lwBaBimXsN/6
ExWDJMkJ/Fq2pu6FG4I6LdhSc88Ga/1OQrLHGnlX1pC6wBMEPA+eGQ4GjSV/EZD0TdVPwEMIqMBE
0LEyGqEh3S5ZTXTkPWgyhufu+iyfaZLiy1vGQQnbGFc6KBvSD49n4VJ7C47KKt9s9Qq5jzpM0X8o
bHR9G6uXCa64SXTT5ig4IHa0te4374F2F7kF+xgmfRVAWQ7oZ0jYJFv+WO1782kgYPmW9CFihOT7
NCJrDqWMeSNXHCtCWeYufVV1ZMexsf6nk4hPoSnW7OpKoNjs/AEe8YDDyUoYK4zQaInbrZHGxev5
LV060O0DKQNIkAYuVN4VKGHhuGeNIsWlej0IaL2SGNXbCAvunY+KWW2iBR0++hnCUbyf3Pj1AxPt
Yv4AA4iDnD0KfwnPokj92aKI6sIYa56Dfi4OsQA3bOPnjhxVjJ7aEZ0y/Ok1CD+8HadOB2oeKQnC
lrvMY9jhPAGVZ2UgcJVELlVS7PEY2fRU20MKrM9uB0waIQgI3SF4jwyuuNfUsUXrnjTIZmUrxEJM
eiOvVXRqxCT/0jt53meq/TNf0somSI35O6nDZ8LweOB/88orUooDAlt9qt5IcWKgKJUEc33AYbBY
MJ86PefFEiGQMaHvovhdfZKOQXu8ncSrZ5cDJyjGzoV+9fk2uUiNL2QrVHj37enZodHdLRiLZaFm
PSmdFpETLuTw8KNObsgXphT+ysSjnGdHRwn4nxVJ5q+x3Gk2SRFY0dgVPSXjVwRfqOcMvVTzrWvI
wJ4LpXSjchDo485Bhsrgf1idJr5YSxEGotSZJLsGMpBhTz37aq2guJNwV+bbbBwuLimlqHVFqpvB
3gUxD9zA23bxhQYx8Du4xG3auyOOm4mahz0KTRVph13BVFpXmfmgQGSSp0dJGnKluzeqHRlsz01s
fT8o00guQGOsjeCqwEP+5DOHh1gykN8OxaNqUYE2BSI0ZAtF7P7cYXh87+1JEHf4/hp1h4lgjtHj
7QmZx0KJbULlGx0kc4VGXWlUdI1z6yyx939mZnwjvrwph8n7X6At8TiX9G7g7vR07MF7mzpg3GWW
rd77ytnZE2C+2Z/8Sw6F5SlQStIc7+mqu3MOUULKqMAF0Ag485KIxEDmDzpsh7w5mp/Hztu19Od0
BT8CpI47iFqDzvpzMPVUBFn8/LKJRb9+G1TnStdWbJbp0sU6aaILqtUoDmpKCSndgzYhScCEiGgq
BMU59a6+OiFpUnfj70QAjrkL6kRxxJ42IR8CDvANesY2z2OM320YBtN9a2IGrWI3goBgNHHOpvfW
B6CaWUop61WjPFV8NjwptdgAhLW8W/y1DQoJWUUueb4UpGknLtOg9WlTP27+yy5CdsXLHw1Qe9VR
3N9gXfnYO4qhrExReLFQ2JtdufVZgVOrHS1PmkJjLihAoNmWn6YwVcZJnjbria3afd5SJ8jdsrzd
Oxibk5HLa4gbin+HDRfrPgWp1m5y1j1+ewSCuE1qfX0eSYjDkUB05AJL9jtd1d5RzZ85I/u33hB+
rJuX34CBqBqpZDt0RV2jm0NBg4n9FrGsDHObZ9xZekYHiaN+D9tjF4ttGzeRT/3OCPo/LTiKf4Od
FoWKolbWsh8a0c+dDeOUWNO2LYm1KYDwjRUTRXmqOhP1wNGWT6c6NB7GjHFnMe5kLpUHSmHRReQB
aIAObM9sqKf2LJa44OoIjzZAS/DlSUfTmSotLMbXGyxnV6OsaOTjWR+7SvJmR4lOCWE1cDJJh06K
551b3c2udYCy15mdNtc61kx3iu4aBnr+Jqk13V9H+2PLEGaZoqHpBbWB1HIyTwQJC/pFDGMYTq6p
UAJ1GvGcFzolIwZjZ6mMiQIPpohAGY2Qd66Ihw4Ve+Udni21KJDhgeyQCqaHEC9z+t06iiHpsKl2
+eRqKnkgk7JKkUEuoJPDa8Tm7okQ5vk7gmUw6EL8RoYtX7iETQTsxOgiTbsIS/9Vupqa1KkvZnap
MF/oXCTBn0la1bhve1G+lZJzd6RvY4UwoGh4vrGWN2Rorer8n9no8P09Vt9LDf6KvriyaaazcUfU
DoxaJQtxS+5sO/R9NOdL9+6gY+1z2jj6fk+zYdIR5gJTqH8HTOwV4nfFfIoiXMbj7qH6st0P+oqU
+9wcanSoDCicCjpD17F+je7WGeFGVPs453yMqP4Rwb27w0OzNnCf8XTI1lAGvbE6PnKeHYgB01fV
BMY5y+hjBXIyV8zTGUlSCu32lFeFs0nqf+sLV+TiTh8TY4N3tEmm6Qu5HL5aImmvbTa7Jh1yeuQ9
+ulsYCx76eokdlk4XAShaoa6g5iEaA3Gb3OpltHA34mWIyjg9ojFFaU6aQxZi7ocENekMg5AiZy0
XNEINbEwLsNT9AdyfFGVmmuDbYYvSkBp+q6Chgn9nu+TPRyU1xam19wkkH/LikR5AdMhdXL4Wijr
FQnXyvlurfYn/jrW+i/iLh/q9sW6JWxPzWvo82PVx3EBD5bAqo07O8fkQgYbxECjGSMaXZsv67ke
75WSGWPdbN851AXH0JiCT7jM/29yqcWcfn/RZZy1RRRmkBocPkdhvmYT3GSSiZgsc55MWcaN/TW2
kN6BdXKcl20De2KVe+72exS5uvA3f1YwS2iFheXMo7AWJ1iRPzu3EFg9ouMEBdhrhSw9aCJLnyzv
ac528huxFDjzY9gSHYG/+utZoinhqoPG8Au6aTrqJUNyrKtbhpw71ZXrEX7giVz4Y9kcSeH633kg
DNOX9eRtxPzS2tNhFuGu/Htr4caqM2TK34ANTvZJVpeDuZsaN+DrmUEHEmIn8bqPTPGgw+8v8/nC
hPpyFkF4B4fyoEPniFMbKYsIvjGtkSeFDebg3LsZF0Eu+1XN92Cupok3zCQvRpAcCEWwL6RIw2I+
yMhczOgb7hT5XfkeOz/4Ms7gmIYZBadhEB8cMmpt2yluVaePCFlUITJYlzjbpk7LAAXfJjFshYKe
EIY610CbRFo4nSHlr2uOPx1KI8NujrWosHfTjUghsPR9xpoJFer/l9Z2MoGAN3aepUzp19AkkWA2
3KBXZE3eesDqh0F06MJ2kRdwbYJLKNtXB10yeBpZTdxT5YF232JssSo+SOin+kBC6BI271OrcDEx
wCG5Jo+eX8EQGVKwQZxUexhIMNrSiaLJC+VEbjZYryNWtko6fqgFcR07zSFiY1462ydMwbCJYTP+
898wHQsOG7uRWbx62ZODprNBeMcggkjQl8VazIj8Q5UP7T1TLgmoqp79SU+0IH0NkB2hJ3xFarN1
fOl6nOVeJd/wIGvyVjuUpDg/7986YAM2tMwW8Gu7ovwE6VKgW0h71kbriXDNpgLx4ml6DGqO2BWV
Kc2c7ym6YZweUlZKz9WZYHlCt6Du6aAF3hy2scVZGybPtcvIYNHxKHjyQvtd7SWIVZjMmXWct5d4
Noo/Kz1xafVno5PTxVqb2QLdCrO0C9wn6Og3YqaawCDtdFQ8cJ8DHYe1fxQQv6dlPsbk1+Q/5Cal
tlTtXvhXzZlgJDYWzDTduIpxIR2djADslTqpVGym1fhpCwo8tcMj2Qa+SrWrv5pcJ/B07WlCiHYA
6dN8gvYM0SchUKNmmuTIepig9GKnB7ZotxEjDfD4ccRfybwRbn1FhrGtjAUrMk/i2Y0+ewb0xP94
LaECA5GsU2dyq9+NCp+kRdH7PXioCJ+b/MHpDDBs2pOs2qtAAQsLDr3EBSZt8HwSrqQTDuMuKMSB
QmJMeXyucAWKNORokbY2MZLR3I2pBnDqa8eLjofJkoGmc1EJ1a6/FsRky76KlVuUQWCOTShG073F
QbC9tvebqKCfus2CB5uNAXwdYngO7AQHJHVvpZ5ZFdBHtjF5PFHt7XKiB45tkHxwL/K7Zc2wGeLS
jtDJd+pXx788M5ZhNE9xtshVrDxDQ8zsmGkyzLLztdWf38OKCpORrl8SwpbslkYwU+9TljO1xsj5
BkeoOY3qlO7ZHwVlHgDGE8zQLLuqrWPl9XIqMtQdWNntXehPr/e8tRM3kQH9EbIU+/5dAW7wYoWX
/TPdIknEFoVTz71yxIkjv1dbNSb+qwc16zvxwQ0XgJLdhv9PLX7Xm62ZtrbWEycz8yNxIETL3v6g
zAyHAQP11jSpkqHrQZ+7u280RFXGwPkk8VuIqKZoK5/Tk9tmLnZFF0QP10qEgJqE3C4NK4xdb2uR
LLp/17TW6nCV77oalF+ZOc3aBRQUpqfbZkH3CTExKdnQhusxV5wRyzB/jHdZ6FBJg6UbkAhPfGMF
XnLYbqomeQbW8OgOlV6UZyX6HsVwaSgjYkaKODWpVmyw84Uc9Q0yi60yraxxMD7d3olTecTHI0lO
LU0QpZv2Lo+4I4wwbCeILag1U7y3KTGTEtZh/r9GSrVBE9NEhnWm7XryUIRwkpHE3HI9yGazszy1
VI9fuV1WAe4135YjdryevpS93FWJ2xoD1mpZ/O5V47Ljix2Y4/+t2lk1gxBqIkXHaJoXlG9SMaAv
beGNDA/JX8CXAMAwVPXRVmW8tGiJccNj2KZJE+ryZNx+MhQMIoDzo4mWHYIsbUpFPozf3GNJFZ2h
YKKecBU6rMbbkw9PJFvLmnUo4xeZmcyfCSlhMEq1I5kPiGX2KPX/2Gp58sIORROKEGxhq68ZQEgp
ZyqYVHSKodTafOdaQoW6MUuI6GPUj7gJHy1ZfAzXCnxEVzMl5t69oafM4Ozyn16N8ru2U1IxoL0h
jAKW/RwlH93iHUyoP8lsl4yOo+FFRT/6JvaMxW/qWsU/lNWt5B3F/AhCdXdn3PRk7U/6ibzppXmu
j9Ihqi4m5bYZf18ryN6VpIHzNZCV+SODZP/0JEm6Sf5ITVPAV1qEe4MVXQrwkbDlOCUJSjPK5K7+
PeWGFD4IJfNFEotzilhDkE4ePG/E3BMKK6I2yloaIs+LpKn2SdVcve5b/GGLbi5JpkttDwxcE3s3
4nlFuVVURJB0Vc4s1v6eH6m90AY6p8qzpSNEzU7EbSQhzOW03bGrF35175KJ0lvpBLBeWfSsr6Ms
uiyyyzVhPE+KW1Z4QVuJ3r8pNHTJbbjDFnsgONH9c0HalDePn2RRp2T7zb/b2F/ZZz3SXFp6WR9+
JrZtj4zGAisVbop2QocBXSgOirhq18dz42qoYEAsbmZ3FeKHYuekm14Qqy7XGCxiwDQ2Ji5BZAt7
w9h0c5RYdBy4Z6ScMdEVKqmTBH8dZXT+42qIa/W5NorPkpwoym3Z18EuKKR5t/unESJHux/SX178
6D/ulP6Ti6/cHKbqJeBtv4JLgzQyS8NtAstbeOGeJJhLeRmiSgARPgB313voZc/VVZIWdhj7v/B0
vYNpw2rTBYTk7vZw+XuP41BHCxICL/7QuOBl1bgp5+CUPF/EtCUJ0jZfoChzMRs/YDDjHqW+yhd+
xUc9ZJHBRTj15mwbKqgbuHKbmz2NJ41Xk/KB4QG5dx/UuHYXZ9fLcKRj8Abw9z0Fq0cvp7Aw4emT
kBw97fPQanIThcjpZmxayhuSk5CIhGUwqOkwsAb+Y0NQMFUKtod/a5SAC2VCmkCYxwNH9tvuMmOS
S4RpXrI3VEKcoxAvjJMXxpLWidvk08VhpEM5JD7pBVj5cAOKQvj8NVGLbfmmJuWpGDHEt3LZpbxj
6LrODQ2CgiPkb/bqFF46H5qc3Ykocw49FWl5kiMG9BYGy/F4wz+9x177NnAIG2Y1JHhczTcrg4aV
bjReJTz5bnaofagoEmVbjcsKjOftXXdbs0UJeg0Jnd/oZgZyxAT5nW2IEFUE9GNYJKfA1w+dxSfl
BtR2Lbs1cnvnOi/z3A2PhbCoA7Uzp5YEh5nHumLITmAxaWqnIa8ylajTNFg5YVlU3PICUfpAITrY
oqy20G/8FeZkn/sPpbSITxZduYCXBW9yv6hA8aylOZkqL5/TSIaOtXs8KALzbeWPmVtNlCzYU7s2
1xNNcXCFQ0cLE9OF9QisbVDC1lCH+nvcdZxvtK2tYFmMcGyUhdb388J256Ao9zghHd/DJY8bmqyv
RLW3ywlaFHn8kaQWlzF/as+EXO8G6pOFGewgNWIiQNZqrJqz8LHVnya1yTn7nfohDz5naL2PAGam
RkSceSu+uTw3L0ppuvlZOsvI9E0UajBbyhQG0AZCxr9i5dlB284U2UyqOEzeDZAM7I9oHLiqeB37
hs2gZRv779fD+CiVU1iVx43/h54uMQ+jHk/h/PVoqfVU9nF9OOXfgZHXkNH/fjbgx5yBsq0IsD2i
/uCJYZ24L5mhWffRq3NTo6d7JmrnS0N7Ohw1Nhrg+IY5Yf+ypTgCPIBxRK4BrZTv2c+VG6Y6ozuE
rMyvJCAMrDE3Gs3nNt50Nvif9TKCRXw9x3Whjr1YgCcPrY9nJzTh8NveJeVJQZYTsusZzetYR1Xb
bF2rROkoiEu1TvP+W6+Wm0AyJHN5fsms5F5IJyEAolshh8mYYz8w2w7qz3SelfdWs3laTl8f/lQf
xi0QkWD9CMMS+8C2TZOX8qswVrYyWdnGEWuozWWIWIcMA5daBZDQJAUtaF2pR5lGonSz13Dcxjml
/yWU6yA3RPHlu+Bd9pYaWx4JQg0PTOjZZ3E94kg8qQKFOGzVVE4e0SmudfeO6Bncno4v2R1D6nAt
vvYafwfzWc20sC4dJvderALYxc6H2AtM+g2rFrhv5sO9Pj81wQpBuX7n6pRqbipeWsLHwybhHHAx
itKXTvNXASPEn8uXlWyn7csEYfQBs1bw4v3ZKvgQm6Md/QdJ+6NPQKZxcn1jwH9GCpJKBTto/mje
wbPyj5/+lk7nAVkkVZr4FoGj182CYzWKMaZuSYGJPJ8a+vc97FoRBxPJ1yMJ+qVlO3W+w/YyLWDB
F1WosAtVL7iPt1x5MtoyRV/mm6nDxZuu3EJggMWwQTUiBTdBEvLnreEWcX7hv7nNq3ldHKWnJyPb
70ygky4npGzWKYkG+PoQnf7NhzJTlezLVvuZmrwwhQCf0/r2FaslOwmY8ke2b3dyNSiQ0in3z4mV
nsTubxYjMdzJD/KjxUuAGVFc1/3upseXJDBmTewKIz8oFVoK6PYUXIu17aNT7Yb9vRRr0nLxXWW5
MssG0gz/WC7GXY+A/metjtoYP3Lm7L1lXOZGj/dA4rPHBCNgzwxM6XtLxTALcCJL2Nc/PASW0/3e
C55sSnwSkRDqLPFLC6H24fH43qwQ8cKcjsEAX8Rb5fEdSw2EgtaAXaPLMCLzfh5tcIOtGwI0V6xW
9pDtvfji1Ql6yGaPEamdMhcgbGw0NxJ8F5N+oiVo6cul6pxdpHIgA/aEXIjmgv2wQ9rvuEdn55ae
PQUf49eaoXeKD55KkghExWpIbWSR7SJ6Bj8J1mZ8oemUwV7j0A12i/h8CThak/oBYrebkSgAjk1f
ET6p8d06HoFKR865YrWT/iPKXmMDCZjeCebw5O6LjE8s9TuyCCHzA2cCx6xOxBthS+KBVkQ5wIGh
mFWhYMjPDHmj2ax7i4gUkNNPS1tyx3YR78PaGJFQ1H52PSs8Hx9mmBw6JdGiLzBsvHrF188dhDGk
aTpdeGmBZx6xto1+ovYItDMDpnBEE030EtwudxT14Za64GC9KpygGOjJQUPGbHhVXdmKAnfQOoam
DklZ+k0Y0AG0Ofx/vN1zDLmXLOQEmRh6o1mUJNTxKd5f0Kl9l53i02mwDD6jG9Pc1DeH6Q+OkGXZ
QgCOLl/ynMCyqzJ5eUVFnLftN/vNieOIZsVN6ancr2Dqlhslhm4H81DqanHLYpGYQpxJX7FqtYZ0
O3TQheX2BOdOPB+QOe6NEBhofkG+vyWYwLYengT+e7wQxkAT7w7OsFxU2qDtO2MdfjT1nIIYO7wh
k6uWbD0z8oeC8I7BBXZF1EDUoYGvOW+yl1f6s85asDO344XDdwJkcidwSQLIfk5QQlKHcIyRVTKT
rJxno4IPgeIbI3g6cuiZPQdjaXlGKsoHYDhBNXbkkQ1tvtQ4/UDtn0SHtZFA6g1+ZWzPg42dZSff
i1uOP8PSvpMnBXjV48cnHVzdg1zDatT52c00oIPPJ8yD4y7LmPpX2gcLrsV8QWvM36JDrZfq7853
jpA5MmmKeheEz0VN6Br5VqdbZs83x2SyXiqVTjN/D9KxrDsZmeF111vAfb6Ls6GZ7hN7yYr9q2Hq
y3tUxZvXOh2+4/6V9lH55gKChYsThMCayqZRWVFYHa7feU6vs521ymhHMh9opic9IHOMCQuYWXv9
BUQY2d/FpLJd9nA1+TV+IX3eDPOkavffBGel+o5tfFG4+VdQNMNv9DIikn+8F25//wvimfy434m6
aB98NOn/0cSdgHWgGeDU2SAIbvifW/oxJ4RZ8EmorSkpqBvgoioOe4v99inaEllYEY5IXDFv+uWy
AfwNqXd1wSj1urnt90zzoncd1wV29vzJNRVVcG7kLE8OtpbVC+enkxEPftdHJolgI2QwFvvHf685
BTPiul2VXeTL41B7iMzQUbaYdZP4K2UBJ+gJhpVO43vhspDHrUlD1Cymy9iYtajq+jTDEOaRR3kl
8tIQrCrFGGz+VzShzYoXeGtA3TPttpscxjn1P40UD8UljK/5gsfgRZZjzEKIbRyqr28SMOWok7Ig
i/q4uqrGTZLQl68aHOPbAnDpxYZRzB5H8tw0bz72d5dWTwXODjbsokMuqNKKqdyoXYJhkQKJ1xfS
PKaZartvWIIWOFcyjmvuF+2052VV0/NEyHG42irSFOHuyE3Rbm9lVEZpdgXkmVtJBBGB137I6LB1
BOqgtpDESNIiuIJ2+mKpqCgLpejp721SsfSm/yBXdUxv96rwcmub6AfZ0u/BLyjYdIQIm3IntDyk
+xD/RUucRWO92w01m4kVRUBMxtXJB0HXPWlNVaSG27dMVhRm+GfhSUbWmTR+ee+f/61J/P0RGlut
8w3F5091HmTuf4ZuN/ZUNDyF8r7ynKeCGrR8XPtprWNwdO08eK47Nve6PkUunbEjsE3TaFr0mRyj
4hj6XN8GfCHDdGVhFg2szhmxDZxR6AlBlq77TSfnET7H+Hi67pqefYONY2JBW7DYfmQHzmEGEro4
Q4LmYyu4blFN1WS1B52zRTuURlIZ7KW55MfW7XiuUAOVmfH/yFWRoXoKFi00K1+EvzOVekox53bh
RI2e/OQv7pg7903xH1c2ls0xTNzk8iEndxuvabvbPYlyYtCGOCZCswKoppCRJwMf/3k14LzGvZur
ChN/JjpSTcardX8j5aJMtsBAP0x49J9B+wSp4tbE3X508PnPSkWrGmiikjYNNrwElJa9JAXI7xCs
5dsTCk5yeSEt3BTdm8QPhBsA41ivEV5GNVs5DCbaSd4TMUNt6nhrspgI6GwSxDdDYKMxkcPmD5F8
66OpMP82C/r/nBRjnpDqPvUcPBfj0cX3E7L8/ESJCW/SkQdJgFcgyBcTbSCETboUYURcKh8e0vkR
JlDLDaloLCwHpJF39AAFNqbmbz5kCh1EOt2qO08PHUdiYteX+cKKe1o+ibNCdm+S9OKTU7991coZ
xVFyin5Vw+cciP/rcv6J6BZGVS5yn8CHCjjpVDtm4dj8Q70D1Nf6WPT0ddw66iBBn8y79IARjEwy
QLcq7UWl3o+6p8dI9OocspOdyr0B5+TdW8CG1V9KIPd6Sy6TQTpn8cDf6aS/UnNhFLFkcdF4R3ga
ZCp680TXtR0KCy8ytcvF1gRNVZGv/F2cPSqBQ+rAhlNb7l2sjmk0Sfg1CFGoLhLVOwYNrnjGS0M8
h3mQ/2kGec1HA+AStGp495Uh1OX0/qg5SzVrL6WtL3VWEuzE9AucoJrktWZ5rmMWDhZeMYkoogFO
k2i/QnE+aDV9j4d7Ya6KkyKmOgpUarFo5pP4vcIhdQSxfO0VdJOcFrg+QyFEULB04SdS6eInLjlP
csyuPp5M8hFg/36eYpOtUN1MleTLINC1q6gsxRZp8cKnU+WIQ8bby+PS0kk1/Y4vpgL4rtl+Z68o
Q7M+HDslYmeM+i5H1D6/nUD0dOHiksiV6+SnRuiErWSlFrMRcUtYtcFx323rOPagXJOXVlNA/dnv
8TLa5I4MWjzYh0VuVinOUseX7pKXUXD9DwZR1s8KwBi+1dUzwM7/9E1HQrULG8w/Lqd7pE7u7CEf
9RuB8Lg3nfg6nSsvq6GvaXvGdQTiCGw5aQ4KlNWV/uVH1Sm3QQ486jkhm4RZLb1kkMcgChEYo7lV
hcwMPftMzq7jjj2iATbEGby28S8HcCQ53HWvVRgRzn2n94kgqik3MMgEt1/QBSk2ujDdIk2iEdMa
JOgu/kIC7m2YGBNgJ0LbVgMYSO1KyRiqNXxAXldxfUaYADS7SAaSGBIO3oRjI5waHMtn38gNKsna
FH4OKiwvYteJlUKUhRvTdYQ9g+bBIkYAbF/X9sQ/qUUDeeG8+72Wkshdaa1yCtInQB7XDeDNecCA
ZsXzGtgZNv8OtZ/F/PdtCvu+dDiTIg2tGSfPN2YsvtGIfX0wzOC7tLjcPIY+L5wuw8RbwbIPP18c
kMwi/5Rdb8dgytdR1a0CiNcyQ0swHeesYuSI6m2NTroCrwPI9jLwyuF1JcDuZKsKNZvNUzBIEXSt
v5JLwxMddp4+mvLvR91ybkNZBT/vhJMFanxPpkbrWaavHd9bDJipxTehxkQiricTj3wDhyuuokpa
v8LivEXN4K1SC7UfxSx8vJtwtF0csHFzxLv0Kg32PTyJBMrYeQU/S+s5V6e0x3C98ciNcGOALTsn
3txcKiWydrGw4gVoHXm9lE4NJA3PAjwr3IcGSkogomgum4EEQ/hBdNdcIpSmA+GCuTyY7BQyn3lA
Z3y94LGkrZ+PE+X6meNaskrA5qNnNY7E67IzVtU0zSFYSflHu16Suntl82Xzmf4oY+ZcoLP9jayl
DjHd3StA2+DvHginOrR9yN5utl1FyDmUTUOzITjy7JGxA1PqDeIOBbyZF1J+x5/HYobcoG0TmySA
bj2FG7VPMNAtiiR7T/ZUoY3+nZTI5+7fshGzF0JfsPdYf/PQ6/HL5G6jKOmdudm5J6o3NWI82ed+
POv600Nb16X3MgkYNheLiVzwYu/bQn3lgXZPwvh19g+0IBKtoUEEg+NmG71KVJn16L+ht82gn+F2
3iaTcHiqp5VoHQmeBfu6G4xI0u0UyBKL7sMmxRqc0t2IMijG7pwizCUSq/KNNwaPl66IGtKXugjq
IU4jbTWTeU1EJNNwRBF4qw0d5f0OGwfWSlzCImhDmSNVTokpD3wHUWBGyx9xMZKxtZGE5SdQsdEf
qq4ARPEyoL/Da1+evMVZCKx6AJ2es8qqXoNRcsTvsDtwcSs1rIz2rOgYQ1XtI2PfJ7v7Iju9XzkI
dh1t+UR8DW57CaJShf6DzMl7HbniM7JrCdZEPYhvRrU/VLZPA5TRUGgv4w0Wip+m+llonUMNPXVg
sMkj3OPA6/JaZa7O3oJFUvIPbGPJNSwO6DzC7iQXGgqoF6wDvJPEBbBQIcdFWTHsOCpYFLAexftD
N51KNWkYqx9lYvGpm8NU3rMnC5W4b6YlC0ry7iC6o9km56vRTNi4kg8u++fBSLFpvUqE+F51BSFy
ijvYyjcQv5XOwRRi5cnItUksWlTpsFMz5G5ZUTr25faZZ0ouBY3LBt+GdXuscccqu5zOHxXpqafR
fl758L0X+UCS4UBXPmFyJB2dKwbSevZGYTKOwleXcDlOh/C3OdSRv4QBbgGhY4vy4PMuC6eRxebX
Xmjm/uHo6eohHBgjKl8p1Gq5vtLxFoIBjTQyt5ShEqrZkruaeohHwfX/JJjZPZU5uuKenKdvnZKX
tDpAVx+bmo6acLOcSNGu/27HChVfjNULGa847iXH8G/zyMHwPmPP0GPp92YQa6pndbapJQTcP+89
AgqiDt1nJKixCfXjbTrDPgEY/cJNHgA+GP9ytxVyr7MwWxgB1Fah6NLw+vSk7kcdz6ngQpSRP8dt
zSB/E5Vmsy6Nv936EO8vd48IqrBUImJo8h7DCFI/joXtfqc2xRDVHSsxVGfC4+D2OioXd+bTmrPU
5ajbwvZXPgU6G4Xscuk8Pp/fAmz320T0NsgfhgcOedQLo38klK8cFTL9zPI2xAUKfA0KpRfHxg0d
zxiqekcsAFNPX84Y+w37AHHYRFCsGmxo4qR+f3yWs+0uK4XhHWitXUM0oJiJK0Av/F1YxxhBEYKr
5bHtGUNVBIMpirx5Nt6MNTMbXuaBqS8RmkVVtNk3TkGyaMH+njaQJTMWVxBl9TWUU+FvD3Bts959
FwtPn5TEWWcJ3iMXa6OxeaewCqKbZokrn2i5DuM3Re9tdNPkqIZS1Sr6GAR8dP2ym25tJI1woWW7
KqYslKotL+T9o17mEJIHC1N5dV/9ia9Iqz6k1LRpyFPEcXoV8hioH0TFYNtzric6/AssIKvhLPph
t3/zRgWeGpsruB6YtJFRw/PYvrKtVVEW9gE7QtY8lwBSrrNFapfIFm+S+oBCFOpApAmmUFNd6esi
a7hFKQQzJPkrHMBfq2f9j/h7A+J6hWlHP48hxUDK1/vcl0dWgbWDr7iycq8vrUS3/BOeA3I+fV/8
ll/T+LqUs/FE5CNETJXRc+m0/IO6hQjUI60azRcrBDJsKC5FOgRwBbiZmSdBW+YKwD3s3nrB7Q/e
A1Io1ilYEUd+/pshsVOb2KrnqOuPqoYfa4yGxB2K2QN11pe58xKZve/YHJ9D6gj34XoAumr0n/Yn
mA+gP3Az05atIKuVp6mZQvHA+JLmqBEvrP+kJ6Pt6GoMZvF+HpAE7bVXFSsmFf6DkBwy+Ar+L8Jz
GN8g6oc6Y1xBOzeX88kRbRX1qQr3GNho0kSNItJWzH8ie3WYHkxEEXK7p8EBQAESJiGUpOdekyWg
OVF0jxfGGwsofk4AOjrCEeNdrhLuXg/FHkL9GGFlX9EWKYxpLu4S5DaQxLXO/B9UoFzPTmbU7Xah
3gn9lT87BeAFmY2j3lomoTuLrYDudkjITM8odxcxLnnLYuS+1e7ZwEQxD558qKbrJKhF0AAxproS
UE5A6iu+/pcVnf17Hb+lbyZ10saM1m4a5dkvmURWtd6tXm7uEPoWUqWjVIziaATAVyjQx3+eKJnL
AwKBRkRrsGWyIr5Or1iuBfHXRU0P2+FCDycU5SX8G77qIMeC3M86vki2RJXgGtsDw90lQlbG5Rht
ETdtKAf1Dk8u4cSlrekYN8/zYLejU6WrA4GQ/fXxplBqK7ZC2LuAJB9KgGQ7l1afzK0/z3TjKdAA
Y40ejXTdZK7Zpks1FDpFiQU4FS5EGctIaKpSupASxChal4EEHLNb8Z2P/rCbKKTY6fcTNzEplHhc
Tfj5TdwejvxQ4l+fnnI+TNZWRRctHY96CHUHJNVCC6UlaTUhJrTXd3qe/U1fXE44UkKr79R4UFS9
fVeWb+8rzDpPuOqwfDRPlmK6fL9tEYUd9u4heYS9wcxa4zI7e36Zb1e90FZ9cdLhv3YA9J6Bmhn5
7eVfXKzu85xwheYtFvDnKNfOL7xglmN+BvXr2WCzB77mbekDqj8YTBZiSbFCK9GJfZx1kd+vDn1I
+yPiXdXRxQoZXq3qr7f2dchippVHbXmuPGLy9KGWkHeIpHEo3mONgsPVA3N4b/GYXyH2nsyZt3S3
D2BvADuDEn5LBr95HL44xZU2KDXXvPVUtBU6NSZ2VLyYDVHfAuDJpjNrovodOFsn2QCQRcxYXpPu
niUcBi2yb5zChVstEtJONbh2FMD0bO4EHSQ+SQ88vxZxlO0u1GRlEzr8srLOjK2tJ0xEOcKLvf/+
WrX/XI30SxvRKba7PePS76Ms9OQWqEqVH3YYxPrGHt6+d5YkrUI6TPJ7d+8cvAkde8/TNZ6Zunmz
Oy9lf1BfaAzxfqiqYsJlJ8+SHkVQbj/7kL/oNQ7jl2iRAewQKyfqiPT5bjSYzfIlWdcjMBqxLsd3
1Qxv9n9G5H9nQrgUIjgyNjr4CdVo9kw7MMz2LYSh2qejm4pIJUkbEwCfZ5lzuLYgu5ZIUTn71ZqQ
supMLQsADRD+NHKbLnw/dAmQXONOi3GuYANmnhGwKXyIMCvTIRdpzoy5SabYy5pBZYpNNduOiSlo
r21WjCPE2hUS8J+UewV1IYtEmzLXe6iX/AvppZBDuzQ9ZU36bo8AIHRX4TrkG3sFE7FNcxDB8dhN
9XCV/kqyLM3qYtdAQRe5DHoXCRCiKVqY2oatT8pDAbwiAcwJO55PnV9m0TBJ/v5OIDqfl97Fmig5
KuMj6XQ53VZU12eyFQqX6AYFrLG+arJA+c7arMDG33TZY4zuFlCcv+TXyHx8KvwhBbQdzkpB3Uzj
71uzC7wLvEvQ7vVZM/onSGeNEq0dFqzMX+ku9uouZ1YBoxxp3Ud+175GR+LQL5o06WJ4vS6O7cC0
W2Sm+cP6F3RTlWflgGijCZbNs7wOf7Ykye1XZEb9PGkYk5eAKXsz4JVmhl9CE91PvL73a4yS+fLw
Xh1KLcMgOYGowm/KoVk2b7uG5JiZipFoqPjQySHkrsikNJQZf2Zqma/6eGPyG5cJl0iMsOkhNPrl
8vTQ4W8TvFXx0XRaityQiibF790fY5F5covT7Khu6K8DA9UG7bTqksVVWbbTDhpsEisTKQdtUVpT
ZjMGilaEpFJk6Yf6xGxu2+HG0lVEeHLslLvJQJu3fkcB3XK+mdNNuiDvxhGALwpLFo0zA7RftvFW
2igaiL+x6UF5Zg78KS3dWDCvuxyDJ689y3kKYsupIUz0RyAaZ/E+bhZbQbItj8VR0SEQuBChWOEp
AbZGxsxqy80wx5GdDcKc5mE3VWjrPXhRRJ0tjit4ZOw4J8boyPHCX8my2AeMwo6u0r4j4KpcmowV
js/Ap3wFT5NbhV9QXE5CqDrQ01C6UJJAPPig3Sw3ot/757jp17Jjmg63+BSRhMhVrOxvbTof+acG
JsonfRC25hwgNLIILMHkorsFv8cFKeCdyaumF+wyFOLsQFZytGowKtQkRka2CZs67ytNDt8r3n6T
Uj9Fu8MLjdRFGuKllvWTQwCcfZpMVG0MYRz8zpwZreU221d4LO4NJ44RBpfwAVkoKfVu5loxx+gQ
nEB5FvOE9t+It4XmYfH7k1joi3qjN81JsQNIXv0jvlhbaF5BaR8Qpr9NZSwD2/OaKwX9X8LgTyGi
VMfvs4hhB1BO7G0j++J6om5HyUrWYFnv1IL/T5MySU4b4V8wbmoTpKI6/Qh2dRu2bdxviwufHxHu
d3dm2dDt7q8SrbG3Ord+wVaTUTNSAw/ELs+FlHTU56ONKgsws2YWh/cuMtoRg1kXeFXhb+gAgBKS
Sll0hX4g9aGjnm6CqDArh4FRYPNy/YuiQ0FSkAbX+/aD6imAJEZZUVD3a2EQm2pkA+rBKguu3L5+
2DsyBGXiMvQmJplBoc6lG16MmcJd/jcOdAbRpF0z93Cp5YVLOgJ5Gec+t/2+fZrv649GlrMipySW
+b4YlCMysl9UMLb8CLWFoIcDxQL8dQ9Z3/45zyMteofuSl0vong81/GyVItQcFXQd+yK20E/7d0D
Y9jLDgPr67yW7xHX9wRDa6uVOboQYr1BpZMgnfsFZ/LEYxH0XufQWpECvSNY8qXutGqhzg03tqQZ
9RxctK3ZapQDNcuuZOv3dJnDMlXCd0o/CbZ8wRl7ULnivHmNH0iRpbGBO7bAxr17pPgOn+rrDaKp
dFYkEr09+zclVkp+3fM/kBV+uvBFZf4U4Srmcsz8/doNP2BUu6B9EZwPcV4hUHi03nJQAVSXTl0J
UymZojlsXkHVXkUBuQJNZLwT2EeU4H1gUO1NQRUvIkW9vx1H9neotjqoziD3x1s6BxEr68tCSFBW
xBCHpf89u/oaEvY+NXnONnnHZx+uO155R9Kw+wy74Q4xruNytlqzEGn0x0jwKJMXvjKbs2WBrsPi
hnddH+u35Bv+imipfjHCCenxQCJHeu0JyGuoiucuqelsjA2um8DWC1M7HL2vaW+rZWlBB0M9pQNY
GIOqqKMFcq+Aolj7UKnE3tsgkndObccnNm+BxU/aEFOaewxhwZ8ZRSTvYvnfVuUSW5b5AyQccDeK
nzsCFnc4fod67wQqD79s+zIiFUKWTSr21Uw1U/yG2tScME+zO6elzWbkThW+aL/uswb7V2iZVDv8
5mHbHlAJ3li5qKkVMmTo03oB4p7BZOPP0ZXyuEgauEooeMLfOtl5CsgjWLXygUDYuWS8bfTLytCp
yravucCuDt1pCYpvQdHmhVCjthlwwG2nNswFKE+HzUMXmlAZjVT4C5D69+Q7HUL5fuWTaJb7M7E4
i5g0gssNjGJCq1R9bC8RyFTfF6NjDYV/nMIA4NC84ENDVgqN41SLSzv1UDjd17q9MPJ4IxG/n7JH
Pf8bdYQg+/PEPbKLtPeOTHWdvrH8UIbMp2a12sjd7glMjF0HhIKgmsROXouM3GlE3dqpYH3o2b01
2nHxIwOTFUZulA356gW/Cy28I0NwXQcOoWhP9VF5TxXkDWwP/U5jup0LuaNnRMvApo6MgDQmL3/x
RtfauNYy7zpnV4RT/dD0laWcKVVCdPBjIuUusNSRAJB/3JzvqShyIKbk/uY82MZOF69Tvbei/O9R
ZgoyKrbkEC0yKHWtGkflnn5qtdwZnEHsHPUGEI0vyoBrhmUJ8WmZw0RGrCyTv9ehVrEXq7KQ37dO
Kf0E8XiXYI9WcwxFZGicNSmfuLccTCySnf1wvzamaZSbLefUYRLn1Kcz8BR+DkCukKK3InVH+nCh
HX/mbKqZ44XualyW08OImUl/Qnbi8pipuGlo11QNFcqOxuj0UuNDsngaGmSUj1vRV0Z01wS/lwa+
GPCinqb9NFQmy4M7RdPNwLCmD9fLkUBMJPtMAMOiECOKpiu/Ejp0JC0AXvU+qEj0Ksqqjt2pYCRI
A1ieWbzqwq5cPffPD/tL44q2uiESQAaIX/LIE7ZDpsSubFH3FpKSzKAc6bS4/2xTFyO2Tc5CXu88
6stzV6OsR8zJKyxvz6wNfBf5eEoHpvZmq9/JwF6sb+hUcv7nlvOtuiXN6pyLD33pk3RUYM9it1Z2
E1u2EOjkhTSfG3RBUPx4rhGE8nazfR+bMhIif28pvZRPhCAcW1Gf+PCNIttzz+EbeE/KeKrW5xT6
qXag45PrHfJWPN48ewf4Iofh2EWnkm48gKLPyzfT2+jDzGrS81zLJ8WP2li+/KZsSXGy0rPgPVG1
U6U8Sj+nuwwtTxUUzqiFjsHJ3LlEF5u+QmL5G2pmj+CnCPQghon/z4GanNN4D6AUP+IZ7fxGHRJe
V5fcs6oWvui9jWDYtvxW7L2aClRK/6jKNZ1dOiD9uXOX1Gt3Jytv9r9ooGYYIzhRDjhDzRTYJy3o
WTvwFDho+rjF41DR6FLA4wXT4kJhJR/IgV381QoZoDCjBAYaF0AewSFs4O81ra0wUZN3wuOEK78G
O3yltomXMQqaP1Zv6Ih9b6ngaREPlOkstErR2eTcj0/qp8j3UyoFOiA/YUVIU2+CW1G86SGx5d9x
WKmMqZG+42TMd/MTWG0i8ADqEhv3gXprxrg8rH2wGGbcWPvIR2f8J0ELqXQ1w2+uDOh/xvmpklE1
ds2zvUVVpdQQ51dPv7ucQdUSgPoll8wT+dEjyy224dDWD5nt4JxqZco/YLkrV9AZjBYj+bFe6g6R
ACULLWoaKkTlU/sUA6xHwZIKAZ2R3RJXAjXFLgp1h//DVhiKFlFSVNPp8mIAwo+AdjX44EkeSzPz
4SyTv6uWhAWmtgUAA5w4cffTgcmw7d2uGDBBhnRXNwajIADap0yeejZVN3GIC7dkiq9bkwiiMY3o
AT7B2hUxLkAu6YZiOqhftufpv9NTPSkwGtXLj8n9cOiQYAyUI8LgXz2tNsc0b/kcy9aA1ftcYbfN
/3JJOPYm2ThDoFoQOOv6dQrcI3XDOX2h54d4s+kXPEelKiQr89Ev8Oxem5P82jktNltlYldTrrCH
k79Irj3Z5uvWgKuCoEYtaRXgh77DyA6e1CBrsOviacFfFgtL0XTGa282ujqpzgYV2qeL6/Y03SMg
X8SOJq8ivvzf20UIIS9Tfr/mEos1mwjjt7vzSIIOLn0UnVj0Z1kHmdptLCNSkunEfaxMKRRCFZED
Bfh+UfP9rBCdXsILQ6i/ZSNYlmqXGhgmUxQ6Pf6sv4nyht0aOCUIeTjoeqA2oYyqoSOP/sqKiyGh
fXy6iLjOfi3d/cTDkMY9Oh6o5YTU1UDjOq374XicbkvgjHT1jcI2wy5H6JAdvFNouSXjgK+FQGdD
25xDT+vesOn1R96W62VMnK3dKjNPbJJ07iYr34B2p60sJZtBSbxTeMnv+EgBtpUOlE0ejzmN9jin
Wl9uUNn8On2yhrWxiIq91O1QhbPJnz8XCpxzNvuXaf3CitGHX3j3NeDOt1JBRiwz2Jex7ksoHrqk
oLXnXzbgM2flEbub2tyNcczololaWDvR0EG1bCXHiPh3TFTU97ACym1bwqBymv1o8Jmi4tXnFCvd
OLL91kwe3aKa9D+UaXfh8S547rZ+EmIIzJBKwTpZ77pLBr3JOJSQUSNdGUQ2/JAgeF0dIBRtkaT0
KykK+lnfQUYHGDBeoLpf0PiRWrfH7Iw4B1hNp/FXOdPbIhT6j/gZtunIuTE+1GOXukcGipODZfBn
/7jcghWFA4gtqiIwba2RQsbg3VAOCCGbfLlAF6WRAIYu5f9Fyk/8FASsR5rgKiQdOhgLOa062WHH
akGOC51T1qF9dmSPcRG2KzzOLL3HxyzW+mY84iNumLqjgCxb1fsk9xGnnEJPnSOKLLvVw8goHcTf
lAU0eNlFMHVq8YBpm4Ym54q5F+iV00f9JVNVAfZNQTyWzR9hH9s0d5Tgc1kUnLKSwmQygCRbGnZy
rTdcgcI9+80vDPZTM7oZ9+LFyQqpKB4q8SIJHQS7T6MmOpFx4sIPGH3MmiGofNX4ykX93GUGlltA
42rW/zLLleH1kFREE3uFEWQqLTYBBDg595oqqCoI4jCeGZHxns9uhVh/1WLnnh1aMZk3VkDA8ZZN
nLoTzYgYswBSN2FlvXGW7uEgr1lySWG9M0KhV5vzzE1EW1ALrwzlP3pUWhn0GFnr82rL0+EE7VOB
c0dSQOYsYxmBr8J9uNgV5l6PpJ7AQjy8KfIsyM14Yq2Ts4Vp8YGJtfAb7T11xN3qCW4xo3GANR+7
e/9mmdoyL/8k+im2rUyTt5OWz8C8hXKy2LU1ZP8I7uNFkyYBpGA55y4kyhTerxqjKk90SCgTIEJM
/esemZSIdg5AtFDtzjnn+S7QvYnw5Uw1mIozHK4fXuuqYwKH0AOD8X/rZWcNqiQ88bRQGrDQj1V9
ZnlKUCc+KIV3XymzQ7JBvr9yvrFS95JeQLDhtc3f7JqIwIQAh8r5PEyQofOwZrHYu5aeiodY0evG
pCu4BaZgWjRLtNHkY0F9YhKEFXWbpVMJdzYSQ2ku0WVv2g4jep0Tm2zuV4owHitlVtpPDoVBaqAv
gCz0IdLxe9MP3g5ue/Aa505GvT9mBE340LDGGSSAczDsMKud+TSFqkxvQWm+0czNSLssXyQfUYm5
9XKWzUtl6puhz6NtGUqxv98ja3u0TE9OY6umWY49Dv8QytwSpCAKwyDaAZAVvy8+KBHR3WEEoy+N
NUJN9LNZXl70LB+MCdJ9+3+AFxA7U9rVvgx+grVIdztXKbxcqs1DcDfRFkfAxnV/jPAVckaja6Z2
dsbWSejn3k5Da8REC6L1XLTgeQ0R5QwMhYUtMuWEt+ZowGS6dhFCVGJQ6Wu9gJyF5s3Puf5Qplox
GNZzUESzDIJ5QVuqE7KT2cR8lNmHQhPsqLHbHgYrW5iF0ytn46JBNVybL1DlUssy9/CkDu+v3Tyi
fzlzV/H6W9tEWooAigb+yg4/wqAOxYlffGqzzJVjdMUGi5zWCTvf4IyBQ0hAroxlPMzyWszDWahb
ODrmw68xZm84vmdgL/4e8HX4zq00OMMECFPvoKjXPmfHPwPrdL3Nrheb3Bkj+lT72b/K4cDqqKOV
roCSzn00SIhUT+z4cUbMow4Bc+aoaRnj2KKdSSFt+jO1OxJkPyGd4Spqzfud1D8Q9+E+tbYqD7QP
3mx5J59Qxvn7o5y6vmCiN7wGMjDNWqey3jYUOST9NJY1+EyTcEoeDVtb0As30JdDjbKYfSZ2eKLP
Jh4zy9LcMXgD5DEQSGUeToVWNKvlF2Fapmu5OjOx2W/Snd/gzMy2AxlIsVgPPf7J2n92MDvk6xYE
UNzy6QGafHh+rY9NNv5qgk6s9bdIiDNDLQdosf6NMsQs9kkVLYcR58H6dLD+mN9DviGtLzZwXUS5
NMpZq/IC/x9gGbKLHqQQfqohI+RlJo0qlzJYDkVNwSth+hGo477t7aziaUzr0mKt+f4JP5lFIWS8
tCN25NJ020ReQALYaarm5qhcZ2mHc08Vf+d5CT+k+GoemR8xAgkAsBuGivweidIvd90RpFmpkmV9
28jB1LcLuQcUdt7rhnPRwoN1AWqgTeG9SQuYNBCTkuJkBpzMn9+hUHyEVJihfiA4ZOw8pBLAycDX
lrjB4ZjeDW4KnYIY0568dx4fgEZuEP3VqeQdIuAUNwdXDFxgU6Xw9Ba5fh5EQRD1SHywJDe9414k
bxBNvyqeiWL5kHWZFgEf0zaEjkiGTR+ZYnpeF339tdLFfizbPxhkSsIrPHXvn/P2Hz+QrGZy939b
RkToQG2RLh+R3n20IEfwZ96JNFytOOQjoPtajYHjikdXjHPYsUtmLhUQWDpzEqG8pKJn4FpMioKH
SbKaaLkfzLbjXObAmfvIt3YTihTxLbIBdQECF3gpD0/k2PH8hDGfAP0nkCEo9zR3ScizmVIHivdR
SkRme9aPXaYkkc3aZoPElf0qpJsYJN5QcgQJi2XoxL5koOu0KJbSu5HUITxfh3tCEAIl6AoAM3Hq
dYHSKWcB7+DjG/GFLy3c+9az510ks2F27/5ZnOihp3Mz68qH5jlW7kzHOQVl8C1305wA9t9f7jCw
5w9INB8M3uCetTrQr8nLFzi5NYUE69Wj7/YmiPnmgxYmTesg0HOLdjIPxRX7jHuPEhd0Y9/esImI
I2LEgwdgK0QWsqJqiUf7yEbBt5tkDWRmL/6D4j3nFKLrRd2bEXRyMilrSRUgQs6zCoUheXFM462U
bByvoXNa7hMtgeFoiPrJySBV/u65fCabYpRRNslTrlhCezHZf386gE7xaZGTYJvKEcParmZ/DG7I
8ADkuP4bxmNQHa4jaDpfubb2pbpYDcOHjBJy7YsR4jTrWmfuGu2oYIQJu9ei5duCTK6bRtdZhJS5
geI0LsxJ5hl8tdfV8cwpBA+HdIfDmWgB+y3HpYEWuf8CfKUIddL59qYiou+liPZ7BVrJEC+3qFtU
Ng8GVTMWEpFcU08JdLMkhFpbY/E/RafKKjRX8RShOUssr3q5ATLAqcT6PS8LYXG2TApkdnfotKVD
uXnKKcPaWZkHGLtd6pjYu0IfsC6RzMACNdwpSPWfY1hDgPbDqPVrGeX6moMRqh+n+sgHpJ0iFjzI
i/Zc0SR0etgwi98PalsgqB4KNb1MK5Oy7a6DhWR7McHRvReo/OgA4I3gykx37pMt1Itb0oFbTsjN
Xp3AUt1bvmNshmVvvpdR2HZhdhWfSK3EPg15q6TXtvK/El0QdU+CNJIkOEM9lTZ7HVy+DuqCk4t/
Wm3pPB23MotNsIlfu9iggIN4iW3sYlERCkH/5VM+A/wk/mnt557nQ9YI39CmXwY6wvuz+ZvQi5ej
UjNkR30V8bUf5zyNFvFxel6CNW60i24LBsDdCSdoIjfoE7fLXMjbvJOMx2BN3geOLXZELrQJOT+1
uNVwPFIXfrRNqtQQ/XwWjyqY6JfJYw2ejuc0av5KoCcvClpC36Bxj91RDsYy7bpcyOz7LrwKE8SZ
FRgifvHI3H6r/j1dakDw/0JMgul8uFY9Ywaldr4wSgOz8G4/WdJHZ9cb+RvQF3aFapjZ4T+Ar0q+
H7CMx0/iKF7dYQEV7dLfp398F17WUzw/v1orvNg36NZRYaeIt8wPcBKPXhOoe+Ielky5yeWhH2MW
J+xCRozltOpd4/ZTmTT/cgL+V6J61rLglLFdJVv/o6rPC8I8LMAWM3SOhU1PhZ3W8FpcXE8kSzXp
ijyJj6bTYcp5oXGI+nDAAYSUGX+h1PIYds7gx1a69QYnEh+0K8EyiwcBfJiNzgZU6aNDjPDjXk7q
nz8ouCtl8LYBxK74JzI8lv+C+xhE9uWYSOaTyYeMkxny5O//vPKx4hjv7SUF11RnYlEErP4HrtCe
WzC4Q/6QNYcsgbBn6c/3at0myxqkcmYBL8vKnRBjk8njOAJQ9Fk7aiUJeXsCvTqWtoDTmCU8t+an
ClTTNxPSMty0edEodY7L9o6fEcIZaNGBY80sLoq61OmUWJkG7VRQN60KHuMNHWykOWxdmG/QGWHv
YBxxx+dDonzpFqWFUHzbzMfe+X25OxCqY0ag13ZfNMXicelpn5UtD+1iJVp2SVPRsXVpOFqZzbW+
jKpIQZKgxcMMfb2YUnqW/KTT9ZJySKQhpNiCe2jM+VSIuyqdXaGmkVpiXDL5qErM2VMVQGCpGIYC
kslhhLWKXBZ7Q224N2eA2hZm83QlFTOpQ84WAxHpTLVyGGFudW8NJ3Kr9HjExHhdDOvHIH3P9Mmu
ZTyaceqYbaPd3pVo7MdCYZUEjmRns1rPSNq214V6DOQH44BD2QaCqj9TMVwEEc80K3oeU1lpiqjh
08IC5ZwfCfRzesy61hFigytwWfmtjBgjNqBnE62BowyT18TKw612muP/vJjfrAM3qZcOxRob9P7b
QmgG6VH5LLM99njM55btPy9UEeQEch4NC0FWAF8Mvm8alGJ8ROkw+w5Rrzr52/FncwhXzceilYvi
9PYv9+F1Zd2TkIPKIVY9pZTEFD08P6SgBqK44k8ZZZKTYhvLs6FMbeAPaNt4Kq3Ix2aojCYBu49i
WA1F3TY/8IGHgDdxK9kxoBY6Od7Mgy/aWET/XPE5TF65ujCt2vd/yIEKXkcXLwNwwCImnTPjuxeF
WZcHHaixsCTH9ykHqQmA/s6VVYDWXayGmkWAWYs5rDXaV3eEEuvaI0V/r+mpL0OCUKyC866wwz7O
KTUxyxZLI+k/j/WMn5hATm8p35MUC6x2WQbmW8xnkNMrsOPInMq5NVlokxDYqBp4mfHN8R2K3kQu
73Pp+dzhSWWR/haQNQrths6VRIvyNt3K43EMOIm9T4KjiAt7vefNzbKOpDJwH+3QG+/Tk3bidyWC
AnhqmZhw8OTVf0Jj/LVm95dQ/pty5P+tRvscDiZ3V8/6xL5J+yGDR2dNc4xGpmGF528pwawxbz5n
iY9t0q6NL4jPm8h0GqIqy6VWCcUOFiPjYniXhPOXb5dNTw28UAzFlIfK8kXWhdhCq39xQfbqcnyb
QG6tmvIRcq8Yqp6GEMOEbS4L01Gi+aEoNa1+i56VIP9ESxXd4Fw6EwSlH5+PgqN7sYaJKtpPPPGn
7UsTWc6pQfGTRL2EWHodoxfTx3EJ6l2yyTF8TChoPopaSBEaPl4LvNl3EH8N1L7TGS9Nyk4lTVjG
zAKfUB+gJepLpKX/DA/Uz0Xsr7ZpHUi9OsLVnhOlQWibfZ14oOZ/dIXocgk4B6v5FB18V48nxQ7p
3ZyY/qCVDbRsbtjoJcG03Cm14Q8CvHVcGr9MIZ4N/vyPUyHtCExyrP8v0UJ6XyVDU0zkVwGeQCuF
JkgixNGoWigmpWEjx2v/OrLxqZX1ZFb3pvBCbSGJ2dV7DLY4kVHrfNmrn6Vep2nYAo1LwEKhg0Yv
bCci2oOX3keqKEf60ZNMORLiUv+Opx5Tjo4wBqCPYU1BrNiBy69kfnfGS6HQUS0B08kbvi8R/3LJ
jarFbN/F+qBciq204bw+bPNprzHLYTq7M/EtYEM3GTYxDLejlAKL9ptXbkLs6tryC2cJLPV6f2vO
JwLrxiHY2AybQTookfdcGqOOiSVMSSuXAYUJJrb0h/B1Qa9UxGfJCdqDFwFc5YpMdW9UGZw02sL9
2Yjezqv19VePpeEwbeui5YJoUPzpr/Dn7tFncufjQdC1iCB36DAGOQM+fF1PW6koz5mzbUaycsKl
yCP9ctaMDsPKZ+52dC1KzAAskLc/l8l7x9QEonwIy3qU9/bU/LkfIeS+TMOxzAz/ar9LYznuKQy3
NFxgdbmESNUoNAZsT7rLiVLfzAAv/G97kcZmemj1ivUPFHM+xF4nYMdsVztCapjUFOGoC0a2/UIB
Fx9SndmOGotEHyKXTkcmIm9G2Ft1H4WHi56MombNJBWqlUClvRnZZx7F8zjxA/1JVdDxQ0idJhtV
7KENzLBfaFU6Fv7JZ6NC1XSoQmErneeJWx93WnNfMzaEOKOtN2PJdlgig5zTVVHatRv15xSyU3Cs
TkphaxdmgZBzGaxno/IZOJeOB8hTGB0HF34uHWvhbsZJb4w6J2B5BOyQr8kS7ftj6Ebf/sB4ZD1J
aatPAKk15Q1kL7vjHTQ2q/8uC+2BlgWG/g+9pELV3MXjwL9HUdE2C+bTnZ2Jf3fej2+PnzLas8W6
A9BsQyjvSGRWTqqAPMv9UsxsQhcxQNguTrEBEaWd9JS2/chb/X8to9I6WDFThsxZdJotq1ims753
INM1iHXP+RiB72AWzeFHB1k8Tjp3qdFTSRSodt43Mlfy+fAe96rXq7TfrWBIPaI3vHSAgXWmUj9E
ctHPwa+D6tiOZ22siwgx0OoQ93D4aEe6KQpdS/27zFZMojU/Y+1eQjpSXiP06RT/s41T4uqgUBeH
e+EPNmo8Yod1fz5MgYkjUxJ0Zcd7sTCQmgQkywGgHHyrMloPfKYq44butI6+Nr08SBtSR9C2oZud
85OOOh8GROMPGtaOsqcrf8Q/fe3KNF4vz3iC8ShwVD+Okx1ImmXEsefwuOrZjUQu6Y9J07qfirF9
ZTMw3mdKDtTRHbbo/DlXnDYhykpvNQyA7bZKvfb9SJjuF0/uZW7xw6/E6yceWp1qtomt+osZNf6k
HkK99FRnrk0WGSqEJT1HqmwFd7owvK8CB6jSg8vWM07pHIglr9uJ/gC2cyq0k0D9UyABZmPzVPno
qkMCqaX7S0EY5d28zN1SmU7n09v20o5wdUymQ/kIwUfeRoWplwidVyzzsE6EgUoGo2mru7ZjMJSG
GPdQpszSW8z59sazu+6CCSWD52MvPLFNxrsKyw73Kq5qN9Kqwn+4rW9AklzbDB+4mCLiuA9h+9Gl
lrZ3a5Hi2K6VZywNbDd+O81YSdw8ArSh+UKzGy3r4clHjPgrd1ct5rt/cymUgTm54jhx27dxudEz
LCsg/FaklzbeYVqPeYK2IwLqzDaGw+xzglx/eF/a9/oaKKJFEYW3RFflUNVBuhXB5JIva6wfVNBJ
sW4hDWGBqpzKcDuzw6gZI3DOfuwfXKGccDQyMGPBKFprialjKLhaA6oUvxM2ORK9DfKljceJU+bU
id/0ZR6/sZJwnU5NmDvDtwK4abMNAzoUS6VjgRPIBnf2AH2RwfKNFo3G3tM25GSpIqrcwNjIFFrD
6V7bJDAzTORppzA3LMHuLl1/9uaiXdXyqvEfgKueqJbpZccPpfyWK1qA1DmX+X5aV++ppqTR7eDL
zGp5IeSap+4BC2XRSPk55s5cE1mEMne/rdme1xWYs5JYbkyJ6uuGE/I914/Uz1B3YLfYIBqy57OB
tigykjg/YHm5Z9Wj2No0daEd83Nx93Nu5To23u2e7Jba/eR3GB0+2Dkciy294Q6nUoj2Z+nMSCJ0
+Td0U1ayUQzeevqdQnjR/AvSVQhhE/WatqgaNYa+zsr/qKln7ca+Bz9l+Y+SO9ANTbYuxnH/8xx0
Jk3s6vA3xuX9cvpR6K0Tm+xx9ivRKewIOZ4seZZKoz0YljhCbyqiqbLMqwkQIRlkqqMYP2t7BzzZ
MoeDr8cXrtP58WeN2soVtCbWDUWlWRvNKfXPZ7QYIRmY8fYmui3VvposMDGqqlfeZrUZnlMCegdi
vrrKmYONPu8o15lbXNDd+IkvPKgL5Z5R0QIAKYOMFkzAOZBH2M8OROLmGGXJ1+SpSPlBFUi2dO8z
c/apD9Q5J2i1aMYhIqFhbPUoacYhogKkhtzEqo1umQQWtUG4lkbf8HpfXoZGwqlGrhbJ+9ze98Sj
gH9xmKibDF/nNY/nkkQcw52XZgsaPfqANuBsJJ2C+yFGpofcY5yYq3Cy3zh0E9ZHM2anP8rSDUvh
K9s4iI5PG0jZMkYp58DusdPfGgWFtN63xKsSuTXl97z7HOY2iBJ2CgXD7n7jjvgtv9veSWIhlq+M
a2yaGe5TrLcPfXw/nzTYb1/mNhJcScKwl3vfyXRNi0Z2cwZIcbe7wCykONk6y3epcY5j3CW3dqHs
T0bA4OP97vsiLWmYbj7rF9dKDgJPEMf8GoLBUXUzsGjrUboqcaQ8gNVxtdRLMSrLK+Wu3S+pGKun
4UZu25BsZzVWhItiGBGc7HyHtY34jd0PdY34D4OajxCQiEdW1Lx8FrojLfjikGrVtbvU7r3WWLmH
neM7i3yFkxohUPiOpiAFXRu8xIwHUs+2bOUTJn2w+a0TcUbMiodVQrCo/UF7yqpC8/bYyxF2z3qT
Q7jl3/jqTmMJOEIbQwYYpOADPG1vr43YeVDKmGU8CTGhWFuhxkGfM9S05BcojHiyEQ3fn2FC9oFR
18FwCrmW4R69BmIY4ziBMj1QSJg3TY5d+f8DJh26IaXQh8fhIfm37MaPE3Xhzzbea+qs9dSjLyWT
3DDSwveHD2cZ2Do4OWc8Taha3qSduMdAvU8/K+D0ZxfYmY97JV3gPn93fkP+Ot6Q/rmWG+r1yZbA
lnS7EwghxjBhsIKl0TWAyEc9k0K8jSb19IdOmbJKt7IH8mvpDZ/Ktzj1RKruOnlZ3osTB3tEaR4/
1oTTbOMuyRz4bmitZkOGTweb15SLFIvTQPR4xzrALnzJ0DtzJcNA0pji/ujKwnba3WGZiPxxvA//
b1H2PSWR961DraW2AHjCibWayKcal4xuJKgD8r7iqb1f7bD++1Oal4Q7bIaz5kt4Pf2f5tPv+7TE
m92I6lGOWi+v4is/DUk5AayOHl4r7iLoB/h4jucu+YpzLh7PEOS+Zl5SkFWDVWcNDcc3Du+BUi1A
RNVvTq4n0gPlEy9hArAEje2Z9OGdjSaI8BuwaOnEWdCcOox2mxd716o7s+JEtCOg3cGPXL2gPUA9
UGnW77sTYUT+rpQz9bGcvpsjBL+0nzjLn3zSJ3Bw0Mxfk/nVNRKnnfNSXbLSkZs9T9pLPYe0PsaJ
zX2S1kQgj9x+a0lo2VBFvAOtKDxnXUEad7mF1fpX2VoC+I6aSZJOeJFNqxETk99kp8jnzH7+a9ro
VOR+mKdI1vY4NLNlKTpCqRnVsIRfVSvg2ss5q1EdIcgsMbkwPzoLZePD1WIWAYVXb7pDw2DjEJDS
sxY3YdNsyxOKCbZy8m2X4YNBdTwHN8YbLCWEhsPTZxFgana0RPWbrLCDG5OHobJ9vKluPFfmah2u
wosb/t26YF1+LukGlEcQ5h2SYP72XmPL2eK/8pBz+nhkpg5tpJfn0NLTovcPS7T8CsDNU1XvP/OV
GZgGGxhiU/eEaBFvERCFyuDzAd9CP+yTbHXKd4rPzTBF/ifwj5KSgbbDcCO98tzULlcp0kSNZVZ/
rEU6dDwImWv78JEEwTRUeY2ceR0QvYGiMztO0wE4TLwUIUXR1vuc9oO+wduca/cUOwlIgx5YmNpL
MMHtmHsJxhoW0M2mdk5qmC7R+tgvOlXullBo5hI14q75rzVs4SLEx7SEhOwg2xXbzS+lSU3Q8AwL
6qBcKk5StuHZ5UbkgkxvfEfgWFldD/ORigdtcH66ofcrh981YXE9Pka3dw4MxYngwGf0FN7/zTE7
nmum/Uhz983owePwQRsTzhzMUUThH1zEZF6bKzfIOKqr/YC6sYvhSVMVnFYZ7dFRWPqVdFQotVGp
pLzjltVweyaPpHaDdHdrVTjvRilygVb9pdLrrDTi62SmCpQvJeExrMgBGmpedaT+v/XEF+Gnmzbu
iuclk0A2D4g16oDBvXqhb9TvXfgXa3iHjvlFgWD5mvgRx9NKXn2MiPcwe0OhPQRB13I8VcxJyViL
Qd0xEp+xUtdiOa3Xq+V1p0WZ3Ixl/nFOq2jLKau2uhuflLi/OVdekAYK5AAwlH5h9HzYRSSw39wu
q0t+zZ41aQowXgB7uZJFygn9w6nlQOVghp/qmqN58Ugi62QR7V6QLHC0+rdxJpwmx3zq0ieHAFHN
In7TmcKN2V1P7f6ZWpkY4PQgEEI/alrhOqBS4CSibXcgDJVVQOBSsDo4uG7W4i4H8W2q2q/cwohZ
2HbkowOBGUzIiKQcKqT8FOhCHMPM4mKaMGX2nMQLshC/mN95gPDUktgjXyEwLx8FR4hD9ehoHP3O
b332PWd/qajzTjdRYC5jO8hIAXqo3acOtWR19nJ5MkpWedu2lTvOQj+kco1CBuR9SgOD3llgr0oR
4UIB7zzKrqE9mEe5FTg8c4712EBS2wbb3pUSahXyy0R0PuVmFjffoG0yC3m8E27RMnBmjvwIvjE6
xtKlFKVA1o6fu86MNNl0ti2QMF0LqutSsqLq5YITT7p0SrtCyYd5InzHnRpfWBAsn+rov4GbwDfD
BdPal1II0f/5tn8UdnmgfUzB389gEes4BfKy5Uj3bnSsW4I2JdJ9ttkXbJiq2rzAdB2ILiVcRz0d
DZUEVbLA2atlytDxUpAbVj+3NbS5oZW78ygn3dYId8Lpb9IkHkdNpYYlNmfvdIn7C3Et2AzSLYj2
04IMlEx1UHHNfeJdzCHiPzKElu9pehUJNpl8i4cnM+KoLmVSutNZ7rPPsFcKYrghnUGevHBNV2Xm
U4bDd6fDB/7bSgDZ3c3B3YLbD2UYp00chi+y9BatT7PXDa1zF7eqwJImI3A3oOgqOCAW9MyHpzgI
qL9zX0T2t/LbP64qAmsEE96Y588LzLz2OogWbjzxPdQ8y1zkvQajwQJbWVNQtW38jRHj7Tj8AP9c
De4bQmcQ2o8z9K1GI/2mmQdD/O0f5ePDfzkynEvmEWfThwpRQC2aIhX2bTmLfOBec53ScqZMe8Kj
KLM6B8IkyZZVC8U64mG2KJ0ss8uoxM6HVyMKYT2aWsOY79tD3VtqdBX+oe5OMTMfujtdD71zeszv
5aE3odg84ECmVED4f6ULmIBDUVhgmNVtU6PUeXTEP2VQE4Mk9ktDylY6OEYU1KMkAX12usddlStX
GPgZ8vVK7/qcSHXFersGwjaQ6oPN5lQWIfOtvegmIvQ3E7XiMvJefeHNO8GghXtxO26z9/o8N9pl
GcTwUABizdlq8PSVJ4dwKtr7hIvdSP3PthxbSoapQpJ0uzMPABpAa+4gkTEpBN3SUGr4W+wbitVM
XL3FoKb5uMFppDIeqIQoRR29JryYPOzPyUvDBNM62SUVpIdts49FARNu1h3vfZbDyrzBJ1Z+cD22
Rr8KTybhSRc122Hy7wQIITTYbFXBPQEvsoPokHVUEGxiGtGMRVpX96DiK2Y78TDV59twQcx70cgK
1ZZFnThktQIDw5wf8aKtSx5A/jSNJZQcSdmptcdirMJT4E3ztPA7iZUS4rGMa5btWHqFC8tq8Hqa
FIUlEe+JCaEEclOlumlJocAxrcUDhG/0GsTFCebdYaWo0Nz684JLQvILc3uL9YcAl2YGvrPVEmMX
IrwscXGQ9uH2+vRv8OpyOEmWDDZC5mW/u7xIuLE89UXb5TDyhh+Z2ubURBNaZZvUIrVo9/bA9VXW
m+MykUSanZ5G7xjv6I4voJfAMp8qYk4fbWiZWOcj/E3mn7+wbTb2i8aJKBZOGzjmSs39WDR7Zz7k
oWY2Er7dsAOWMjAuARroIG0MxJBENgJ9eK8J0iu3lqqB1ADtmlMVHINSFwVjNxKUzTvvFwvvYTw5
BHJhCIUstYIY2ovhUuleZkfx4Z64nQpFtzjh0Cao3VfhkTcI7TJYPdqNowAdSDLhfX4fs0XjXRtD
DGY0FyKnFS2OkDARhVk5pI/u8qEjF1JatOsnHDd6HNPrpEdV+E/fmiUGa5gazArodfkWcS4J55dA
kCYh3f8elu4iN4Sj89x/OP/7taA1GobpuN0NOP6R7xmTMyHI+JX9HXYd9PiOHuHR012FXn3Rql6X
uKvIq8xSgyQH1aiTh8O71XmUFPYYCO7KKXfBXu28/DjvjR2FbOPyK9RG/zDemCV7v+aaUkjtlp7+
LI9CdYKnyNIrkXUbKZfhOqliGwdccO0HeveEVcs4LDvq0iPVs5yFsIyEFdRRBe1Ibx4/FUtrLI7K
yzN+rfcUb6DU4PFKxloCoZ7nAsXfq269nvDf3x3EKvK+FP/5GzlGB2EG1SvLaqXwi23SbgS0JeUX
eFp+ZMI7XQzpMMouYlQq3FM8yzSVs5Brvn3HQqwRcSE2FLInVGLd95nvVlAkpkfoK5+4Cd9iGoz2
YaCbFCacoofPVjpoKWBJOlCUnYb9eYok/R/D/8HmoSX0xXrsX7BkLai+5KeR7wrqXPyWU2VxMSgH
aAa5+tT1kPkxFzA/Z/jjyYwpx/iRm8NQMW+7WGBlWOMBcJklDUR7yR1HJQR+q0Xnz7Lrc0+f/kqj
ocNd81XGtacbh7HeWWL8lPLnjQyeJvueTlKW1cjZjHRZwFWfVsANUYLnTaNM4j+La2T1WVD1T/pl
5xzJ2ldu7zeA4DLIzhyqMVP3zTpO6q+fZmis1nkD/PcpZ42EEszqkgF8EJ3fqSO8F98GofQLgU+p
wUqfibNqfubqloxBcQE8XJ4AUOdrhU5Ow0GhX3ljIymL41ZO6zDcKz2+AogL4XchBxjIzqzxZZkR
DxmS4NiSWaGJhEzc3TmWY+A7sRh/JMdmUbw0aeh7hJT5nCJq5AT5+sTCX+5IcfPLVXxn3k3wQedq
OgxlnqpWgp9wrf7DLQ5mmzZ0luCUnZz1X8NFeOrmi6IN7VCMidkcXmKmFb3QYPfEKOJQO8EPboO0
Jzf0dF2xnxLdJj6kBPzyKpBtLn8exbIrJ6EbekjgDJPe41oum9hQLpYisE0mf8fLkaTkFbUJyrR8
tXhFxp0bir26myXR/TPCTkzqxwm9lhMsHn9zoOpFfWs63NRzAUpfPe4qoBUv4dS3mt5aV7x3HMtp
xgFxXYIjd1VI5/dA0BA9UqZPDywtHooivWewINKkYqu2sGlffj7bH3Oe++lbXKKKM/e9OUitvLQR
9snE4bl0a4Ndpj/YLja6VBMgGIu8RTqDUADpDyX155QSGuVwP2/sMKjM3rvLXGcIB6QPdkaSP7UX
AU9JXjM/+7dc9yCBY9Xzi8pu0kxzUZMypXVR5aQPFEXLkCHSnKgGRMGuHdPOmN0cfFgYwcQAFq0i
55tkX7jo9JWQzdiEGaGlE1U2OTDt7uPVQIFcRfWgmVc8jh2ulIiH/rv/L1RNkJP63gAplmcblTND
ytTSYsJTwBnccztOG93VaGHi03DlkNf9LCgu8WHl2SRJ/MUMcE0pPLr1xeSLiUvYot82AjhlfmEI
mhp9jVmVNeTBi9mHWvwyuI61XlaB2jeACq2gt/fV6cLcQkt00Vm7hyxfMBWJETlY8l69pDndF3vQ
kPVeCOVtsite/wWP072ZRENbCTJPf/jmY9ogdNKejG8glop1Na9O03poHXfxpTBiqOQxQNSNUhlg
V4GEshBM+eVRLII6hzfzDlu8tFg80peY1Y3Lxag2emk2gUau9oQIlpHCSkiqXRdHoO3wKdlLTfvG
P4VbxlNDhrVR1+lTZZ209lEAOOSg5Jtj7HM5KqEhg5xoobFUDZTT+3gQjTOH/T+0eZzD76qn4Xj+
pzr1tgzdW/sWiKsMgtsSMGdY4KJpdoa9SLkU8JjMlCxi3tFCouUDZZAwkNHiy+1obnwqVBabu34r
Njavs8CStCWz1IbckOERwr0+gIw5a/Vw67Mu7xHuVNeOnVMQcmPPN5P6GImJyBEE6LPPxvG4RliI
lcKEDT7O1TQngr4xj50hRXQkEyCcLcu3QXDwOf5cviABB4XeIkXCQbP/2j7deBZImY7JrbtTZC1y
RBVyjXsYCLdetFiDPe6hq/3DBh6ldIOAGFxRH/zkYV8jHe1oSQgfZCNWXo0kxemIiCbgX1di/iKH
XQbNwxY4GbtfiHnCHyRUNCZgoICZyp1Cj6jZhMM99HyTjFW/yIekffIkp170EVZHMPIRkHjBoRm/
tYrXD9af5QsH+aAsHsolvuWedzP4qYO7wNJSPvGGpbmagmG8UiBjZaEIPNkW7Z61YmHvbTcTFg0R
Su76c37wBAhwf4ElNtD0xa+prQwarBx2LjHbBm4X/xeAm6YE6y2VOoCXQWSi3+8/CvpZxrIoedz0
wbyr40nu4gMy3WJicFVVmGjyGNSSMjwT4stiTTYX8bbhQ7zOOwhHfXiCbR8kZa1OTit2tVZv6hGN
F6EwYTL8XPnYdkNLUGe3kR8gUmHiUpqot2lPhQGN2sL/+UakY4Wd4kqpKaqKzI4YvD5OQSrf8iIp
6lbWEjATnwbB2y47GcHM67MK7+4ImWtO/rQ58rE2rz50rw7KhyfBdPrdcR5bTpwTjRUu9HxcRO3F
E9sqjzaKzCixC6OtcB1pTfggIkc6CkC3YuqWmhorjBGrMg8hDBahPcukLV9w/K83CvTc7hDP4a/y
yWTL0X5f6LHKtNvZ3XQmoJIjs+U1JSlAHmzs/ANjKNrCWKdz4ITb2XIVvikzWLo2/zATNQ2FOqJU
GnIY/nzbzKYrIj3gPCIqWGCm9F8/sZ1tNIvwtIovTUYU6l+BqN4BT/V3iH3wabygJfDEpO9VT1GH
2+0THyO005ShvnDuDDl7L+moiHrRvdaVkkCTf5cX3iI0SYkmolR3OOSymUBxc/ZxYBZKBVSD3SQ3
yQuMJde66NdW2/zEUN9cMHlOx9Vd1RWidjKAs5lEGOUf4pZuqtgIDj7wrz4ERv8chF665r/d3WnA
558qwIxP8HNHqpAAnwXN8svQgTXSygS9yvEgtY+GX/HCn9PgssXI2Jxaq/dEsZHuw1Oy2sljNZxV
43FYcw3I8ZHgyi8YwvqyLwDRs7Rc5pPyBizDsc3cXb+iSKqAmtYCoscxDbQvNovefRalZ0aX015h
Dwck2ZD4OU7DOIyEz6/yL8jdgGSvE5SJ6Xjie2qioSykoqFk/fEs6jcnVx0RItJMZVAg2n0NE9Zk
/S9kaHQwBLXaVoXlJoJfSigEHQtapHwx1jVSCeZ6b7xAQ5/OfpPbyu36x21YFpHwteWAbZf2/jU/
8w7tlu9ASMtxLHh4p9XHnogDCGsUqgKZihyhcH81nsSvsefSELfruHddmtvtqTHQScqYzDyfVa/F
oXuuJihHpAhaFbT/wTGDkaAklG2oac6uRxRm5OjOIbe1bvbXSXsRWettFkmVZT7AIzQ1p2sF+6uw
sS64MKqKecV/ATa7zPqBEzSGMfVjP9H80a5Htj7v8qJ9MSA0yb2L49ldWOG1jOd5sSjyH+tgP9Wc
W0LKlwREexhvnSsAgIqvY7WJiemSs1skOSFYNGhEEdKNs3J5cOuGp0QlwkHINngZen/8m3jsefhR
H9yFWYpU7oGG4GV/pTdtx14Sr9bZrxMXZtfA3vXb1AF2iJQ9sHGrDD3/smaVXoEHUyVrVlcvobGl
O4AQ80OjJjXJcSUTpJGmwM0doRBO+h5uyKJ7CSg66zDxwWojxIbte6Ts/yuGEG04idbAWA9M2Ed/
+9v+05Ze8LykhsBX/SgybADHVpnkhjeZOnmQjUat2B9tjBY+0MZVr3ld5E/eiThmQWDGIQx/coGj
KIHsdMTT3HUOvynUI2grnMWtXeFYfh70ANGwtfufyUkADlVAX/b24blEd+weeLbLXKObQtqtQj+c
KrGIYfIm2o8S10T292f2Msal6sEiBWid9GKdhdciVshzXukJDgvx/U90VGUsCF0necxZn3SfuowN
iDy74E7mwBzUQ07/Bpg8yd3dXuIWNR5aHWqsvQ0Nvg8FKAFZKmMLJeHmA49aWR2yXPXJlYnVl9Pm
X51pXoARTgJmDPNj0TQZXb8KqqG2kTY46OB9F2gU8YrPgqSzb+/hSIySpOX2wUfqhS75EdPFT52A
/rB0BHvWsqAPvD0rcyiOPIvlR3vaAVpvCgq+DXYDRGyyMb4EVMqOin24LuMmg6kCM0EU2OypjGDB
PJmKWYEeZiGZWUo6jYpDe3iaPbC2qQaY082dRMnpiLmOzgDpaCRfroDwgYELvK9lYaNw39XphiBD
ygkYfavo0vuz/kAObemVmlBnz2YqgqA6o0J2vqlfTRUNZMvCvNgkCba46XsUrlmUqOHXc09eLKp5
gVjUBgNfI1fA0Wpnzr982oQi5vylhTAeE4/HLdMIvIsijDU8z9YUQK7l0hBZNd3Z8y4IyWfgJ761
rVGuX7svDng8dY2h2GOcUvoMqIK7MwKjS6c6wBiPf6eSpMDdY1zGrgzkh+2JSryI6sMtKEEOTHtl
vJLndkhq51B0ebVVl3dZFUPPHZMvxbOV9nfvVApJEgAaG5Y4VHk3DzjUFi+Bq2ajw9EklTEpyibG
GSDnqQ3uYB/nUnlVCpTT7+1zt9P+tSJqbSovRHCyvea0Q62t6byhf/yvdPeT1T2erNK82yMpldhf
AfhqkPImRCZ1W9LWe8h9S37ituCOPk+5bCFUx/m6JRZ9Ux3Iks75i5E2B7Jvsm4RkVo5so097bY4
jO1t5Cic5R6lVyvK/vJyJ1r0Szoaf59WwpyrAnK5GoT+RNDQN2KmHDgq0Fpef6qfw7+9JIGp6YZb
WWp6DSSzK3SqTKR0DP54dNr7xbGhSpOd6cDEoONQtua/iMCnrBD/C/DANmbjxj78Vcpok3HdcMdr
cne6p8bwSyMYVsa1o773OCjjpQN+6btVetuSKTatBu565svdGxXGFnMJMcc37pV3v2321ZrSogoX
qt/EUDt/iXa/fl+xw9YAYJ+qNLRF9RIuGZ1vXdrF0E3Geug5TNuw9raxVZ+ayrmsM9OH1B+KcYI2
/6g1Q3e05AHXNXn4PeDbd/jEcZU5kClOwTSiOYkttR7pcL/3YrJZ/mGLBxBTHd72LjYLusUSgJw0
bXI43PtHpm6BizFgsonbYEJ00FM+YOx877MqHAjtGkhywqp72y2/Trmgqx1908SOk5Fxd7KZ6n9H
AeiiHDhyRYiB1gP7+tg+0iU5rFsIbBQOSbJ7b7D4dX7GSpyGx1xB9JCoo5vR6k8C5RW4FxKUbl9N
UFEHGVbXU3CmHidK/U6U9/2FzmtV0J1UCiJ/BFi5pAs72DP80EpdV6kJ/Ynhr31wPJdfjgucLJYm
d5JTcbqlAvwUJbZc4kkXsF8+RLZLC88wAAiccJxF/IV7Pf3akHoPO3644DUxrlixceu+vsuRlDQ+
JyU9zBqmgfbJAwQPBTi3xd97FfnvXw6A/BU94AbdGQME+Z4TSy8bKDW34evQskd1SFpF7vAsa6tw
bh21LFfA9hZamQrfUoa8Q1OtmOYSrGKCkqx//ernriECw0R8yhk1LmDo1LZetoo9Rd36QtUg9Hu/
Hjo5zJnBSeNkj19LF0AT2lJTYhlOVeALyyTmA5E5Xpn0NRsaaP5wCSJc2uPpD58eZuwlRhG4iQR/
PhM962gYke4pTj/nNGIArCa0bJ3JbsvHueDzQyG1kJod9dUy+zqXBp2csX+dsf0J47Q54sN0Wf7l
OgTdEn+DEdusQRCl6oxXit3MXOJhv2nVQ2KvHiS7BD7Gl3l/9/3yUhMFRfXi2wPFhkY6+5cW754c
MXS5a676mYqEa7+F3AW7IDR67NBnU8lSkXa6WmDuwp2EDygXY1m/tQUwZRE9NNEqk0yNjK/yACqq
TFBQWZ1mkCF4JMpd4fmqDnW+OuRiHd5zZXEmP4QXxlnLxK5rf8Z2RbwpnNfwNQkJO7XB3sEEXki5
4ULydQqU7uBEJ1TbWL9Vd8mIAhUZBY3dLk8aahPn5Vb4Cd4G5e2FH7Ajq1DmfK6eWyxSwnJx5ny5
Ov3zgRBlDvM95HBYVnI0AdgxPtQxGaLYzViFL31HEhxdxMkXaLgrr2FzVRto84PA906g060gjJ4A
62VMC45Bg6rVwpH9R/y/56QT2vFodsTj8BQF6svXZLhOQJIy6XTqJ9EuuF51aqgsP6azUetlDWA1
wLVSfHZYNAmCUwhm3rGsILat0jiXfTOh5C095DDX51fM67oh/BshzgDFcit4RsfYOwn7wPPONhYI
iuYXAHiDKcI4miHT62xLBPazNWIrBfv8zmoXdi0HIm6wylAXzucTnB8cAT78i0A4Wzo1DLcaIXO8
ooz96jX145JWYs0vjr64wTR8CEZaganjxrvWhV0BemlaP0WT9tmI8ajz81sE1WB/QifnpFc11hQf
Z3N2iYog0Klzzill2wob7JWr6TpMKs0v4rRNS3pdzt7V+PLZBgX9ZAkIyCvcu+zngcHoE+DsbJtw
lpULqGfgkr/SoaZuzTaFLbhsT1AGGL84cALI7i6Tec1h2z0MKdkYpjsY0LUP02oS3Dz/N2k2jZgz
cPcFH9hF77/W1fHf0/8g3cyn7mqMkI2j/FHC1o2SEvBCHnD9GEl5opiVipWV7W1LBwC1W158BSB3
cGWBcq2iDcjMzItJR8a//Hj1fSwk8ieU9NcC8Sg3DyP2wuqQFQfNW53z/BQmrnwXKjlpiig/OTA0
qU3hfi3KNhY7zMLunpfn8WpOjyFzLUduqpro+PTmK0EWRQhpVP8Nxht5sETKHoRKCDQBIPnUyHpX
L/d+Q8uaNtRv9Zn6Iixt44iiCjJ7+Ii6gr2GZ/7o64vCmhr91nTBTNaoEaB8hLWDstYjHZeceFbf
kdij+/bFp5HOm2Y8zCafL5rjON85UO54sCx8xz0LYYmv2j+Ar3ghHLdnA6+b+CFMNGlEq6Npku9Z
MSBIPh6tH3M7edeoPIRNVmhGdJvSDUpuyW4kI+3IpiJPSzV5ITeTSZ9DII8q9amfwfnZIK5WAfqX
KsNjNW08lp0zB5VB9Mz12y5FeSe/mhZJ32/TaD7MnW5MCaOUZTTZDl0rUZ/4fHddEmlcg+tEIdoo
vUCdiwGS/+E0khQZ8u07+9/02E4Axqnm1tA0jJjs9XE5UWMyuvmgc8GlK5nSuPNq9jdhIU9JCL88
QbJTzhD4lKB7e338BUAJKQoO9FB4Nud2eziLoZoTf9fIC4lzMw7jECNHqqiBDzLk9R1W6EVf1Fv7
eStOg8jOOj0e+5TkTizK/mPnfJrTfKxAN67ntPPgNVBzs1PqXXv6443htoG1u4fUYQdZKmdWOi9A
txWLAkodQfWN1E1jbwhueIyhLAREzbSD9oOzWj8toyZkJVW2pBnbtHo/opcTdHAtlI69GfwkTECJ
58I1J2YG+dW3HZAII+pqAcREsQwIDWNq9SJzlPnF2C068fZ3nKnai32vsC55sAVXJOnJN4jZ0JK5
CmxBaoALJ8AuqL6W3sqrCWvSYcI0dxiiU5APckT6R5L0uQyuahQDKKbNsVgEkhDgwwZyYgU/argl
XujJ46qRmV9jranfCNUAQY+/lMbl1Vw5iM5VfVG3Pn7PzZY6RaSjULbJtRjddLkGgfA7QBNo6UoN
ZOw9O9oUNoxvDwVa3D8BcIHqfPs19F9c1OuhXfUmIY+YI+HgzbniwuQz6XrcFiCD895yWyxLGJbm
d86rkbVNvTCMEqt7I0wrQpLtqtsutpXsZD5BVMG4sMZC/XFmdq/Z2rBjpYQW5rrpoG+VGXuHSCO0
RDydrACDTFBvWGMlukDgaAbQNhQ5zO/F9iCTuvf5tpXA0zIQPfXaPS0OFMi6CcBM8/OpnFFrYCfS
cnuZwP/nn+DuS0zoPeU42ED82QyUaGCjwoy8OqBbLUEPyIt+POPDkGEHJe3C7nqIIhsSjR4ArJ84
VpeX/VuFOcZ3S7nqZpJlLjwTjw8iHpl2g+fjMCkNuP0MrWJjq+vlw5K3wr8K/fE2ObN5FEftncKM
xeakkPDiqVbl0+H/GC9ygxxLwzspWpOO37MKQCdYx/GK7RuwO2fBQMArDsPn470mm9XxDQeSqzFZ
v2sUjHGUggJMZLRBoHIzQLZGED7dkdewKTBkox1d9Tu0clMl7QCAkwCe5uKsSXAMRzcNCBLLDVF8
xZwHA7dyWLIwccTBl9vjOQ1wPs8eE8pgT/Ynr3Kys5YmnptgB00lcd2TDVdaziCb/sf3X9a4PCPv
MM9ZIzyEl1RnX2z0c0EMDk+s7I0QsY7KFINRz+le9W7BXMwtMI0tUDe2XjgJK+I/zNHcwyJ82Fk2
dB+fcixw3aNZtbWGBMBrB2k9wXtmLg9b9DWIEk8XcKfgw2b6HZYy+cB0OzFrcx898ok5ESug3nA2
dQXu3d47XnSMbrnd5tn2bNa6Qf9eJ+DEJEi0+HiNG/63DtMm/GOLxYwis2yYe+nzp+W/3Gwu8HpT
262MMYNHYo5R6BTiGsjgNOuBA8VQLIQHs+3XRLPnghF2sLVW0A+Kvi/uwhvV+xaQO9h5qHWij1W0
+wN9SdLPrWeCxsMoKQGHa4i3gFV5/wau54oPCReHdb7B+VogjhscDz0tUJbY8GSheWJWULnr1Nmh
HIgCcQEOOdLNVb67B7CDHcLUJAqxlaYsgEH3Orllns0C6zP8G19tGG1Vk702DEloL0S1bOz591vf
Et+cYfXG4DVgaXHbMl8WoLUYJ6CjguGdnzPVfPYy/6ehsKaNjMxXA9FBosi616iiYCD79YzZzU6k
vTjAm7Vrsc6d0E2x33C8+gqbcvIrrpds+gplJ1o+tKM8driW56jB1Igo1Z26Rvt67T/3Flpup7u2
NB3wcFhaQyX0WXLUCWoXJkNskuBuujX2UyJLHlXeQlErq5fgYU1EXfDGKWkTuU9+K2sHKTxMBa6E
axFpSGCKQF16uYpeAy/nFiZrHPwqFJQYrrg5IB2HGxjouM4cRrqMHs5qZZygF7gs3c1MQIhqNdpb
cXVBqaeGSL/S+CW92Uf4oATNLUF+8DdrQ9trRoRfthAtC46P//5iqS4pA2+ztUpHm51ljH7YA+sT
EUwvPm/3YV25/9l2Ngi5N3WuNhI6cjaEQC2MR78z9ERIkrA50RV6xux3SJ2x/gSGly045dbp2nYw
Xej41vF7jxtyfAdPq/WB6wyVBK1FQAVnqIlSqmzVQgR74bkprmckL34lzKeBLZZMTDGG8qRctZBL
a7Aa76BtzzlPF5xol4poFsDFTfmRRMtPjtTncigylhc6pV/QEddFG9XIThPP3dJLVQNt915mMuOP
08rjaDkrsGmn1xn1yytjV6VxlVhBZuG3fT0ZJ0JSRqCfBHqsdnGDIi6msQfy7KLTAdTW+UIUCaWv
pikdd9eyUTOEEY10klOMQodtsWlim9qLwyRtnxovjq8F7o//vPUL+fTbJycBR+RXhLnDs/39sE0V
JUzQ1235i7kipHBYljOzRSGXziIfYQHT+5Fa1u/1puHPoCNyVs6xQI+g6hTtYVs2g+RGl7FsHKcQ
P2S9HvItD903zHn6tgJhPKU9I/K2R9y3S/YwbQbn10VTYpOyzaXxh60OVmCECFDyWgTalphO0d7o
zgK6RuuF8RUWkA3hkrb9DZYqyMUFqJzs3GwTUlH3hWEyJfm/DrBiSRe95naBys9afa3rH/XcIrXD
T53L+Z//C2xG7EF6ppjZdTAFWk5op35IfRsmPOz8MlW2Ei00tGOofy9Kj51IRef2GCAy/PQSRhef
GVLY8dKBfuLQeHQ42zK3KcxTry2QwQ4jTAW3xLRVV7X+zh6IbqkWNdOJcy2zJKSzQQMgW8lQQk6J
SrIlbAluupeR4znGdc/gz1oEnp3UHDXBvP6POwkAiBPP3KH0o8Cu3G9Op/jOeVqiLFvWWvOCbMoF
DME3Eh87J5RF+DY6LGndhbTiAWk+nfR4VTEuKyl9EfPdexGsOgEqaRap03CtU7dS27asxP/gZoVP
HsRGNJBP+mFFVWEdmZ4jKY9Azv2ixKaZQ1BJFCGBW+0xUNaFZ/wWZEVRWrfdel3XN4z9VkalpIsh
s4KsB8RshLVf2QNgBzTHpYRTJf3yhoc+pXaaNrm/gv23hUkI4pfhAuY0KiPVxoFP0911tBJmEP5E
cLOMtdk/O9/zKFn4e+oq9yy7+fKnE8FjD3veg8rf9lSpAh4Rg40AwvQNI2ZxYq3uQw1IlKBn1GEo
BmE0bX1hsRYsMcNzXyAF0eZoD6gyMST6mmPVgxjDXFJ9L7OMYxzWOXZBooDpdbscXrFVsNYGo3h/
h/DSSNWaKPnKSe/0svATzf9LrSnZpHsR1ZhfmNUPDmtySqXSKLW5hgQ3BHXMpCh0rN2TYCNr+F+z
0/E63e2Gfxv2FnK6Ab99IMx8jkobAW67ID/UEIPQ8VwXZO+sNB52QPE2X7OxUOXPw7VarWL8vBRQ
9/8eMtGkrm4OU4FHlb/Ck6nLP7zJjqSLAFnOUKeHlqwmKADitYF5lPVtVem1rsoJkTvbDeo1F9+J
o3340N7l4R9Ol6wlVcajhHmZLfI/22+DA1eQ9kbJlbUbrGGXXcoD5jCCup6hT4664C5zGguKEN+d
2S0yO0CmGf8Vv92z46XlDTQjzc3RQts+7cYAF4w8YnxpvJxdMEbHBM4DpHL17yga1TpLHUdC5kwL
a8wJ6P8GHHY6CS4JzGjszQM5HVqmbaMEmWghqR0c0QSyL9q+0TL2t8Om8sR8n1GvZSx0884ToXaO
n8Tpj9/n/OWieyuPidDB6OyCj9nGjyKCX1VMvbe+5o9RjUCDBRwsoxy1rPyB8SYRl1rPgMvpFPSZ
EW+bbBB43brWHi5KQtH1FPhJSZBfbC2MrnZfhMwnKOX6BYKsyIgHnwH4s9Ug9dYNhnBXH6jDifB+
eXxqQ9HTOCbengXpe5NldmlDIxiw4oHf8ekDseIoxh8g2Mgkaw73foJHJzEM9gOfYwSe9v3sZM2i
w/uI+XL3Qke2L2aVbjtHEswJp9qC36Zff09IqvL83njEis+g9PGMxd2gEmWZ2rKWD5PFUTbyiDtw
HvfjtE3AfUK7C+xk/j0qzxqgWfWN5Lw5Ie4BdSY26m8zUVxNDVHok/0Bf6VH7V3a0CtxCSlzd+HG
vjEiMQScxPeAvHHLxN46pv2/MIfD89eMFNRhTDBdyPLdA00aG0w3xQBDm5G1iqIX2O3vaTgdJpHk
CD0M+0W2o90b5MSZZZiAN5k0RZHn3Zln7uA1qet4kCLUsP5tMkwiYerjq6iVocw7ocOR2Ow4WMEr
PPpYGgZAkwlx7Sy4jqCAYOuHpZhxC5Uyx+ht3a+u2IJ1VmRKfz0MkckFN4O9EdllW8P8rVVBpgn/
i3AfQDSeD6EFPvZEQJh/p/QMv9R7TPqPScVEOPuyGufx6SYPruojVV5+RchA1JSfQooSWUNLyg7w
mODFequ4EbUyCrEw28eC8uHzF9HJ1H/+ud3vYCIF/VHEybVnfzJVUBZBF1+UTWlF8++yQe03IGnW
O5hGXnRu45GKZLPyo5OZoYO4wPo8be090Fhm4xG+9MEw4ayLhz8BuYKhzPA1PCl9bF+pUT+bLf0K
1dGdz7LOq6Dkxg0yeahyf5JdSvcL3kds4KZlfpWzjtfOi8CbAfkjpXKPWQvlWSW/GBFDsijMOjus
tQBVqXP4piBb0TNgYEANJx3m/qpBf435XGTuGb7O0SlPwkBEelUHQ6+F/ig0Rtsop+3C94aIU45d
fRTKDRdtKm4hrY6WM6o9DDAh24zd/oT+rrhyoX4/7MCnXcZD2IJ3rI67001OMs297M0ASWGzs6g+
zAcXTf2RcNtQVlAlaV/67XgoO/jQp8JN3imeHiYlYOeaoJtcS+wrgE6Xh10YaEDALcY8spSuAko8
SWaa7N1rhkyIYm1DhSKF4Zhkuk4tp9Wc7yVYRDfQ5Pb+JXQP/W3DAY0UQylNDUImRzD5O6afe/3I
WGRtdBFwNTJsiNBpWSK0mnIEzO9QIvQGosIsQQ19VLOshbYoBRjm3jcYbLyj3N1u4A4v44fxGbpY
JDFwcjvkxPTW68vyGW9hUPBrXT1p0XTfsJH7d2qMsid7tQX1KNO9TfDK0elKA/4C4YUzPt/p4WKb
GXTU+sadKdl/CM2oPcR5rlME1OeyYavc6GGHe5UyBG2kzEhvq+zm/Ex+rsaVKrmOH1mxoFfc8fKf
HFYANARpFBmQOOLB2dxgMOlXBgCJvo4XmRMRDtr6y9ptXKrriRVjO0F42UkDms3unGKIsCX/vlXr
XlUNv6Ku93cBGS7SnLkTnxYeMtt2twYf21XzL0hUWu+ed7gqu2mg02kaaDG3ev84VG6SlyTP4t1X
132ktacGtg/xLUZbVsnSrIl0FOjUhJRKwroXQ6/05ApfoZalMSDvw9o60unwsNMPmKPrHQWO5xcW
dey6VTg7PCYy9lcBKqYnLEiIA3O/+FG17TPA0TF5GpyARwK7QzbOt45w1IEHz/ZZAML2fl5RhvKk
I2R2NgDPd0/z6KRRg29AXcJuCHd1VRhUUr2pdwtgKSfJfWyXiK2NJj7Md1zl1y/PORk2GH2gRavZ
InSPRXQb8TWkfnLjv/7LCk0k9XNLK5mTenxfsLX9BM14h4YnzP3Y6fSOGhD1CGlSQMhqLRxuVIDl
HSZbDU6b+qkjD9dNY1OB+zMxYsry60Kq7O2a2GSBNeMhCCwahrgiIcBGQ0lfxC5mZYGV0CMaVTVa
zJNUebYVF0FP99cfvXhwn7jh99evBlpefmIV5+pUmJvGRguUHTYX7JrrVSoxNR3XfgCSF9cQDvrp
cEurWWqQnvhCgmP7Lsi0pPkH8YynUoN2P/hFg9o1J6B9pIkLDgVHG4nm9Wlr9rqcOUOs62XWjFFw
WaQgK5STVBISdCqagQVPGWXJoR8+56nu1g5ogx1SWZZkjQotJIulXF0ZAoVN1jASsMmEAmNJqIzQ
NSUkOOfjCHE+iRPnchShtH+hAGdBO/Lu/BjKqQyj1zIBeKPdCE6x4G/rEb6qjMCLZdSg3/ooRpJM
t+IxTx3sp1MeK9/IP1aYBgRz8WQzI3nNNTVM/ockLJZ2mNvvi8431mfkkI99rGRYU+gIexYkqN97
qCFJ2lwqrZo2NIEyb1xuz0t1TzW5LYuUz8VJxLxKSEWEWDtgAT6/QQufgPN05952kvH1oTz1HsII
zPDlT587eAr65Bpey02slgbt5pJ75Oj/ttduYlrBE1bTmQul+Lgdn1uGI3j2oLmCs07HSY3jpIH/
38WDFWSTmCbUrItvE55RU8nqFSZfgHA9PDbSQlglFlJeywMImW7flwI4b1FkFP8oAN1pUXtfOOm8
igl43xwyukXjzB8wveCFoiWzdcvktWi2HT1n/ZAfhjXTnTpcF0ch2D9gdtylB5GmKCx5YGJRcE+4
2PMGBjf/Y7BKfJaiFpdaoHxDsrZJOH5yFZT/4p6MEX47+nriazAQ/G26CLgiIvxgjZDG8MvRMrpq
JwepCSE39O3OI4RVXFYxy4Mh7XRS/PrEiqP6jzJiEnv/vK+MKSsZBe1z1oNdXVhXMGH3y15nU2UQ
ks3h3PV/2ecRIgcyMD8595MJOp0SoIO9xqbjIN0b6qMyZOd4b6EjCRQMYNGazO/c74N7GuRcpj5Q
FaljkKWBuN/xIQRbEJIKCzyFfy8h6AM2YDDLqqDMy2MaxBANoZZYG9nSeakYB2STXhULzQQYMaOX
Qkg8onBTPKiv7JEFou+PYLN4jjqpUt98uN2R2IWZ1MKdSwPm6orxWwK77tGpd9hZ2w/o3g/gVodG
6yuncRLta7k2tJm7Sal9mN0JRXQPqL7rD8gxnYibI4EsPQwqvZ9C7u7+1MmNkIHocs0FVNptpAri
FKvq8nSXwmEyalP4TeLxAahIfMSPYqM14KD3RGRzAIdeZRLGWagHLPRae/W5yJnUAE6ojYfKA5uD
WayZj/6bB8KXDrKJ/RPWUhTOM4aX3xPbbwOoRc+sRNdw5EzkVgNuQTKdCQ2Kv8ZelR3u3PiCkruY
j8ayLCIXWxZ8xzeNX5JWpeftMKKDSHcpw5AnzgzyM98+OWfaVnP9LP4+qu/5Ft14jqBlP54DSvrf
NhFuP/oVbTldBKh8TIahnHaSxtBRVJIzlEW0SzcWdN71KU7Dhcb/o3m1MEW7cGGsAXDtSV3e8xc0
gQoJ+SBser5wih57tpbLr9KCez75dyMeyS5qLqJz7xfpJkVnQWFtA/L08/IjfgjFH/M/CpoQJucZ
62C4yb77hdNP1HI3IB33Uw94O2ABp4Z0S/TjOoeclXkjBMS+CTLcyGl+5QD8n85wJ5zmafPMt3oR
XFyIhcxCnLVkaA9FlEewm0uXi0PbweV0XmD4MzV1J1v60OAXgwU8QxN317BcqHa4aHJRpAsv8HgH
XYpkq7N3cTrh4vVaz/OhIHZam3oWVxYNhA7lp8MJBj790VTmCMZKPa/SMjlq0by8l965XnDYQk+M
f4AnWYrqg0WZ8lqBQVMzOVH9go6cEorvqT+04KyuYVu/Y2p7VToljW+DA/onivA/F+CUq4LheinO
0N5JRXu439jxPe9fj15A7fHytOYzPCvmtwd4Df/rA3+L7MbdAATmYa6i7TouIjLwp5XZC49J8Ln2
Tp9xj6vsuOBsyrxc99G04QqW0BtMqWknju0MyCWrSjIj9ReCHKa/8qK92Blr19GkmEaG6FqISndQ
CehWEd3Mnx2wt56byNyyb+02DZwBY3mfOt9i5zUEKpp5VzUL322TBN/WHPcJHhDWqcE0KMDeG1v+
kAOwqbmUZ7hdcDInAiKuiONhv0uMCD3yXCTwCrz0DA6eMKnoKxUfseV64fsTqfY4iXXTml2KvT6H
hEtWeQnfGD10a6TpyoSyCONep188w9MizSaYriMOzDaxmV/csUcofXf539IYjqw7l8UB3EVrco1g
7tv71OFt5u5YlnaSeyXWxx1KdjWSktsAu9SidAQUSieRNmcYHdQ8IXR2O+x2Ei43TIuMx3axM5Pi
mnNWl/moBmIy+I/gCRw9HEeMuK/iu/YSYbCV/NIhre9wKZwOWxq/Drvm5ZTPTkkjHJGkdxXky2d0
VyKSejSIZDVM5ZlXxJUjTY6Di8l7vIrQWi5SIrbIQ97rvZfhLcHDHQile1CDYYkon6VaodyWUaZw
u1jDGTA0XzJubuKIHZcRhn1IeppYK/IFFvPnf9p0XkiEnfn9Z+4J0Et7V7c2J4ZlDPGWWejcSkSN
SAf7ErsRA+umcPkkvQRg2rIGnigvUfePy/bvILqnlZu7dhyh9Ppai2QQJSEsP9hCRur5KW40g40I
2csv0auXEXXjzzC1y7WdfuAp0IAPw0rZn4GX3URjZS9+Tp1iEBdim61I+V36oq10k7OVSSEB9vb5
q+aSmgUcCl9D6gkTabmkLGlHnz8/ZrJVqF6PFbPU5jcn3f2Aer2Xh3hyPWfwRxADrMQIkwA1GlR8
5VwCWrKhonYyNmhXlynxpU/2s0iN21D7S3dyWdtyuzFcHlSbmrCSH0yaUmNwz3AoMc41D5zsPUrZ
x1Gll52tA4xWdf37KXYFC7CAuNFJDDTU7kXT/yplImvg52nJ78gMZ6O+y8bVqkc7prKBgQpZ+8h9
FHnY8RSbK3rL2fnO0mbldhvjOkRsbFeBR3tS/F4HJVwg74nyTb1TEyAJMl4EMyd1tJ9gvV16ysqh
oZBMuBtg/Uz2mz4BoC+GootA0nY2TLm/mP35ZasI4UFAhCytVAY5cNIAReOA9tqf/oAOtynMFx8R
vREM7JhEKDg6bYk++QD2w6jkOJI9RF3ztW/3eb2E4UYQahV0Pqdzjjj2neMmTHLFkx726HDkDmxC
KNt1lnTmApKU/Ug70XkSjAkztar1xCdxZlgDnE25DTxaTy1qcpsz3vJmYTKW3HxgtQw2OCIBvSY6
65QRx4DRquuRlQ/SvOEz9FpJ9W4IBBmvK1J0cXXEmzg0zw2I5MrF8Jh6VtfQCrsB/riKfyEToMu8
Kr3bNf/beOuOfoNOvJbUJTXkZ3yCeBqh2ZVqu3+MptysqLD/KYvo2lBci9GtZi6sy2kAyVkMiGsS
+lrCmm10/qYMEume/a2MFkBStBL7Sj44KxNm5tEREDrImyTQbfdnhxaftCI3NpXMJVpjyF5DTHSL
uH3C70p0z55V8uiEPH6N2qOUoOsbnY9k12bNfHY6Td4tXSdhfG0CuQ7Ht2j99wZ9S4kfxU+sLfd+
u680bcFc4Xt1Nf2w0Bbx2VHJqU+U4mFwvfZL4IDy2UulJxx9oDvp8xTmMVedL7ULEKkZroHrXDfm
J0KOqJgIZ/sYaLFIm9xQXypIeldTlBz2C5gl1JmKJiCuOynSxyG5GnuJjwPgKxKNvUZr9r4dpNeE
DzhY5ArjFbmiHzf8yiyHAPgFtSFRr6V5E2xgkTlpnTxH1r76hv+fmuTm1U1niYIBqQxsnFjmEgZp
b5YoZML+WQ3XWRJq3ViReAa//xboe4H0BVEaFUgen7LvStGq0m0UcY0Guxlp+rV1d3vlrpu9WK+k
lqOvZ0y5Qxl0j4ickRaNf+s4M/baiUNRo4jcGfqsPAThBSnjPkiEwVZ00ABrygYp8trRNdgWKwM6
5qDuFgjFTDTGccFzcJu0QW0YJYAmQvj35DcMBY6tslNEtnw6j2Us+5wsMEcrC6Fb4LUgaix1gVWW
HISsUXD4wfPOD80s6kViJ7lyhtSsB/m1HHljrTAOl8/SvlRElytjkDl6ZvRTAbfDUB1JoOpHsLEY
MaAp6w4Qvehh85oJFveE5lHrLqEeBzGLAu/g3VJsxmTt11uVFzK62WHavvnbvGLA2dxQ5kz3fOL0
iWEl/nrsJs2u5GG671PCjAK8YBWypPQhoTXXQBPzvmTpWIT00llwIP+//ZgFmmuVEMHameBhEFDM
l6wAZq6maA2iau6IRNRQDf5nuFaZ9JOCj4gFtOEHeX8P1539gf+1asFJEZISV/Vait5XbCMriFla
bi9FVHbbb5rd4pAYlNJRVMP+nJFC+R3giPQJ76mZokb3hepa6crDzKHydlofxttVUqbBtecBF0fl
VKdoHqtl3hLPXjqKE49F105qWjSrfB1f0HsboSAgmcuc3CbPqeV+P3/I/jcuOLgAUY8ok7NYF83O
9BJe/jgz8yWzFMDLe+dXdmBNlnIRbujCjp4yB4bP4G2ueRFm8Gw5hbBW4t/seIQqS+z8RLL7cb6W
S8l8TgVhoSTmg0wpXtGpT+tGwUXuPUH3R3TK4jnu95viXkrrbji9iY9dG8mC0ZL2Y8P7aEFPBPU7
tqh72Tal2dNzCLlPlIiX/CtGJwp+PeNSBydJA0EcefpPK/sveo3yWmYs0R0SbakptrN5ys2Ur91T
R8n5Cr0TXQiH9hJb7UxfMeW6DIBQknLZKSYqxYo6x6MbQm0x1yJG6s/FySmdrSxiLmy6oyUrDhDJ
0q7CyDvkK0OIBN61UP1/coOeNVyxzPxLHlvTy4+MQ1vlJ5okIj8V8IH9J0vkVkUZ+MpX7RmIQ61l
SXeVhZ/hYvQokJUrBpXMMW3sSwSZ/N7+mGFuAbtpR2GyIhENcydRAeO+YwFF+JoFDxsao4yIkRLs
d6HsuZon83AXnriWuUdbukmCxZXftUY4zV0nBFl+ufEWXQLJVLpvXrZGLeoVOI0107Jk3B7KH0jw
62lSgFRt7JVXd4KbW2JeGPF4UER2mS6AABeYGNmrgN5sGrvIu1V93LkbUf/2fllLO6VeiM1ms5JK
z2FlcRpM/lK0ZYfgMWusJ2xCWg8GqNffoNdxvzDCHbOqgPJv0etg7vkCOw+bBu5UzyxSRATPfHH4
Rt76FAFgAonn7ykWvnmBjCE4esLWqpju0JdvRn9WVRClAT8BeEUgOR+dtHCIaSVIQHHDB7hejuTr
0qFmOcoM3ObHn5Ebvd+kd4P2ThjXQTKawd8bCUz7KNMnBFAC/9cHO3+xHVYjkJ6uFNGatP5ySXm4
3fLVR25ISWTXqW4PNMYieEMr/xFf3/AQZ6xK0QL5TSNIC/xkEzH/dTOA+oX/NjSR7h2tGfpa33Zm
P7oOUEHLPgZEETF2aahAyovzTVROrZqGq6MTcqounLWIAYJSkvJk+rKtjgaUtxK6mAejW/NFEHmz
WFkbSrAX1IO39U0B25DkeRFKogjsfZVJPmD8eQeXFkHhEJ46muvLIrXRp7CL3tDyrbRND2/BMzLQ
lw61qEgqQynZ6k0vCMcvW7u3SMZAFSkT7ZD6x6a7rw6uTJfguNLDZe+g9oDUUTFBVj+PdK6DO0Kk
U5f575wyD1rzqT1STdwguOxUTEuX62N1P4Q89mREfPz0mrdbOOOVMSMvm9BKpPHeGeNlwxUxYC3Q
8jrNGrlstZ2EcJycFRy/B2H4Xg0Yh5Ya+W/CYIFpLawMcybzMUq/tDYuXZ06KUw6tssKWB3JKF9m
gyKrJ/ZgMiOyG1vofFsptAkpUNuOq6n7MZQIc4pelgcrlf99NPG0cel4nCoKc3+7s3hMjmh4Ud84
eLq5Uu6vrxbJwgO+3gNZ3mnUbxAQxsyP76qFiVUJupLmMHU2vs7M4EhI+ND9ixlLCL9fDOxD8Ntc
8QHhWbJN7pGfSH0BU7BwlZCkbBhQkfiqzQJ7UKXEJotqCDzDp7uHE9jG5NVf0skGmiPW+Hc6fLFn
JrqL4gq1Pq5fffhZ9JQkRYl/LamZvPTHokHL4CoJJldEl6obu88kNqktLENo9IA2Y7d8IsmkZo9y
4dS+3MnT002rv4VsEynxpask2bfOsED9bM9FihfbdEWicdeIGz58+St95+0vvd6iY4KoZMQlfD3z
KX6kNJtQnA+GoQNXWSrRd+o6EFYT3PF7+gSKfeJmqTgBgFGHm4hLTOVFNoylfyg4wg2EcLEs8+D7
sDRgDfgRwGHWR5Ax69zNBiq8OvmUwCpMhEbnhJUJyySPGVCwjGDNW+6SaX+1xqKsPGZadLU7HL6K
vjNoyETTAzx81M66XXqg0aQsBd2Q2qM8wV8Xoxl0N1KbdM/iQPnUbYa8Ym9EDUYsM+Z24g8kZ5TG
6+PhzBPNpvgcEcxMhOHIbsBs1oRsPijRSH/DVfew/XvnJoMOxFjMBP/JS4k/IbYEE2zaJDnKMJvt
o8wmBqZEJX++QuVN3Kyug6Vw1YwKUykq/2x21LdgJ+lDIk3JKPWnoj+9iCcUB8uqe2NuQidXeBBf
Tm7+QyGNrfXAuFn/pQAMKs2wKBjp4io+KMNqcbfTRbupDd40VTIMP929FJPmmPjR4vdiJKSnupCn
iNs1yuXB2XaDa+mE22sa3H/+vTgFV4SAQ/OQnXQeZwnm7jHJGP9vqQlV2TedW+NBBZ3TGoKiK/6h
ijkBuok9BuK8V6O8nd+1KgUtEReEVD0s3jeVyV1aOBoPVxTUsCZ0iVg3kFFbTRp9MMZfbPHYZfKR
bEAO4wvSpJgOPk8IZRquo3Kh2Uuuct6o/Iq57yo46AjRg3B/iCbB0oOMn/1GBw5dw4Yh06ydC8Hs
TyAFqjfRwftwGosW4x2qXcCkXCSlMR31cCHEd3tmcU9Ry6UBmAANAVaeP0Hlm7mPJKRv3SiVxDpq
mQ1xoY3Fw46m9RD0yOuzE8QEzztd1JKT4TuYAqW/E1oC6erZKJj/0YUBrWviBi9fP1IarQtLWAlS
ldgt0chpqyktPfUFcgaoMqW6fIqnQcNRakbPw0TyMzzsGqKDwctP4RuPkEDysjagObHka4iT3wC2
VGdk3tR+pcrdafPyzXsXxqr/YqYyxC85zAvp9entJI2lV4zXNY7rBAjga9j2V/cKJjKWcBegI3ly
huJzOS3BQYCMZd2D5ql/gsdxYhWYKvcSnn2rchM3HfVQaTgy+kacjAPDM2Qteqg06h2QGsbrdD3D
qtC0jkb60kgwUvoqxYPLWt77ZjLhqW5PvZH8RuNizBfoAtKQySuWij1AUigczJIXkKySfyF7wKi1
R1BH9cW7BAJvEkfNOH4lpYcMKW9hAk3bF6Se8gP39ia1npaVw3nviROXGRlX7UjcDS5T2gZ/Cc6O
JpNtQLGLdhl2pMoF8XpmKiPNbsqfm/1Fln1XzuL8p9QOtIhLxyK7M3eN1Gh4ehH3xfrPdemoSDRr
I0LawZQHFiJR6uLDSZdt82rlMCONuyWYh2IfHFEI6Na+A2IBoSItJ7mgyJCaUwXgMRi3DtEgnmFk
1TArTdfODYw/MZs49aICa5Na1D8Zzc0vTtiRjJOQaoWIPhqrMICux8JKeo1i/U06tupy5jvBnXtk
EgYrrE4SGWKshl4PAnZa5pNdXJgtcCK+HRnejjuOwurIZpbtL9uPWIKAnQ91IKoQ574LaReDvdt1
Q9ajnTapwCVY1Q36vEIU7CGwZqSSLp3Hy8QTaHU3zu8nB0LrFaeQAkcWkykrCDu1ADFQJ1pen1WS
xr+GWAHZ1jwFurInCKuA306AMLZwvvL4oIpi19en3J4kmWG+I4nEbi6PRiNUtxt54s8dWR/G0JUI
GZfnRftQVDbw9OgdQmnQcSAqY/QwxNDuZ+HVt2IxCtMEmZpbodvTbuDabBbVQerGGcxfkUzh8lUI
JPHwZ1tOZYMwUKdArSVzmHrXOCDESBUh/ShQpj4Xhp6LIwSqdkUFkBi8tu5jwFdLvjXkQSd6+Pwn
Nw0trBkK680h+RE4Ponic8RMo9GnO4Angc9VTb64VSjx3SfcyX3l5cPedV/b1yllTmjRjs7u4uDy
7PyYcZwNlhWTZF5btbVYcF3btCNc97TalmyETCYhgAjh5m+vemy2uu6dhqawEIWXscTA5KwQmCS6
4eoMkV/hIBv/UPU1acedzLCFyUohc0SH4aDqbh+iKNac6Crc93BG09x8iPOoHMe5bh/eZM4qAJTa
IGIHIe1GXuNACVCgf/jJAUJvIMnC25hXNhpDRXyrPZhXsTeV+y7BeiAsoUbZtnIvCSq547sA9B0A
giP/xN918lKQ5pWeAtntYs/pAxXPPuLrzv7QpcFnJopk2+VIQ9Elm34yr+dx0qbjUyv9bVL7vIXa
moQdFUcVc7aNhGk5hetEonPe1Vnb9E6ejZEzh3JG4Ucg2jI0/7u826jlOGyOqhMaqBAw0szhbp2I
boDBvaWcDLAd+Wr6X5zYevfx/kjqsAfVOSKdV+fWZ5jHfknGgwtagMaYA8+pfDWqmNhdovaIroMx
WACKy07hjK58hTMu3VtQl7vH2LnAVDckstVNFU8ggkiy2PlPfB/iediCC+Z7+H76qoWlUO0Hg/wi
rsUB3ib0JDrOr2odGdT2ouk++JmEZOAFGWky+xyCJJJIkP9p9xeWtXwOp9JrNZ45J0+Rj+CVAhQX
0Yv1XnlzzNqX4CCxwpui/TrnZsm/YSkUaXYZ8/g4ucHOKasb2Bdqx9c8x9KCWY2xgx6+QQr1WSzS
rjDCqUJM54VDVsoxrghoyhdMmUcqOCy2FPITQy84VYJ8JbHR0ODh/8ajn22OZSE277v91jXCj8vi
10DEOQmaURmgHXYCZgM9OdaTF+lOiHNfKeaUYZ3tFcQdnp1fdt3mXyXYL7PtKZHZdzN9xy+EdAdf
R6/EzDEQ+0q5ePcwX0lUSEiCzdOBNQaRbugnAiKAXjIgRW4WgLMwEh+H90muYxoUUqemNSZ55Vi0
9SLVUq7UJUsk28X/gI3HCVGIrkcQjzCJPkQgUbUxwuHc/Fn4xDgXyP+R3p2oSjDCyXKaYTGw9eie
ACdcDvpmq4ZwERf+WMbbpR68uDnwEfXXl1Q6L+BqWBaGTvqrM5enJC1cYaRBWITiA2/77Bi2Mlh5
pNAFO/INymu6e53ShWG/C+HdjSZ9VUcbFByfP28YlDZpsE44sW7VNrq3/0tBajlD+J0rtqqIvVoW
UB2jzqF0ipCBg6kF55SVj+q+T3rYuW9Cv4au3b3XcTc5GGU/mK0arPBL2PZM4sWDeGrTvUetJChN
iVl4AmFJbhJ0zT9VoH+RPcgyiNOM8L8VMTe/tfghGZXTwqW1RL6AzuB7puALWpZvOPdHCZXe8zlJ
iCAu3FnTC44sp/gTIgjvZ6MQlP6vvD0T2u37ndjTb8SQSme3jTDukEmIGCEBBDbLaAbqozC+LPko
GRQInXG6vJYIsY4OgFXDlchrwr9iVFHIMHIcABSJfbyFF8REVofHPveC3l2n4oXisBJanqEqJVIW
s/z92EcL0HSsC/qqd96HRhEHVQbM7TUoLOcAdn4xkh0Jm773kgWBulBOKf/vjZnBjJxqAXxq7nFt
g9CDlftvdVNDZwXGJ07WRJ6mxJCmoyihxBlQfML+YU2oxoTbmnDLF98iJWoG5/moCjMoKWq32k1Y
Lq+iUkhY6llH3D93F1crebvtvgexeW7rzIrDrlytceIoP4ZPG2/L/2dOIhWjHnY+29ekvJEBRSXx
d7AEv/D9V0xuOtH0M13AIzby0nhHmJlyvjRXtAUfDr1IJVfpdfD6ico2Buu3LSx2chvFXXmOVbTD
lI8spzJHGHsK6pdlVGQvTLKsYHt/6RDyxyWvlhNBAlo5f4z+vw5J3tCiD4M4USIzGyi+9GZwt6Kj
ccU9p5OKprw2wzzb7dudN/OR9EySA01c5VR/oqsLsjpVN/YxF/K900aVoO/5f9Jv8fg2W6++V9MC
AQtIzG2XazGkXTOil9fHMTJq8MymeSCSnhmR1UnM9V0t3E/h6uMpp9ZbCONEia8pEC10iE6XfU1k
2vOhvAJAFzUXVSrpV/JI7p5U5BezAb9BbeIf5OXdZPdBP1re+EZ2jLfqataua28zmz+DJ3aOUIa2
DN2O1skORRoJs1Qp0r1jawrmSXFb4hlxRnRnUK8TVucan/Aq4tHLcsfxwcsvO6DYEse4N9XvHF1k
Zybi/TDPzgEvAimaqkcA2RPlTMCHl5wGokZrN8IzTwYOOSSXkIBPYJkdPWqUeOm6CEtKqxNaeMOV
dxwed72r7hZ98xBAAj5vJqBXgymgKL9+EQgDwULxtCebHVsN+qfJDw0BE/ezKG+O4oE5/LCj8YVs
m8rM8VbqcaMs+MKZDwC5GBGDufuElwE+vWpfqTxjmi54btPf3v1sbNVs3IgrLMDdHntt7wa4wBVX
E1AC0FO4aC1hI7CsXfYIHGi/MwDELeGqtaM2R5NF6Tb0h5h6NtwDOY5nfSMRFlpgY4siptZ+x7fF
Ed8+Q5F48uFE1BSFN5FRJBjEs7y1TeSxBn1fYFukpEd8iVjlyzEoCPju6Xrhmdjpx4fYX3HNPiiZ
w2jiZS09zpCz4F7lWi4atppWxFsvG0adSUyRfQ9h4tIsWrB/d52vSrK1LQ6dlG7vklsE5CkJ6fm1
JlOWvFfhRCy/UdP8EpxHyTVCsZ8kVF52VZeQJ3KWiheEkpNLGWXuBgpdOX5nQ0xRjUes2sxsqrDY
+wzDF7yOQnYzGXFbTYBm/lTqnvgW5GVqLpT9GcB0NZSdflDxpmiV5zpIgfmk0dNykVzjwc+IfxkL
j4FDmjDWOZwZTLGJvjg+2yYH/VevsEQ/Dzd4f8+4mzyvTpMZV2EC1j94ITBgDgoPIgc2Qag3OSt1
KthoDvZ+EHVZxu6l/Pac/YFoBqQZ8flX1FCJzjA/LAQFvNa6tPRpF6uz5mxTCP+N6Cs6y2YlEs1K
U1S8ywq8mCyKux0OcHQseZm4udRRgyUSOttND1oHqeohlZzNImtnEAeDksyAauBY2E5ClySqatYl
aPlRE8mN0eTda4RB5A/cHsqfXDve6AL6ISbX3q4GAKUgS9Dsh2vm/LM8bez5u3/MCOROTK/ANqAc
hch1ca4cw2Ib4FGRYKSlUFb0V2Z9lgVI3xdDmuTYHgi5jLfUcutrBDfDFMM9jKtiVnUouyk8Fbbn
mTyuBRVnJxkvWB5KsaBYHc+LEluhEVxL+I2wOVe8djY01dlI/ib7iNlPNO7kH3QOzc8F5iSmzKBo
HDltebvH57lRRk0Rq0aVS59eSfvzErdCb7J0TllxQIQcQqnULRK3MQjpDlgOAfz0QEEeNUkk+E9r
1JQMaBWjH+V9KSZ4lGLorFIt/rkBjiJ9/Yc7xGe1UHcnKhHNUXUeMt4cHOVHor/RYCdS1jKdydl9
OjQwRjpjr5opwghCaB1de8PjzpOUpfglIFWadQVW3SrLoNudJUw8zwpF2SOdHaxBO0EwMPaP+t6a
9dsx3RPYXb7OMTmRFO9qrDYZhNcaTfxdaQCKIPOSlU+V9I1iuySEo8CTi1QJ6kET3MBNBTCMAn/I
I0GxLnaZLPsSrBZEkgDdAJ0qyru3lvGIfoUb/HMfPTPJAo4ZT1AtPndpHv3KPjO0Od2/uRSkaJ4x
OsVAlliw1eUHNdFmdgNTeeUqCdW2qlbT0SEUTlMw27ngHG2xMzzRDmh083t/Rwk+XJjY+q6XftvS
n1J8Kxkb5RXSnv/YL6XZy4PJ7Vfj52elWE1dxS1FMhDROtgWncGHrHx7isu+isL9+00DARTxNVeE
GAvminiEvevsBPTuGxJki9sa/6Uike59otBLhSt6AAnDjTwlG39EqotUV6MRoOrmIeflJaSJmz/J
awOikVg/FQnh0bD623eoKOxXM96MWzyZujAUL85pWmUWFvpl2DLGt+25g5QBGX/hsAM+3MNJ9bWk
8lvNaRs5I6FGM3sf72zNhHgCEG/RwRVm/a7pyiv8HEP6m7x+3i/S1rwV5/8i9umgk2jBzdyV+srl
kjoMzUsgOWVS59UzGuZmIQaN6I1komzPp0FMp/1j93NMkTJwUG/TQf1bM6kseRGDD7cT3zEbJIMU
v8SWv8UIBO+vUMPKkyl8Pxgnu8AK0iyME5A20RtQWPpe5DG6xQtDX+ewfgAK7wbWFMGA47ISJ27s
dUoyk8x0Xo/B8s+/Av8MZLvO+xZDLUbandvqtU31MCULJixFjuNqM895v7qLGdw/4Ml0KVWl0lQM
k0Y+EXQeaQdSqFXkb88RpD+QeN93tvqTYfzPx9U6EIZx1j5f3ViTN+mMnVvBsBkqPT+c/6NGnT7B
eTCLshzJ6Odnl5ppnCQrF8iN35Y1zb3p9s27bhneAvzokpgDNHRv9uSHdevF5oRsMDwAzsnGQQ5c
E08gS3KE889JkrwsJhkfhvIOw2IreNiwOBgEC96gBHlBO1IeIdiQ23AHeM5CtWjPw4CZibX5Snvg
IInKgQ2bThSxlfXODk6FX2PmD7Oed3Xx3q4DBB7VI4T9NffibHaMcqix3Ha6476ea0zrHABU9CBD
Wlw+CU0AFyNrh3b1ZH+NLJondS3e2AWd/GVtSra3/YJhnydMk0cboI3hjlfN9bTfHkHb26bKfitZ
7faTOOgJX/zYP94Lr5wSsZu9wbAIESbKjVYP/m6u3bpj0u+BL383CTE+MDmkFy7GJZWiZrrVcPdr
MpbXxUd0lcaFttU7/stSCjOmVT0i2ZvVDEpSlo2osJSKS6TihmWoMxXjwzal/adp86qk2VofiuVJ
Z3wnHxtk5xPT28j92HjztoYg9sARWS+WPDMl4W5IL6pc+JGHroHlIzYfIahoIgnLurkO+Js5q1z1
G/INfspgK7gXZgy6TZxRFHfqfD6wjfi4IOKRq7jk4mbpjKx3Syf6IGuJiPM8zMi4+T5gfSAjIork
9ZvloNTWurWefon8qubLxZYE0V1KUdcKCEINBiHOU8VUfH6rFFjaAGJ+YNbqBila4+vjZpTqAoxn
mUeiHlvHIKB0BarwqsfwK/ShEFi2ETdG9Bczgq/pRe8XX7kY2sXXn13NzMmqxFONj+NxkKFk/JLF
sKslvQ414+Eu/4bSxY5D7WDRtXegim2jopFwkOLxJZ1MOyBx/ckVBIGQgy/Wj51wYtRJt37YRAzZ
s4qkIBEH0/a4EsDGSMqD/6ncF3LEonKsaije/wyILK97s7MUdnvWfWstpTkU59DLmMdDLWfJTXRr
9cml2HKF0TIDhNG6Hf9AtXdZSAsWwW3H+zbgZUxd4UEVFD0V8y7k/vD+DdMrEP0RkE7MeSB0N2nS
5sMV/5kHyICdta4yMnbmUT84XsJxXZgpCDMqNFl6A6CQ6iGUVeczZ5oA8/pDo7EtrWaNjODVWvX/
DebBFjG3txQEpDKpna2H+KFUVnJaYcmnaBms1G0x6gEe8YJD0RGimopTTnAAA6u1GYtwh5yG/fmE
v5ETH+jAtaEW5k+vY/b9Rg8fPruvN0qVgAsLq2jdM9z2gWmzt2144p+IkWzUZC+I0ykCkeHXaD6N
Yi1QkDgp9zkis9hAfHtetqNwB2cL59a3ufhF42b8Ra9NchE83eMJulntoRhOLNUmPumS6WdEe8GY
vGw45oU81ArfRDMcB7XT7S1Vcrvq1LK/mtNSdrsMUAVyJqLlZ3fzIKQ0t6c1CCFB6L4eqNObxWWx
w4z8vFJUkipaUL8t7LPfgq7VY5xhMauGJyMHRWATzcojigF1hNHt4k/7h2mIEuFxbYiX6fouOk0g
78vz5tWdniIVOiH6hp34lslvwDFhJhaMrWeaC1uRnfug1o5FIKyV5sp1MsW337uJe0s8qANdF9Z7
LSIQENOOwkx9RSEzhYQ+VB/oSTZOHsNs0mHKkruK46u+M2l11XSnLTor2Zj63iNSTvbha72ohlB9
ZymHekVrs78sbe/HUoktYGcq7CrFNYEzBwd76B3dpgvQC+2JJz08so1xg1QmesO11AM05tNkFzrU
x/z2lqSy3ZuJCNBqJJriaP//ec3CecDL9568STB2sFH4nuVfEUTcZRItGAcMlkwjpUATHGi8MORW
Co4FgHy6Wo0DpHzyRJPevey35LFPP91yexetgxyV/0hlUbdlUV43U9duCWnx7z+gzCnJUbf/8PCm
LGou1iz0RTe6GF79DVVEwmXo6QKEtcZ65D0qF2dnKGcg7tOgYoThDtBdvaU08rWqwFTpSfa9o1Qb
ha6ISdgVXzBjFVA/wljyHzhiv/kJuKsN+Hx3luS1Zb6VheYL7w0lBFc+60ptpwINqf1pDTbwvm0W
rI+pLAx5fujvcSdNtWH9BhE/BZP3wBQzEJg9+NGQFKrJgnlmkgawvwn8jxZKb9O6k2/LqDDI1es5
mXE45fIL0dPBRJH3cDKQgTZZ9HN4eUhQi1Wb4ABg4E4mOUM90vbUpHBp8R5kp9z0+/v00IzoTMvI
JBEKDsJiWP/xP3pfoIdYlU0Sbc19giziMfNZBK8txdMjDxdGYB8Okuj2ZPZH9tIUBh2md6Q6NM1A
WTGDWjCVv29c7ZLmTW3FHAh+4Hy6CnehHksmWj7Xa/qvX+7JK6MjaPauNiUktObDZ/lnDkc9uxNS
fylKEfwH0Vs1UrxoweTSTbJpSxYQaU1rXrN6pU95AxmztknXcoGjZ8prwFgrwoXmTQ0uVqSSoxtU
/SwbajzX+OMo15BbQZKEQFbiwhbIhY6c/VW95PZZA5qjbVnz4ItAJHk8mcZD9rYpe+e0gSes5AT/
RfvG3xA6VhF1gFwRHtAGPArS4FWObxFuk/FZLGfxkbFmTIaTrYvvF0qOs5l6prpjYOBsTEcPrj3d
tAGw7Ozne4mlTs885R/pYH9dyl/dj8mlpJJnIeA+AJauGjed4dC14rq0s01Cls7uQJYGENHwcz3p
xG3PrbzsAaXn6cN7UrmHHtp3B6MasD/6vKzxzMvmHVKHtHlMyJrTkZE0iL98nJgFCqnPowAGThMz
KBeW5TMw9vhrC08EgYe14We0wBp3OUC9GrCbwMmWOFQAVZZD/JftJbepEuXOABj4/H8u1Q41BulC
zVxFsRyiJo4x3YHMH8wKVYErIMJ8v4flbeMLf5rlFZHjPFbFQvaNUS++kx0KJ5Sh4EOvmt6DIs+O
+qoBUVLN7GNEKSupjrdTD2hdQj+t53WX3g4gCpAK1Gs+/AGGhaPCDS7E9Wu3zT8UVylhBjgHGo1i
PD4U5O1CkOKwV2tx8NWHGexrt4xQDDoZvfYd/hxZsh7LC7g+0cgf88QTB1G+mmC5s4tLADQ9RGR/
ZRiCCwWhIKkdoyCL7thbFWZkTI0UAo/qAOeBxhgzfVNuvsAATa9/0ZTH05x6dcbnyKXMwwm2tyEI
ErFs277N7f5S7AQb89+5o4v+GegnzSwOHwxTIaJ2z3JuJ98rn+6xs+ftSfRQkOFfoXkb3xBK+Rm7
zpACaZHUtUoQy4U0qcvF1gaAtGFhAC0h+jVBgRlCArE+BauaLAPYVZmN92Mo+UDcbdODCZzLrlN7
oMYfZAMWFhU8kpmQyKNYnc6Jx55cKb13eJwnKmV5awkHTW30nzPKhyr89phD9INpb6Js7FJ3D8yy
2BSPJ2HUiq55XsF5WAYYwS04lyVg3L5kA+Knw+cBGhGkEMfYhGOcSxDJ9ypGPoxGADp8ykXjjvh3
FHiYEWDCiNXkCtQeDEZ5qSC9sMwLuGZRBuZsuvUOd0vELytO7W/SNWLwa/DHBEnlmb7VLWh7hu7v
ZG7v9S9rwLtaoxYe0YY5fUGSdm5+xx7RkJ1sranAEI1LqFuSGtPv7TD2D21cJnEok1wzvAKo+EOt
KuZ7ayaf06N8Vi+73fXpRWplpX8c/s+iTmwv1nIVjFUL+ACCThdPdI/8lT+mSheId98kClizPKV+
rURhAFEAL++OaSm1cMh9tvkhvyuvHeg2vsRhoHx8ls3ydnzqwOHDrIzuGy3wgC2bBtFNLeQYz1O4
uYymsF4myd4kPTB5CDmcS/xsMn6+IDT/qyoNXEGa+cbr7SA4s2GcaEE3u6m6dONfDY9rgiIIUQ9l
uAg+aO+jjxevMSsj+Yu5uYmqDNgmRTVqJHku2UpnBZLVJnBIHrZ4j7MrhES3qIyC+b+g9PT7YFer
JzePbxQAr9pzet1TX1vWUli+URkoz1DYoAfB+40E74Xq6nuO1a6YxQxduioSVo7qH1VV+Mute4ug
lfyQXtWXlYpk+UHPTj10yuDJCL2VQyhCZeZLhC1iL6/5fUseDId1cTjggR0EUT8JejpKWVAcVaTd
w/oIUiJXkS9zmA/9+X32qiBcx8Iqh3YUBUcPs84X7K+CYICw8FPwQMlinp6nW6ptk38TeWIG9haB
VVSBPBuQayZ+oAmSRMzugB/3HfpEIf6eCsjWIQU+9Jze+N9+ZvGpjqEoM/cDfARfar4fZdmLbde9
6laxTOdXMZXAgZXZwq9pShzThNCPVYCzRbXGJ7J6iS6zZFCZmPpTIc4h28fpM/qLHwPWcr72ixev
Z9Dqk5UzGVcbOsIkIjEFUedw+74tXgAz9Popc6CuwB8EOG+fKA9olOApd4PWIaoRMYgRBPhYsq/N
08+HuFupwscUrmM58N3jA3UGm//+/nNxpG0F9DQahYQQqV9juQLA2IkqS0QubVON0FeavSVRkOl7
ThfiUM0qfN+Ms1GF/1uJQvrOzLu6YfkEmqWLhUal/4JkDGYEw7fVco0mC4GObp/9/J7TnKiiatDS
Yb6m0JHuW0puehBgSF9EESftznh6fMkBv1Xzi+L8OwrceRuC/TBcus4VDJ0i7sVCMSRko97yY8Uw
V09MWNbW/NeG3mdyMYjFpm0q/0HnIy/cM2PdEJ/6DeIRxdUPFrmbO2YgQVGd+IZ2wgCsyZaB2BO1
3WBYFY2DMLAQcMqoMQtK8tiEZk0D/XPpPoqdY9JdYi9si5FtCtKu41o5e2VPhViJiYHXsY0snx/F
plgHEolCkSO2OrDMS99naZSTZ8JcR+QWrwoo2JBeFSwRlkSwmlTbQuXucXG9KVMQbFokTtgLhPB2
k3CA/OkAqDEKIcN56CH+eqaLbn7Rz6NQgqFGEFFo+9NoNQNdOX7zaaRAuVAltlLvHOmChjFJy3yX
CIRXhV9URmfAS+ztTX0GvFXnhY2zgkBOyspgtPmd+73/N6oj8gxJPSEnCEdPYP8Gb8rLVpHSL3RU
NsI4v1Xb3KUu2NDZn93h3hHE9qbly0uW4B+YBGWL+0c6Wu13SgjZrJnwgQEUuE3nQlRMAFgH9/T2
mNsq104xoUDKSfhOhJwcKqDbWh7TMf9DHerxai3X8eDiR2CIbnepI66agZXZPNsqF/fu1t6DDmhp
wDu2fAGNyG0E/Wg/BhDhfwf3wE+SqE9DwVpt5F67rt6dZbh9VqOfd+XB1ELJViVsf339lPjGWoMc
5wxf1+MbfNjfu3k/rkTq5oPzef8xqbEHGKIUb1mfjwFhuKMFwk8J8mtcaxeXEUXPVrwCPh15cu5N
aJjRm4eRsfgTYOO1JXLPtK088qqQNBdBDaaR/5uKHEAw7KdjZfhLy+N+Y4xQ+kfr1alm94rOI9uQ
MF7aiNDSDDVtQy0QXgTgwvqOYDsRElpwz+wrI7v+Mu5qQFG8Sm441c/m+PV6WKjxep9csJl+Ktib
QrzbziL0CLXfdz4LNblyOjos5JcilMs/cVGjEWfPsGcYmnlwLSdoZgslhZod4Onkoo8uuUPEgeGz
LgmHfiob5BE3p8vc5q2x0rVWoNwxM/0nAE7uGApMexiaQef3XGKIUBzSDisnxyatJs6VCgjyavnn
g2csjmK8HIOY8d3JBColvrVGXm6IeM+n/4M5ox9l24c7suz4jho9MruylGFex3FtlLndfkkwjIZZ
icjTaUDs6JnMsoWaK60HVk23WWYQ3A3Lc21nB6VQoJJlvUPPMR7hLQb3zh1QpnU89tBqIqminbEv
Jp6j99mMBPid2T9pWJDWUhm1+G8uMQyv3szPv9mBZeWwRRp1eMr26Kok2cpxxKfMiXXGEzlOC5aY
EeBmwHavnUYbaPrASicZaKs2GHE4P6NNyOgIUs79N0N9nro93nywph7drQV+DR6Q4AXM+qpX/EZD
zEfjsjd8cqEAmRH7ycbFvhGId2ig9tAcpq6tGx5NE6dMBRzA2lxwNja9XyF2bRi7rR3k8DWHzUPx
gytn23+lE4S+dz4wJMhE2kbnAilZ71seG2pdqq379+3vOftzSFKnEbY17a9s9Lr++lbrJBVkvwl/
6Dznrih4iQuWx8GRl7YHtxADcbEabsiaaEdAHM4R2vcYrKjMIJk7YGngutOTSBLKcIYY0PF55pLu
InCQ6eG6SnTe5HWoEc8q74IEvgS2OAJKBmwDjo/86A0cstO5jg/3uF//ZdpCIVebzh2Ou1DoAlEa
Uv1yg8QCuZq5/TdugrHUmLFAMO5G5ogGXJEpEC05Uoi2SKyKEGMcmagxFjSW9D1Vs3gmyT6Uh9Dp
fo6uHjj72FmA6sgZ+eRzPb0E6AgKmBLYKnvooycv/jLINAHimqgJeDVrS4LePqD8TgEslJjel0NM
6j9GWUR6rsofV3ztes4VOoxmkC+ITp+INMjeU3pa4NYCvcfMrAKmvMElu7NIQ5ZnQ5FSh+8no5N6
M8wPTAITWJa6qi2NQVwJMpHCZXHz41CygZ3sOiSMIS1H7GJ5zUJTaapjIeZr0VsmNcCJGFpvuuwn
wxSjui8P7ym8bgmLciWJuL/Df2Foi2RFKflPBjMqvHLyZAeeviQZ4QlCKgzu6LWW9XXBfD51TGqU
1zZLoqdpaHOLa512jtKFApUJ4FQBfGHM+4NMXvgAYQkUWLqZYHxU6oT1Dr5WeHQXewCbZAKvNRpv
IjTmUzzhp1CDfbyXfznwslCbX+eFP+8U2uTjxn7AQIWztjSgB7yI06yqr8Aqv30U75wCNdhNJan8
sNHeyj208097UHTrYp2m57P3i1ULw3INaIlSX8OQbMiTSZsDZVYRp9boLt8oxEDXrD4KaVmn7DyJ
2OpKzYwY4OsdXDXPQuKf+enmX8RnPAF3lJIUdHPojRrilLFNPJZuqzMRPA+cQIK6l1Qiezp661MZ
bojIBXIt4BWkCWtxosxPQSnbE8uFKsH9gwzpY46EHKxHBRZkc0BjYD8JzpxxI8oie9kPXDenG86T
HXwkxKZmmbzdiLlSTOaAdEqvKNzr/aWopmpfvcVD+wvJKk9ycVXB6PJsLnYSssvTh2dyx0iTmX/a
/aMywByLF9Q1ZeAFx72RTK1FXOSbZUfzOkCOFu3dvqRg8rnXozFoJlen6MEDXIrLTRGnsMeLIOEd
UKnY1AdDGxHTp68N4/ic0iDZzNvqATggRFYcB9PUsLQ6do0M7a+YwOrPSb3AxMjEYvO8H4Tcdy+1
ZvVX00FqWBL/WGZF5x7jhgd74dvt1uzRKTLAkuBtkXSwNVR3o9tZACa+X2Mti4ofba9cU/44oayJ
VQ8JG9y+zqrPevCVtlJM34j+d/iE7CZQZeIEKMaDDbMWie9Bh1AxVo62Zi/3viLioZroZsq74EAp
hW6FHiuTkDp7bnYkNobFWM7f3EfvSWSmuMWExiBzO8Qg024hUNGcCPw9HYH9tmdpqSyQIKW1NFAv
wkDPd2pZJnIcXy+DdApTtbbEBZZiZYQqavV+HyvDEVsEETR0y0qpxir/qp4B5H686FQHu3S1O1c5
mpwvFzHbqmwAzhOsGGoah+9Nnyzf75BtUOJMCoKU7jZ1hUualpMkpEeFH6r73e+RCXf8YjiaP8mG
qpS+QuIXDXivzZ8/zCuaNjERRzY8yhVs7IpB5+YcwM+1AoIXIfSF0Wd3PIfAeSzgLmgb2y7vsyda
M3lAw4IVp5XeMOu2jzxeodKuQVY+1lhBOZkIRpWKAu6PG2+CllE6tvCwcBO33y77CYaghZ/wsQN1
6VGTxfkA4IIba3NlKizO0Z6NCqCb2aMbig1pc/12wcmx7rXVBnlLTnfZUSb2INQeDD91l/ybwBXl
lO4u0PHdw3Btxy5SJfuLgzsQqcQNZU6IvNt8sIo+YzpiNoIPlWxGdajDBNXelNrjK4YyvTWcob44
VxBhdQH54pa4T38KHcz+3i3anlNBpoh02Z13639JdYSAuAf6MDPVgpqbFOPzx9AKVUVMnuprvUHr
XTM0rrEAE1z9lf52XupGcX/Szm+jfA80gDWEFvNr2cnYXn6YMVCtQqO8lw87rmMjqkV7WPO6j3Om
3JSevZdr2C7T+az0WCaw0kP4dKP+sVosJuv5jKGUJrS0ci5RjRPnuJ15jltFsdUtJFyn0DlG21G/
YJB5Myp1ZFFw0gGQzlHfQhvAtDx8pdBAQjeNfUEqU7PCqrkpHkAT+WIFJd940zhIws27wNx4KEq+
ZjmSTfjfxOpsTXBBj5Mgc++s4cXBhs3a6/xKe3DhbswIdbsywW7uno+0GJY5qW5UXo3+H4N724ba
HmnL0HWUQAk3xd6Dyisn1L0xZ9+/+Tm3ZCy6FxtTsksxKwTkuY4kQTWwRMFHtHjKucBvXDKkoQJB
z+X2vCwFwBIwxeHszWfTTnLZChoLByv9Rtc7n/HgCHzadtzmPKSWKfYBmAzNV5ceyH6EOl1Sk8Mh
HpEVWRblab53HMeJd2gDrZoqsJmK1QYJLjYNlaAQZCEaXQtyq7pnbsnqKZE6GrMuqDwwNVTgHrY6
gHludpm8RYdj6JFzvPo+J7TM81ZHV7ytnRgZ9XXK9xBLBNM5ZUbTe4UkrpUuZToe8McqyaucGzvo
0SJRUbeVI47S0eFSP/etsgbxpENOajDnvRCQSNUELsXi2iTcqITHTjA1rht/LtqBONwp9KjIwlzV
+RxIKtOahUwfj4/MESRbRxOf0lgOQTsuDJ0Gw18O4x8jtMB3Od8di2bb9BxhKJqEkW5uCX0c8noa
k9pXDy+QaiRbSyyx9LE36QG6Cq0xusuNZB3XL33aKsV5ztMe+Kl8Re0a3zBgQBCKpTX83LK3c6OV
e6YSWikbZMPbczPUM/pqbrbZsO4PKIeHEuvHaEjR1rSBQAYsjwXm14/k+EZr6iQTX1IcacOeU5MU
2ZGMMfcbFqY+5aafqILpPWSCKIX9kDwgC8greK18thNEXe45PFUoI9JSO8Z/f/xmvJehPa5yneB4
0qE8hc88W7SbkBjS/oZAOp/s70bESMwJvfSwRxZ+koztm3oZd9I5fyC3VCPRH67r1jnBNvO9gHSP
Je/lEKl5VJMXPwBX3D4G1XyAwpVQNjTW9F88gR9yVJL1ucmu965ii2G00aHHlDSsrzq0dVFjCIMS
9yqyfuEuecI3fVk5VfTBRXSdTllv/R+8tpd+oKiSiMaRK78Qafch5ZIJYFu+5Q6/uvB2OP0PYZPW
BR9fnabDJKZTfHTVrDl+Y5Lz0a9T0Xztp+ZgjtUw9wkxrNr9PNNmQ87/NYh9VD6lTQXX+b6wI8rW
Uj2lp78BzvvzBTkhDgearnt0CQIC4mB4zFKVD3+Y7/2Ty5TPlGFRajsf+7/zrd79G/VjDjnwdfvr
i5N+8qBkQsii3kg6IH+xnTsb/ymVM9TOsn8XyjJO6eOHJxbBWP5ARFT7hhoE05OK45EZ3nRJXwme
7kF5ZfC2i6kY+PerOBTZZYx6NYA9whF35vvxkIXBcMhmfk+Esa/c5NIODF+faj6mAyuqqoEWJFke
pzDbLJ6C8CIBy8tmMRVhPXLr1kAJm9oZIrlvqo7PfTjTZWLHwqPxaFHyq3hoEB1bFToXDvxEKwL0
GlBYfrym3FZYgHlulXeHHtzr9sVLIkzf5E83Gw4iyzleNNSX7NbeucRjRRLjo0r3o+h9B8d/U5x2
kwSBT36kQcF5zR2iWX0PoGSZiktFfOg+IfuaNM52hqyyCINdEI6kTzGPIr4XPeyfEL47TTDr25+q
7zC7XSHQu/YRCVw0zKOj4pipmg4x6wItG2AHfIimpemRR+njUSNmtG4Vu8k9yRA+YJF2ycuv7xWD
Jq+RfcG4L+0YS7PmfiAtrZPUQ3L7fM/NE4FENqEsv3bCtzUtliuEp9s4UIdPbMygdFknwb+bU6qu
fop+xDKXCJo3T6GP3KmZNkjlQFNVEra8dGb6Jsvp086oEHCz0o46Y95lLwoq3J0jC1UMb8LGIU27
s8iYrb1BqKKPHDUdMisoX5Fiz9Sd8YsCCa3BJawPQQY5LrIOxY47VzBJy9FSeaBjyWlESpY8cKhw
2m/inZyhMuxK4d8ZAw4Bn2cMkAJpe19Wie88czMp44GaEQGj3riWdV67NoY0V+pd6MCZkjWw2nww
X3FDEhOGIov/A7Qhd7sSuRs7UYQHSg30lHt91s6+e2hlG6nqAroItnCzHqATZowSBMYnO1MSz9Aq
JVgjbn94aTpSrM3UF2jSWElr2Xgccv9A1FXGd8mFp70J99NV+ATnOaQLJHgoBtp7xiMkoarGAtD2
4V8wV9c6LXecZNUnSx532h+MaXpSBhLaXob2K5PXFatBqsF2gig9uys+rbp21FFJ0SkBCDnLI8+0
SKThn1EmpX50dPF6BSP5diajO0RqlOTAnE9lUE8j0xPN+AyM8p+onZdg4Q1VSFt2KVuLTcYjlFaK
hEy4AVB5k1MVjImu3JTX02hBJjVkt4SNwI2bCBqpjVxtJLKf8CYdItdjpkjN9kuoR2MVrzlDfNM/
el90D0ytO/7v2l4m5XrPxl0Cswvnii8+dHxqJxW9aGhCxpz/aEW43sgC8LE0B+oeP4pBOj6D2FN9
4pk+8BUHTWnGYi22jywUbLTAXzOZ+7E8jWDEMbT192OHX6T5R/sd2bjqR4f1sDYDueVOQfZywl+s
EcUdNm68aTa8jvYBy3YwJskxDQnjhH9bn4ywXLKtUoZu9gfOeTek22yjKHfo5y7VV7pv06QX7ol/
fYAH4/tF2DXXzzt400puF3I7pDrmzi4RwgZib43vfl2CygqkBE5PzUOwDUz/Jvy8++ur1EKO+W2w
YuEh8Vvxd15P+C4ai8FlS3l3YVXvcShO4doHE4vzAfg8g39YyaukIPI0hGWw7ocv2AMOxkjmIEZR
odlgRXIZNMk+eQOchc6yTUXVBmglrkuFSUucgq6+dvm/DQgDA5xSGLgAAIRJ8Q93hUq0gaL7boN7
nnwcHIvqN0PA4B4aJ2sxpsv8wETg+cJuKNg53eXhg9l0xp/9MmcNfqgJRhCtRaJT38CiazN3ELoi
ODbyNTBSOPjawos75LiGwlu788NDP36PzlvDtQh05BdZQL1Ee4DkTMyGQxfUu7k/wneI/1xYbP/J
bHRJUmLPc/cc98JO4Q8B4MFQXlhtEFPFmAdaeUeqADAF5d06UzCkStfYqIPF+ShMsXQTTQGCij4/
Zb13NCNDKWjzb4LMBlKcCCXNPAQL2EZUW1CFlUnXk44yvwiJjUXNyTb27XKneJyBSJkU7+k3CpS+
hjiO8cdehEN8jyYdTwjs0DnBL+LQJ8eFjmzybJNIZOOIsgULcO32L5mTnPh3+61OKRe1oMI7IUUb
P9QnDi2sCyp0aI9s8FeOlEohYwS+weR0WrzXEj6KkXWA3L9KUZ10wGMd0HCwmMRskmHwDBShwikL
zPmtwsiEf1Jgjq8eCWPN0MtxJ4jJyX4NI5ftP2tFcZ4i4t/Ti/PidI2Rfbhf3AxWdHB21tZO4fI4
DFCezfFerWz0YiYyTaD9RQMGS+zcGGf2De6nZ2t2sQQFsGH5qzS+uPmgGUIUrsNcmi4v1LaeJAR4
QKd/n1F4mdEcR9eU+By+HTufpkTbI1lg0+63uLxkYQ3C6jBb2G8MWlUa1kJma8WlaE6/6jNaXsZY
Ns3qwCtTp+5q0jGi5noJ6z7ya9XqFElyPU2dBoD4lWDYyive4I3KzO1DV7/RQTwXYXpV7LTR7Ud6
MAzs5OpouSPqwNWqAW2/drDepz83hdBbbl/bpXOWe4/4V6d1JMpUPqD3De8YFnzVHRmJ1g8/dei2
f7Rx8yK+cl/JaBXkoYNJ1ymxikOtoNSDPGUduCQDYrpNE5vOh/jtvcMjyV8LQPO2JUCUhbvM9sNl
DOxssO+YyaaMZvwPMqLNOzNrqvOkjyQqN3xT14ITs7/TC6PIMp4uXma0IxsOqvAjQ3n5pYchh2+2
UjSYWZqCA1/kXf1Vp4YNV4AOpFqFD8T5Z0ELpgB+759p6XQ5ROw8E0/YLJ7EUEEIia5O0nTtXcIP
67ysJKlkIButLGP+IWwkgeV2urD+jL8gsfqCikCjP8dBsAHfROLdl4RjcW/zABU3opk3jpr3AEh0
eITywGz6qLYxTRTsBa4l52X5j/c49LuiF1sNzq2NxshZ1ahSTnKZKU9QRs9Y4kzoy59r7/n2g1dy
e82zrK80HLmTmnEDRBTaQODC8pF1TxLtxtjEuiPuBprdYvI1zsQa/YQxi7USUkUF6MsHQ8WEr5hV
6IZUXXseH3IWqyOJzTRnhQ1zj7HphpgmpuTxDg4iaJgYnykkAs1snGlqZU9gzSBYFG+XiAUDp9OP
i8e5ZxLHip9s8lNCrPGcTJ99UkGvVKxWQtpw24PNWT78Nzz0cTGjlHt6OtpFys6IXfbQ7IExAsrW
XUeCX42wXTKM6RdKXFhOsCo12VoKNdMk8C5yCJbcg2FYYCTEDHmgSiuJTXFChlhDXAw8vmBEQam9
QA4PQpK8dIsgt6SRQPRlBTTds4mnGekpWCHv+Y4jWC/Vzo8+FQSWVTsScCXflUtnGzCwS+66D9V2
3vMm9lkmudyzg/AS77KF+Oponn2aYuGTu7oBI5Hn1x5NyNH6+zbA6OMXrpXn/J8nqFE09GRAwQLx
35pQ1kil/vP0qEm997csEI/cvZaA6tG3+v74x6/5PXHlcf5dN1LTcaETc+jF7L3U55OCe0NoVmJl
8roVIZWNHDf6X2IiTedhnHWAreeC1xuVDxz407sgh6wrG+eKxUajKYT3N9divqI5kuWJhrmzMEnI
QsO8OfSXDZylmViYBMTckXhIUJY6p/scA0UTCx+Ah9136xC8ZUtWs98Q7/qTPAtES+zVHLA60APQ
A0s9x+caVvQsEhpdBWJVnTXINgzHuS7QKdf27AJakJPHHJT4P5dPZzvQFdxiDDbqRolY/LPnuIM+
8cquuxPvSKkI9CDO1ykpDrNDDkzcPLZEXpsrR+Dnm1evuQXoF7rg9CjhsTBPhdbwyxXHO0OXhfsr
Tseh3yJMSUR1sBih+X1OSBE7TMYKsLOcs/xWDCTPIYAGxB2Y5cvferOzCov+ZYxfPdAnxMybusDe
wk2Lcx2nH92OK5S2KvGeqEFYQMfjQKnqHK35lhLsbVk5SHwzoMVmFvi6ykoxr5YSSknOrIB/uIUE
NR3diXl3TIGOlbogh1prgXJijXK4aqxABKCBTK27mIRmM9CIjIGbcFPBa0GtrrYEqSqONXivx4SM
wxZQn81hHSHoGD1AhcjFX4ovWLYhN9aadmz+vGJf8euprhUB+zWOqrm2cxoWmI5hkIQBwkRerSWs
vwpw2frBqyvhoLXZqI2rbj1hDFg+UQ1Z4e/jC3aTdXYRsCbSS1Nq4D2wUKoRxFdBd4+MawPlIxJH
vb4Tc00y79mMkzj0Ift1ABLaAkXqrhNFUGuur/oo/8/GELOJ1EGfZpsuxa6aDfGJBjiauOxFxvJF
RCJAKyIoFR9izSDt85tQNsepavZ6dF+Yo67g9eu/qFZvUkgjhmqZ7aaDeOBtWEi5w8W+onhGPy+H
UCrl67sctiedP6uqHhNTePJoJY/FbQhKPvDDNItU1j+UgSlDEbpold39Uu5BLRuW9NQFwN61qeZX
tsX76NGWf2ym7BWj/WTEIS/sTruOztoX9rBzEa1jYqPJcgOW4TjdbdUnRfzRszc6ugBTneITmc4h
dzCa4it4cmyXQPXprKZSMjVPPL5au2Uhdn+uV1huSnB7yfNJlha7y6HDHH+63vgNa+BPic6SItYu
uH3T0jOh9fU3MpjCgJkEY3/a3Nha45C+FefXmS4gK4zGEhwem5IXhWtUHZV1hjo8ti0gXSoG9+b2
55zB/gQNhIeE/IdgWWrrSO0/A/0H8QECwp+NQdW/0SCzzXvsI0wsm2FwkMBYtgsmvPKp9FilbflF
D18GGlY4jS9Sipycpab61LABEQh7hELl2g+r67P/1vAGDRB+CQ+D4IxrODeRsCm+ac9imZk9Copw
2ajmAvJkfs4LnxAO77L9yW/qbaMWDunr0z5SOKQMLhRzmAAY/WPk0JLbeztIsoSq4Ux5dEZgcmU5
hWd6LmbGzw+IAqje4YvUJqHHyVVpYfVHvFOeTFB8oSsassCWeXnQLwiLl8TordHYkIHDLFhCkYT3
VGiL6ee/VQtjt5VjEFChb6ag17yTZuqpdmkfdM/aI0F/PRPsQfhrvlAQ2oia09Mho5JU1bg5rMa2
CMhMKcDKtB6onTRjxrqLB3j3C+c+lHPX7oS0oFUQ5NKGrJWif/+5W2mogdjSkAh8sFPqhfwN34nn
lEe1cNeoBlNzgFP+aQSbL32fEd2blmu1+ApunMOjiJ+d1eazydRf9Vq6Dxya+zA8PLqQEn46ni6p
kN2Tp57+ClmFrZXdY06ZNazK9wPj+pc4R7/ZSibkrEzOUN479UDjCZneLtSjl2vpC8aMNG6+WJfe
IKgvdPanqVjkliSRYm1/qEbbEHc1BuGscC9/abeDFRg7pms3Hef6cnDiQ0tDig/bSn+acCPMBnLK
wf5KPKh3vavsLnYi9wPNBLySb+HYtMP0rnZl4ZHhZkchsvJbi302VA2+ZCR3wsYqVSXvQPaxf1z6
Bg9ol41XC4UW2y0GHCwsepzErQ2uhatkn+iNyLFOw4g1GCDkL3dfG/shJ2Qm643LWiUY5GEO6p9P
pftKbtyOhzAJfA5dHINbdJcRI5MHF9GjASJwkLGeXgB8VOol4qP7OgkfxUxoWeycRP0brWrAngZv
2Hyx02VSP7qW15R0HNwtfLuE+/2nSnCUy3zlU8uzv7cJvGceNNXixS6/dodxbNMu7sKjatMrOdp5
AWpXFVTGX9/miI3ZBnWPVbCejychfQodahztWDfzyQuFniLq+7OqvoDuRNPqAdxi07f55rnNLEdQ
hBWni4MEYjn0iSWRHRsUvZU6WrLc4t/rOrV/vEkZBsH/39M0HLiK+baBfm9fp+j79j4P+ULz/X1X
vyuecyDf492IRjmh/YEh/NRQZm/iJQwJyeHN3YCCbGfKTcyY/w4G0q19/ELTH2nDrQWNVfjVmh0X
IeDBtzAxvPbFD5l4t/JGzcClkzmPcXK52HVUfcNYP5lOtJ/s7uKOE0d8jhHQru2+XnfRmQ2CPC1t
Aex7cZd+kjnOwDrLz7KTdbav2sg9Zqudo550nD58YJ6Xe9WhYLCmIOXUQrAECarcFZ909gls1Iug
aLqKrwJOE8+xcPzSA3yI4UkrUn3QR9nUxj/C5prnW/ODuBtNaGQILEuFEXWK58+/bqE0TkPN13s7
GandT6vuWzHyBxIEnxAXY1/2LzMokozs1jwrl5gKhBmzeekRdpeWcCiRQyUr4HX9xt0BSO5TQMMG
b004XSpPyyhweKS/NtiwH3dGtos6M8vXuEykdH+UbH8MwEh5tE78jKlk/lm0qw6rqDW1457zlLeS
qsMitY1QQ/FuH5o0GJAZ0XM9l/BU8hAYmgAvyPfcQUMNtW4kkDnSioJ+ke5XO07TSki6cONex2AB
g/0Mpy3/vRfx5iYCDo2G1uza5iyt6a4ATpUJ2HCr1oRHMcUGAMqdq0rX0oBBZtSZm4m4JUHYQv48
PNh7UXCbSgcL7tt6Mcc9+y3+vyuQLlqYuYU4D+K31MWb/Tedn7KVHCd4qsDrVcFutcL5rqHTTjHh
LmLVa9/vsPtznc0BHm9bYUaxUhayUX6KK2Ov2T5J+UVbmbD3dNxPKcYtNM2ZsE4aeTozNZ84ot6P
YYT9A8dUNzPOO7U/WgLZLrbL4IWVzUa5St5+XaZkk6jYl4/VCZBeAOLjz6S72+AVBOhYx8dXTVV4
qG1BQ3XhABC03OwGxCEhowRU5vkn8yGaUb+Oa4HxZg31AlFp3sUhF4P+7YVyv28GsdF5Dk4RAipP
L6fJ2fxwL3usS6/99riPnqkw6ddg+nJybK2N5O8i7d+YrTMPyOi0aDCFWwWFAVKq+QTBDXJGk/Qb
CedFSXXsvwnEhYo1Oj19P7ECFNduUooW0JLJLq+fPXkAU9yuCk9bcG3rdKUzhPBiH6PbE0Voz48y
edpmMx3D4cp0SpksXB3AY+woLfteTiOWvt1C3dy15R6cRKdOw8csO4OMsUM5UE2tbKomods7GLrs
TGgt6r/yqBIQiJdr5DYQxVrDNuXaUkp/91UxwWQv8hXeaadw7h2uu2vo7aWDToYodFU26T27ymZP
rRrW/YBI6KwO4aLorSAISeGUIxXzgYDrUY0JmVldNtR6ARfnzlRhoIZ+sASWZo8mHUxgFAhp2cHZ
wDIgjPjX9kWQsc12DHG8MALzKs9Arh1FBAc9PlEOEdxqaFsCvB+JZokZwkBulK8ARaBa4/7papDX
DJvzDfMPQjeYVBKEOOMS0W74mPk9pNmQTOnBEnFySfd7xJOq99zkoambwPPpwCAr2dF5qZRYkzAc
BISO+pE/SXu5/IDSxUUfmyJA8iYasi6rgoxADaMJ7p/eM9dWtn1YOHTeBxijIrQ1W/FIDSshKJtX
L9DL+065vQ/U9xLJw6rIfDF9PXd79jnBlEtCm2Wyp5qp0msl4sbocf+X3V922D3FPO1cDWBvNrY5
Lh72jOIgMuBLgbkRf6kgxTvC2G82zkUIHfEkhKJhrG5DDVRv6g93Q9cq9tf7vLCVAh+LqWpnXyPj
XuAIxmf0v0+DBB1v+FjAhj7JjyKH7GYaXNR+bUlsYlll5agyZDDUaZPIM7cl+5P0+3/CcPmNgwmf
lJ/7wZeM5N7Ij5PNg3+3hWmgwb/S2CBATw3maPm4bTgBGlEIvBr6NZyhJ4jFXqRJjdYi7dZ1w+Oc
XrE4Rb3ZZgpoeLbj/62O3A5uxdx46ejInkvk9v3owYfNL8qdwR7coqycvSEDG/VvRGHIkjyE22Z2
yqEfe5SMZBmK5uAuAMih98zAUykj4laGm5NK4kVhLh4Nrmpv4ESqlWG8prEfGX68WQ6WxIJPescR
NAchUjoO8KvA8j5SI+co4TQ3qIHqOVBRZJcwvANPziiejXrcSonid8TMZUL3mwIDIc0y3BZor2sz
T7X+kvLynFLkDn7yEO/MLAN5JiGVo0l5VPV3jFnX2ptN0fTqpKYUJ7LlZmY44ZFJQBTOk/AJEuXC
+SCzG7xqzt1v5Xj9x5MVVK8jfiIPkMiNbwHgCDQitbc5QIWvn8Enx2vkuMV95YlYAvxgQ1QRHEPi
1Pa9ls+0Bhoue+rhGPSzyn9pP9+AqT3y7QxbR/NLux3A3WxYY3VuJ//yrD3Wm0IeOYJSPaO1nvCz
Az3FAsrROjYkaKMe7B+2LQSy4292JJYLM7ywBBYkWlYcwUg/5vQ4bDeGS5PfUDV7BZpEoAM1r24Y
oekEIEsQDJn9ZbV4h71NWGsd89Nq6As61GDER4jyzH5t3NpJ3swxWamxZ+Vf8vvUXNGWjN40Jam0
EoqRMG4bs2YJgHgzHJbwPQLSbmUyg1sKyptndAoUW0Ad1Nd7i0xK5FYENghcHxcb32VN9MBVSbu+
cvOuQgmgOC8komPYwrMx6d5n+pTZnB8bIAs+3TgjwCrfGHReyMupN7gU0k9TNQBXOwYf3Z5N+ydj
sMyTYN03z6JuL8+LaH3A5zVGgRsyVKZjEfYN0NlyHbRrAYPGxz5sVQ7gZzS9zSudXRqf1tUBOcF2
7H9exxsQaDN4rjze25IK1jd6lW6MqsNQkyOV3xhcKYc+iJCGaKG23JsuTuFBPIhOjwxT8Euvb95A
Mpv0mxgV95y2HajsKcBwDVpN55y1LNdcy2/PAPm+sUgynGF1lDA0GR3k/hFkGRxRMxW2I/FJrYWy
WcWAyptgTOPB6gd5/2iQWraZB3pklHpHsJ6uoxfd+6Ch61WsfTKioygvE/BwfB9o003sI952MPp/
nJgmKz0h2HiwPg1xSr21XsymMcFaGfF8yN6vuEP6nkklTiPmwMX8YQr8M+Rh4bAvqAltRpWG7XRy
57g/xV2D9OPFborK2FU42tl/k6LlSaAWsybRzrH025CM0hFFa/n5gtv7b7Cb069GQ0dG1f3bErOH
fcGr26wWjE0IndGVztnlX4iP+ebJb/GBLFJ7qp0TBEl/QJXekf0Ln91ZfWMIYLxAfYIlTKgWCKaY
Kc59aYwvDALLBwAAIT7jb/DBaLwanT+1Olk91lq6moHMep9osxHzObTRDWB9vTIGmyj9jK8faVWN
F918WeKKu3/Dx2y/xobjdZRjtR6FL/0GZyL9yov3TJ91nMaF6XpcEgdPtRqqoG8FFNVKajYgjxFo
01c5ItepmtB/BZILmKjxr+5vc0INyD5a77Bt0tCk1YVuq3UqLwAaCrngp8ZILvKRSuzHf/AxmGWg
nl/U3ljBtC3/5V1nZBdgB+yI9G0wc3g+cM8koVW60F88a76A71hjJJWEimvNO7YYHDqOEoEEzj3x
s8QjAKtXsuF2+ytvNuK5M5oMJQglwfDPLs/gwyoo0CGkzIiULTvKNJNRnPe4LZuFHyDjOfezBl8+
V4zJ7mVEbDfokEHT/hP3RDBicHSrCjCrx1O1XWE2BHpxM13gPgXrqOgyepDLspyiESNPT3me8O1W
7IeUuPDn+oiQ/475MjzaeGS7mrElPoQSLxt5ZpjsV678jH8bt27VOdjJIiaBZRbFDsA7Un0a1tLv
tet9kej7mJCrH3R4I3Jznyj6ORr2ACCpSXC2kSIsGlUukkW3xOUtZgJVfaxYIWD10JLmrf45Na2X
QxRTmOdYPVilWHN+t2ttB8OJySlWYqrk00eIhbvTAEVASscuEoJsQnX7EWQfa7MaRrJju/vUKroE
s+7HmzUC7zgr354aXEXtz2jKstP+kizkT2ayXwB2RnElneEBW/niQPaLNQ8rKdcwd3dQ83WpRZD2
wcVfZEdjlUsT7FLozOSsPQt6eysFVLwiaH1Sb9gQ8anP4IUI7XAsAIMMEkNnp9I7j/NblMr505k+
i3xaKsGU/Z1tfZ7q+Z6nUeeyKmHD3BNT/vzfH49gtIqaffgf+qDlWF0nBQ8zSjwnULcovG+sVF2M
50SUGC3E4m81mFQIpw8uRrEZEqUgwOX2+CIqlVcZRyelrnz4ViFMpBrZWdxptiMKmJKiGGJbf8e4
9cAAFZQ6wH5a7MhQ1Sjxoz31y4O/cFcuUHLfXmx4kGjN2JP0korJOM16cyvKtQHEdGcTpXyZ3cIb
GpN1UNSfAw6wp6hLlFYk3/l/H+jhGd43MqyHnsr1JQRhe/NGRns2moofpX+eslP9WITpV8bZBFTR
7BOZ3O2KvStR4+aLz2U7H/soX/3zidGHJUtir6YSYgbGVhv8RkZgcfnb1T+3lGaMwJSudbKeaezp
/lXdTpNXMyMzSLBQv5iF/WaqNY12qIEuYGcIdTGoYxCBeWtymx5rL3rqhndO+rv3D5+hmLlCZBCN
quWhFEcM9qXN04XyqqMVdTYXFgjq7c6/IIu0sNgHb+42rbJmFvrQAgI33abArk5tRrOhkqgKH2rv
L11qLAAhtP9008sUpbwLJSyDzx00FQpy0BIpZi3fTVMXdvCMy4yCZTTeBJb3SAOvDr5ZM0dF21hN
YLv5Cr9hQh7MIbmufbzbNfLdqemzMy7HbvrB3WApKe/3HZhIsl59Rm+En/1Ei2q0lHjdU1u+uZ5Z
c8Pv5ItCqqbPUNOGgV4t2Rdbel/+XbCsfpmoyZWKJgLeRjy4laPJIbgE2yauE0176AQMGkY15eDt
E7ydvjKKjrjHrwVnyR8lUw4g5cTCsF6QG34tGl3yIyJD087TYkPtpWcxk05/csVRHMryUwqVOGyy
Pqyegwu2lJ5ji5LkkDmslQ+FZbvdmiolbghtAOFYw8G+fBaa/CW9gIFH55tvCY6iFTwxZ5QUDD6V
Th4cSi5ferIy/Y2ikTF9rRCk1VLuD3pqydE4s+IY6KTvlS8GnaRbwUxmKiAqpIwUtMiuEhyEDZ4J
MBZxz+IWfUYmV4FO1I8mDV+75ec/bDeDXSSQPCxr9af0dIfZDwS4261rA6wq4veYYp2Oahxp/Mdf
VMd6jvNbmCq8fdSiSKo6kYz7ugE6P89gixGGIgM+MW2DuqtEC5LV93nPSJ1tUyjRBtdRV9zdoHcG
n7GV7yFUhwjqNUGW4QxooEnk8GuCp6k3YR0AfEEBBZvvGb9hsxiEjZDvb+aPwq76VLRl9QfC1emY
JFX7Mc3fCxwN/tPNmvCJhvW2T5av41BjbfyaQK7XJZswb9+cBJYtgcSe26EklAKp7CPWbLqgrj3+
vdH4XSDejkBRw5rFJ1CHfpMFjtm5spAxuwvlO5SLucF5Fgu750QZLgZelgMoVa0cTXmpFhtfVgcR
P6E6a4JE6l7alCeLKDGvg1Z/qs/VNqGNGoi0tdDEJgsaUSO/CfZ1VpLrX8d0F1FRfcb+RAEEbtWd
x7FfjpGlEhEa9cZpnMYUOyC+6smeCoqW923mVhJ6Of2SfkIrst/3kNlBBHh4sRsc2OiCzWtlQmp8
3E9ewXtjIYWMsUr/QmvHF+xhL1vkgzT/Ah8oidPrmCVqOxMXhH3cTVQsDfnJoHq5vqYsUbnN8u6e
hkAv7K17iZSrjD8a/RERj/7+bFqVarcb9KUdfNb9a2UOIHt1z4QbztUckx6g9OLWrWWU6aurPT6q
tGGuBrWP9qGonqSGa3hGYOfuVnJ0Q5Hqlz+ojuTkk1Mq6Ersv0dakPf+prRLCGRHLWLy+CUsWX/5
Gbalh9goDzQ89iLGIto+DiRwD4vOupWq7y08YL8SX80k+WrNYKvvfaKj4AuagqiAGDblt/BNjC4G
y7oMz8U+jwNwQeYMla8L6S6hGyxf5HkwWoEpz/FxKu0p9csWZ6jB9kCAt3rAVwTBpsvrapSwcSLE
rXG9x3edPiKCREX2eL1k2d02ToB46+SKAw9eES/FqjriwZWXVHnWhM+Qanna0RUmwe2601HM0/bK
uW4fMxnjT9CBwthm/PONUzMwE09LeRMnxz6umPesjonWBbYGeCjmo4MLBqFkYeRVjIHs9H8242AP
yMkz3ocH7zOADID74AAEFDaqEjJ/Xlxm932ox3QKqE5KIMaZdvPxIcPzBFWsJWddDU1YCsFG3piU
iuW2rRZv17d0OfWl1aQK7FTKUGclR4QpPsN7a7RgUKBTqPwOrRsnqE+ohbBE3OuIRMkUILt3swV4
YXvRHYNaJQFWWZV/hl/AC86Sthtfd5NVaHUQXuefoQnHD7mUav81oHEIMWgfwoZPFhxcWtt8vXDT
JohVSS8kZ0dw2dBrwdrWaWiHsLvIXg9cSwNA6jtbDifHZ/i2B054zEOzqhIDxDLdB2FtCr+6v8ef
wPcepGqXnaEN8sliMjlLZZKrXgrydlZo9JnmpO6wv/8bnWQXLjAeooPEeZHXpeoUZvFWqBj7M78M
q980VMzxwB2WQFruaa85xfLb/FmeI9YA7VmWMzWWzj9oS+uNlRCh+CVw6f6hfuAXa2flS0okRK2Y
4+g2E4cTgAKvAWeGY/OITaQu3o1/iMA2Cl/tj4nYf80NW2HHvXzWmxhefqs/CqsEY4eAqyXxplUv
DLylo35pALxgPIKsxD12s1aJF8DK6NL3pOEAhyu0jlCOIEH6wUrAyXpPfbi3MPW5fHUUPTsnxl6B
ZAr34zia+/wVPj3DfiZ7p97q8PjolmofLlzxviYGOkQDYGrdtw4/6y3qflzBf3E+ju5HnBaxlEp/
hrEqTv0f8onq+yjFgcOFpwTkvjm8hg45tl46lMwZxlCk6MqDb3nF0ak7khtEg6RwTW/Buf0ruh4N
h8s9xIzIxz/R3DWt6d3hY0TYDf3EeRZD6gPQO01I0SMA50ipEfm+cXHNBL0OVLOEGi2Psi8rIC4P
loF7hb9IiWGZFK8jhYoo36p/XUza3IxAhAvj33MxwvQU0BBAZRfyMpmjxkgX+DcUJDW8lxWcocwj
Q432VGCtxo6b/simFbklJIpLpSnA90aZeMj4Z1yvoaHOvKAyxOOeo7rMS8y7DrRnudj8qXh0H21T
Ez1IC1tT+Kf5yC6PaKcv3CmRf1etiIe8hGMGx68rgzaVUTapfby2QwcG2XtoSitpXJl3vWCMRAdG
LznWRZGtw7NmWRu8hCNA0hg4Ggx8xeel3g3fyli0YRGw1i1t5MsjUfpNvB+3Zrl42tY5Nn0Q7pHf
9FhW1Haiw2n23nfK8hYy9lilJGh+MB43u/UwKj463wePPGH+2vT1jydFdxLtG8HEWeQnlZ+lPxVX
h9w2oI1rhMrbC2+noThXlxw/dvxvGsVruvpInA8tD3BU6oKuybUAVUJCf68ViPRE2rboWZGhvll8
9S0wsuQK76X5C+foEJviL6kkWRbqlKxQRmfuqJSMVJrHvUhjZHoTadr9+Foox2FaGZ55Kv/bhajP
whLEGJfIrDubS+JevjpCI0TqWoQnoRagSf7hNrCkJoBwLFta5toigZPbv2FUDK0MgFLsG60ZpaDD
u7DshQKQ+3HpBwRmVswzfrP0rCOwvePh1U5kpDtp2F++aZ+9T1oD6zL71VDE7BKc5gZBlgEd4gmB
zuge/qSDydytl9+S3TLJ98WDgzMCUDJIEtzBteAF67IfxMNgoRnBQafTqbK+KQV3EA0XqolFu/PQ
e0d5xYZmrYXEagYR2J49mHLqtb96oAcf4RRdomNE3rERXRmagYMsNVKpbd4egj96m3jTvuH9t8gG
/U0e+f6g0cMi2LSRFvOKH4btcrU3gh6ASUqWuawFvfYxGsLbDMTRkvVr3Zv/TqEq7jYq73QRsPDd
IGIWOgLwjfGsQGlGmy6XTUD/QmK/gvBZ04MaQEBOBKs0K0jOT43UHB5Ql8dEC/odNMgm4AJTmck0
7LrEDKXaSKusYUWtaSWYNT2AjIBAnzhmp9A490dGa1IMDjpLhlcfAGcV4VUx1tZdKy6+FEeBpa6Z
prh8UaIy8rQeo30DQUGFL3ecvjqjEfyimSWq8i7vTFZSPXIat/k3I/BJuKig0iWIhdCSSwTulNAx
+klUBD759MvaDdXqnYRDnRUwcrv6iboKHRmjgtXdhDTvgDnsNh9nNokL90d0+b+b9fzweZtV8XNR
8Zoj6QBcqb0KUa+7nErVPp+e7WGYE2VHL3WL/IDiiaLs1vzRWcJwDrfSeDWqSZFrTjLZLEy/FBGl
s22jH17YFs8lkTwQw6Paf+yoy/H3Q/zWCeT1cOIc8pasbVU7tQUUXu5sKQkyd6lhwf1yt3zI7Xoa
AUPOr38AgKb13iSI4ykcjysT24b3TGQgmzTukc5GwWzMXRSvcbTgMmoBKgUKARJEoyat3YJo9dBE
HYEt6zL2dEydmp18yXWRdhOCTOUl6/4Tf1R+I/ZQPnyNqUjZtv0QYG0fqVKAD/45LMOZTZ+dhddO
45hMtIS6gDwvfzBOzKl5B408zwkyknslN96yuQNBNMThD9NnbcYQr3ghEZZ90YrTVmr2pexmcEka
wb3Ulmf5rgjITiiH+uQt4V8rtkkCZSKm0skTwoZq5Jsz/8CKzutIEbHX5/VEVmQSyF+vWO0bIj3a
FiYskzHi5sG1vQbaQLVnKyyJbYYkpPtCTpvJpMMHQfXF0ah9w98dNtQPWEx6UoMUeJ6GAg23k7uv
bwxZW8G0o43PApmlDK9Vf1bNisjzENkBtKQckEGIJR5m+tqW77DrRLLdLyi/XmFexSAaONQ5wUya
36rxSEsNHxZfMvmlCNm4aN6rMJKititmH2eXKwao0zk0VD2Qq15SH2NejJr+lIRPLyHRgqxNdrIk
EikX7dHYp0yIkgz43CHJtjBH2QN5bOJbqLoq/CE7RCrf02h37jPvBHxcelFmugbtim0TQkQoGupm
oUZpLtgHT73Fx9srPcUksXipCyI083y6J19ZMRz9xwZh+Ud463kPA3OxMiSovCGmQ6/av4U6rJ3q
GZbqjluVOE6vbzUu4ctsJ93hRTibfuNr065zyEPaFPq7zAWb6TGRs8iYaZRJqgzvHpImh9d8AYJX
5lVM5LQveLJLy0A8vL98caaX7ZmUC6Y62JpWvRIRb8BUnZrAEaaiI+DZ7TLksU4gnIy245Rkh+V2
hzVrljQ/uCm/2hTS9SbKX6hZ9xwqQfd1hcleJQ0aXQQpY1KOPc+7LecgK9Gy9vMsPmDsJONakJ9U
Q8pNCwYFkXduoABfQ9f25WwxD2gT0mEwq+HX4EDv0WqExrJ1kAeNw/e8f1D1RaqwatOnWiPSkMGK
9pGl7U30HkkfmVGw8hqc6VZLUaFlGX62sdku3tgXtttOtT+Q/n7G0yZzzq50GWontksZQ/QST1ME
JaeRzLnwHq3DCNrUAbkGMZ1jeIzIyjVBLTIHKRhYwI6ELJCuzgOf1eLXKYC9sEUUhbe/uJEjug0d
eCTKOZVWN4Aobayz9IMYCmsoO76tFjzNdWyvtjRHokxXpAoWQG2SQTbq5FKzd+xXxqFnabdUcNzp
cMRIxne288MsssnbJmfMA7QyhbJZrwYlRWiP3Y4Ce3DMvm0vGL+51Axy1OINTVBD+W6nQ4blUbfR
rTzZ1A2sEPPEXva+iZGIFYuyP/QSV12uC2yvhcWpRHZTi6jmMBnbCmm08YWlpZ7/LH5+qI0yvvTb
nUI8P6acu+ExG3Hx0WLnqDRFrq+qsZikb3Tn9U7m3wOTcFawzOjkXCCRgRcDtcGPJldOPWd8h5nQ
wBgYajfagDO3oahcfzNnu4PGAXhm12k4lwR5lmsxMd88C7CO3t12enVDHJpks4vywJVeUZ6iakB+
+KR2x0KIozdmkKMg1FnC23n67P6q+h6gQmsgUTiAoXX0lnvl5Zn24ugXIrYhi43M0Qc+MsXw5gM6
F7vsBeqW3D8PH45bNTmiXLeaDb1+aRFWH9Uek8+lXm2Y6BrGBBWsA7Osfgu/VjolWvR9U2lE8DEd
iXlC1Bf+E+VjcX+95MRG6V/XQGEGr1yd3HCHAnE5VML+oPRmkwpOM4M9a+mH24KB4GtdX27yAR2u
zkjs7glbw3hrispOccAV/l87unZZWTIFQMSwlj6mb9cRtWm7a4tptJgWYilfmDD2PEr77/9Hglca
wkFp5NNMp6eawrkVlyZJvy1PGzIwyHp0ChtOK0aqQ/8B21pAexRm3iTNlPKFbW4pfyI9IBgfsCZL
MDE9HmrEH84fESmeDj/WWFIaUtLcINrtltPZBgcXvJgKqgSYF8WCIoUJmuIwOW+eP/eOzhjx+ghi
NsbPDrzZTCZ6hHoY1jiLzLSsECJlEFx9orcfu0w7Oqd7ZPe88z8nXYfMWAYz++J0WHdoczjUJ//l
JGPLSSPsaG2oAy89BrU7FT8sF2rfp9D1zwbSSbOdDndp6SwmgXJaK29Vrh5q+B3GBsmOU+0wvQNz
s/JBnzMhLucdvupY4FEOcfDc6u6Df9c5Jji+dTQ4Tnn8N0zQ+eSKngeOs0vU36VKaqZ5LM8PqcHv
9qFn6QMFGK9xsOeg3ofxEyU5K2fbnMTzNZTdoixyFvaNTHZEeCMbM5AkKwzuGfnN8VYzoc9ykXrl
+hNNPP10hVBVCS2GjjJiKdc2H6LSPGrJhzQrmXKS4O9oqh/EUflzIbF4OwHyLA43CsZ7wFtctvxS
kzL//BLrjQIBc0trV6m0OihvukJ0X09SgecuDyDuiLjAzDeEmgr4mJCBSM135HAB735mMSO1O9IL
eQABvJFylU03bsNXMTJfFpNkaVfpokTgfdxXR82k9lh4k2F19JL67e1EptYe1mTXA+Uc2bb9aHvz
fZ4g7sIWLuyfQwN0fQP1ZgmfbSYycUCmTHT4J3Rm6TDpbSo4afD1x45rYL2gkqF5gmRS0vtXCEte
5RkgVxAsbjhv1mHV6NdQyoojaektzOktaEWSw29iGf/xiT7JUykGF/K/03KxLR504lP83tncIX6O
CuMoVzbNNS24HBPz+Rknp9rttIO1w5Dw7K/YDA6ArJA7/Q+Tup9kzwu3AHdUEFmHd1IzBvZe8Hgr
N+vM/qvZooyVdwkUfgiLvcezi7MDIndm3snqNPjP67gfPr2CcVEdDWzn6Y4IB8Ea0XS5PBLCZ9ac
HuLQhKe2UVdzJSNiBi8f6UH5tlXTUxly9Cn2Xx6YuRkeT/C08diDCndrC4CiWfyqRNPo7/ZBsIJO
U2Ps1mt8WvPQcyZymez34bc8fv9M+DLZh+5NV72jHYnMLfEbbQzj5GGp5M1YAkERq51SJVpL34m+
DozDgdkphv7KdihEU56SJ1n+ehqqLYpjtXu45o4A9F7fFgRPIycaiWLYcsCMBlWvmjP7v6JEm2CO
8/AGOgIqFnhNFmaUpPIu8l5tdjYozc2MWypoKPEZYiL38lpOCM6kxPMnCdd3Brd26zo3Ygg81z5h
b8PrELCWlNR3nNNo5rTWQQoxmBh884UblMAZPqxuWJ9V191Ke5Vpy0WwmwnxnwcSwss+4KCbogUr
wFdn3D6aJznLDPSO6pHiI3rk2j3UrTj4v+a3uGZKpPcRB+nuteUHsBWBIh6F7jIwesq/e2LMtQif
gv2aRaaXkZOCo2A5oaeFJq4x04EXxSv22qJ4SB9TZzWLE0ytcirdDlslX8Yq9YTs7X53mmdrpDNz
SohSJcnvM2/tBJGVpj1tGQSjcGpN/OPmgpAEgYDX/KThHOWJ/Niv7945xprB9XNw3JloBaNE591Q
fnXsYWJOU5iSfn+B4DsDqywOvgVSRNKCy0rHl0bjMZ1BEWXKUqAy34FSKJ1S8GbSc5cycZUNyig8
NAQy8s8N8/9r+S5wq/yYyPkdjUfBhQX7PHMAVetAJz/6OoLiUMtHfId5pLXOVuALIbngYVsVQzun
RCuJ3yUjherlCLYKpCvi5lSRigi+57+JzmOONqaTNcpHqTnkCdMZ2iUZTNVr6WbiENgHhSqtZkUZ
VnCbtk+8LGYUT8rmuc/PHdrnD9iLCl3b/HzhBePrpIA+fpnoggdJQz1ij4dMnalPfAk8Uw9qAz2V
m4CNhqfzOMjFQXUompFxo3EzQLU3qtq8faXjxidkYjMljIM+YN+Q40AN+mmpmhREHjYgy7qH7Mp5
pe7NUECwjptkDqT/tTtUAIIJaUJdnecK1xMV7BDX1FTHyjKNfoV7GBfR8bg9RiSQUwouZbWzNa/P
dQW89dmLIrelSaucN+zU3ofTcA8w8OekXeBhbLScOAlvTptjt4K3GpMAwzxNZ8yK9KTFmxbutULM
AN2a//n8Bk55o+j7xElc8gOZxM/rpKbE+zDi4uUZ2XRjGwMNTYShletgpQqjamGnniPXS5gCwWL4
SH1SSNB9EWf2uodwp1PvqMwXsMScKHKGqBBi+paz7iS8nzGqHn0nfjYkH5x4cqm8cP4adZYWM9bb
o5OqmT1cvMlYPKttTMJnDfp2fZgLHLgI7Ysf859qC22jaOrpJdPhmwN2Ryx0v5bqKEv7NIf7VxJt
qUfa7miDtq3Gk/3h32NemlbwcwR3ECwKMhrsrz9WVZEpbvpmv3HpbXsjvNt9Rwc14omFRZS3VT0p
mqC/rmY0tOq1dRe9ytnogZS3vOXhLyv5i9j3R0KOBOPf9ag13+7/pdsH1tBKyeS+tR9R2QRI1o4r
RJ3F7/0B/u/EjJaSCdM51BpLrYNhNhuHG8mlRSyuI0g/jUd/Az9l+qfr5+CNKGjMmjapXiA7STtR
T8G/HtF5f4LMbSPKejM5ZD0y3ms3qtpoqxFls6pZlTzLQ6/vaW/KlRRU9aqTlrimqtsH1kBiEia9
Uh0LzTm+5O1YdtqGK2QfeVtcMCQKoVO4tqFIQWntmKA1SSixNeip/S3YW6sVmYrvzgkp9LPGJ9Zy
xsdO2h/bKUpOVRAb801j9gNXsXOS9bFNjLgP4cMDypSfRHkvmk3+0ze7oRRYZUF9jY8wSPdnAsRY
1UCcjvPN/jcbmeaZBtLhdps9vZEgkoIvpGfgwn5fwLeXTnSCoi4PX/Myq9bYTyW+z7nmEl44QWKy
0O3+sDeUxGKF9u7ynFObWRnz9dlqeBTivG/D7wY/FWIEyGH2WpCDeOpdGLLoX2W+dU35WL6Lsmh7
qmtNR8hMKzssGkaH3YrBLBvZZIIadHkR9FL/RpFp23w/y9yl9io58SxV+NLh3LnzlX9usHPh1zX0
iQhevcg9Fx11BrSBUHp/TmUn2rYJY1Utu0F4udpuHG+XmAWoVP/3XPqutG2rXknfdpLzAVpFlnts
e6PJ91A09FzfUpasFayIuh2RyPOkeJWbFmJwWzmlnUh98IGMauYGcTXm0ZOkRlilsv+ZQb3iCpWj
pWv+K+Pv8BV1WUYaha+0UVRg50+DxXNJGc13259FsTsCQ9G3LMLfDcJkFXIDdMA2n1O7NB9uisWv
lmvPwWvL50cq+D6knL9nHSaQluIFe/qUP7pfX8WxD4VIxZOfTyKqUxFQkIJNxF7eU7e+DF0yXS51
BdwAWZyITTHi4l4xgwmLVfZjZ98vPLH61RzgMfThbKAcWQWSiKMuDHAk1YQqZsvzlBRmcOWkEKsQ
PiIlMYJmXk9xzVXfsYWf/Wq5dDpJo7XgEU8mFRCOpqHiRgpk1mzONDeG3wAe3rUxbMsZuRUL4V29
LGxtFwpFxxLcu8TjMHItleo6nkuHnq1rW9NuQShk9Ya4S/mPsEx5WqGL8khnwgsE7H9ibvSJzZVh
3V66YyCZoikD061oLJk4O8dL9qp1+zRw9uBRTwQknyTQuHlBoDTKbV3my6TPypQo1G6IHhmq8571
CU2R/M9dqlw/aMmHxp1usa+C5wBtVS+M6MVFfVXDnPZQeIzOQQM7Uo0WlyL7J4eJu+03RNt/HGdL
AemPn7ZOEjBPmzZU+22D0sNEHdb6k8LPXEohJquZsmJMv/lX2w3U7xnmtj1as/IQfU7WNWuFVwK+
58csBmwuNKrcRcgmUBZxm1KC6FDwqzrQYuiSBKewG79KBbNzqrCMSvRYS1MtGzZCR5Yv/52CO3hZ
JvS6exO8pawmROLxeWXrp/AwpmS/DiCroQRkMHOhTH9zHX/MrNaziFB6NeKNVfZtxGGNFvhQlAU4
ND+1lpotm8O/5IQYn+iH3uzkMrGOib1tKQ4b/p5K/CDini9uz4YvNJ2Ymqet43KQ410W3Rpz8HH9
+/uNcDhsEZKVw77D06IdvfUXaeC8e37X+8/q4bdGoeGuct36pF6orisnVnv9Y9X0GlWfY9aL5TUy
2ZolLfc8Uewi9ksBNpVC6JXnqpiMZnPrWrYVN619S3NPccO6TUhPKIpn3nomLnXq3qe+FjK7CEAz
bEv7EoY44zMDA8V3/MK0q7QhZlUepb92WRJkImLL3GMft5cqn9nFWeB13WAEKqqLPp2wVb3b8PcF
5kdzkEEWmQ4xnJGRzCMk1dhNTqm5YCHCwKuzUgU+t6TPQeUlYhtIio0jR4aKsVm7S244xxgTBEiF
VhN558TMDzish3Sb1U6rEe14cbdOIuGEIjZHr/Ry88mYEQ7+RitjWqMDn9KmkxT+KhP2BywpkG5c
Hfm26ewnK8v3edUfOXOKdg4/ehskiiZmYnW9kS6+Cdu3wxEXCo7SSEl9p7JO8l+2Q9hUUQb1fkcX
F590O9nyO6GIkwEiiP3i9cNyzn1wjpFbwM3wNBX2CITR6AB3vzaEfEjzYi35vgBRB6HlqvNWidAj
Mhe/mJyFQShdI+N4xTnpF4Mba+cnQVsmzYIizl5y3y6OMXV32xXv7TvW1dY455vMjEh3hZeifN9L
TBwSe2f3qqFXhautLDj3MbF4UTF5NxSOvvl8ZZNiMazbARqYuZxy7sZmNBmk+eeeDAnu9Pznv2pq
Bg8gNzs2stkkMcJdmhBwDxjWsH5laZ2MdxLy4M6PaiWyUHGVTNEZ3ffxGKBYEg/Zxa6ZZFOfeSNm
PA1T68TTBK+jQY62Vzb5HqK8M6uiG22xc4r1QX8uHT9VhbzUBUlEjIIPbgHfhzI28mAH9ABOkrMz
UnYfCCOWDTfZciy8CdOHSxUa7ea4QL4ZxUH9jXYfzYBY65HqRdQpFSm9OmQGTOoouWJ7vwWTDC6q
P2gw1fiyzQEBJg85YXJlujHXtRf5XOevS72VYAaC5spLiIZHREv1EmMuZ3P+agZXH33/fdi0ZXuS
QTlRWIMcN2hycRUcKtga1CN6PEC1aP5eoAQLhUDVz1LZjCEAnrGMbK40AR/kPwqytYWZUI7G+gyK
WSmMhqxt63667XL8nGMhuQWUUZbRFqq/lQOFjOGCK2rCv5nRxy+wxlHi12atlX5iR31VrvYrenGW
/o5ZvHD2YOJ5KkdY9z6EG5KBFiWocXcXiZplU0U99R2BdAe2P8mplKAiAsEAh1bgNkCWIb0QSz8m
sY4a+MO9xgLSzTlRgfukY55KCUMAUSy27buzUEqob5R/JVtIAZp8kpASy9bNtnoeuMbUkNxE+1hI
+BEhfTvbNdgwIPHZISuozpToRfC8cUNTN8SONJOs+3sup5C0C0GOo8dPlTsc6Ze6b40Ebj1OYX8u
Gx09QfSHuQBDzv+VWHk3nL8R6u0exXh7YZgcwbn44xxrKu76z3hiubU+qIuWo3StHD3NXwyL8ClC
b7KCSGgS7M69cho+bbf/pVToD9KEb6790ztd26OkL2LHSUpgs5hlrkLivWDafPkfb7HxfuflwyP8
BTyghSRaBDO1RBk4reuFB9kO/KN8YZEd7XVlfilBZoBmpzNJ6sqbXIG6QQr8XBVHbvQCM7PbKWdt
k8nK3xSi2YmXjVlhzAFh8ACJTbmAuHn0+va5dvFIvvthiI7mQqzE1FfXjCKlyDNcCb0H8RS4tEbU
bWcXZk7khra/OVkGJHghmUaK3rTh0VksI6+rvNVTnSBZ9m/JBPrhm+xuQ+pKBCBRbWo4XoQIL488
mMvGyM7WKb6CI8+cWZCr6zK38CpDdDR/gM7qoYBSFQcW7O4lwMAk9RVmk2rwmK/4Q0CiagD8dCVW
aqCjID5L7ih1enLBZ4T04DK6hkfsTly0Ug57d7RFCyMdcJ996GrnzQkQFVRiY+ANK72Y3mPpqVpf
bhFyB+fq92JGSkT3ToU3iAd1Udt0PyDPJuI960hkWX+z15N0W2ZvDtueDMgncjCccLVtBQNlEKuh
QDzvBDR9kEKrrPBn9svsW8MTs6n9pK5N0HjD0+gxpvR8QQIb0WxNnhWrprthiFsgCDS/3+wVBsSr
iEP3O2sTscO07/WFP6fjFHbrn0JQqH3BeEpCmVYSK2n4k9i+oX+U+2ij2sDjcmTRzspmt+JJoYMk
z1UlsgfEhidfeY8RhIyJR/iTdx639Xc67Z2CVX6N67m9fKfXk5en43Wlj93HFKxgAB5RUhdq6VHE
RoPGJgDO0uvLcTLPfIJvaDywVzU2V6519XjUAJHAJ1qF9a1JAJYoGL/hcCmdhp0lO+mj/voPuDRe
5tkqvxPIyd86hy9T0z6rSWDuf0v5OKrax/JdVYoSPEC1TRxNM8cBe0wNDo7/ndjbOwuEPoCtuAX1
5/e8dDf3zcyacn65SSxb3iUD5w7umPWeTNe7JlBejJxT73ydmljhiaOvE7GKvcoSStdDNxKMocHq
BEouLrq6dT+MflingJvNHraimddI/0EdO+boB/Uc/feYxHmnoEhz0LwsUmbShOgfdMhT+XmhKLvb
12A689bB7ECnfjQAAU3qRQn5HJUE5gy+tHxDf8NXgqUeun9C6YQSNAGKdzPOqhcDe48Ehr8Hb4ah
V6Q2sOTkvqCNsPA3pknbZQJf1F+Dvt9ONl773Mmn4hpjPb/NZcl03JwnallIY5QbKM4iSvKKCAkm
l4/At9Lxx86NLGB6rDlTXkk50DHuzALsisxYC0HnY8h3yR+Hs4KILMfH2p83cEHG4Z9xVs2tYKpz
FG3hPXxjo1RqyS/ENkfPSCCwDVVCOz28JbU+CFQgg/5ZjZErORlidCfVDPrpz78HISUJmFbvwF6S
eRHvHmsTBY7BFF0dSUol9ghbc7nxm3dhBmpxLD2b4RD4cpP8fgaHiRjc5b/HeJnxuTGayJY2HX+k
RHtMqRUDYQTI/iRc8J2lsAl8cX7vVX9RVgRu0EmkqYAvXh3NUhMTUIg43OJ8GbhdfWM82rTYapOB
+VhoL55KunAHnyKQtIbk0UfUGAPgl7mKD73DY3cEN2+Wye1RyULg+dn9l2mQ544Dai6Bi/1BVLhP
AL4P9OKgbXQCXmiFPgPmDcF5P2+OU61IIBQBwuNrsdpTl2kmSsWalA4EVoBMBKOqJR0uMCmxyBQW
QYaR3Dh8N0Jok9Q0Z6pJjCrtEIJZ7KUlBaqK9amxZn0WjedbGqxzhjfRHEL13lUrKSTBv9ajrMVM
zWt+jhAgHeHmGL43UfT6XDVI68u89O6y2graHvsttv3hlWPdG3IwVrKdJW1lI3QojJV3bmORpd0l
2kXF4jyutiZn9o/hWc2YB11xgGf96RaUQzhHlbI929ddlRcw3p+1ZEgzdc6ttOq/WukY2Svxal4c
sj724f+sBFPGPBlojGY/9/D3VvJxbpxwaayvdZGe1stGVlx1bProRB3z3nI4t06JKFpBM3rY+hzl
CG3kPiZCWWkgoOPH5jOGUt/oEmZe0J7Pt4Mx2TeltFiIgxbzV/LGr/vTjnghA3WqWlNIq0mXfq4k
sW+QndIU+t3bJWoFtar8Gu6W/bvd2Aulk581LeeQ32F0y7Fno2WCSzLeQ8zOs6BzaZqA8QrSbT+L
3Kb+mgtY2jQgEATgeHgfuUC8aFLjVPP+XjW3JyQYV1l6smQ3ElZBpV4xjalHK1j9JAFUIH4nJapQ
03qhLG70OGVnlbrNC3o8MqU2QkxvrNaRPLNZkIMzI03NckUNXwcdLclJSx0ajN2OwBnPFjVJW2CQ
hgmpooKDaX6LQUzhRasvtOgl10wiKdTQWDA8pV384cU+6Wx0s3zeC6rSeB9W6r8WGY/aA8sp+31L
hEz7Rl1jXAoj98uk3nJNeoRh1wciTEXEIrRnhd0PqSmzj5OrmmqppvMMOgxv2No8wAwugpKuZXy5
SSOEhkvfbxOLlqpxLUTuPZHRYZQVKPeyo4TQnMft8lsNZ56J5rHPl72WgHNvcuHGpzk45uam76QT
ZsvH8sf9osPfoY3ZK8G4kKZlR3IKYmfl/KCH1cxQ0qlVstctXCEW+1Tz+cJJGBAweysWlYunqRRI
XQ7WKz6hdUa/1PffodKkC+hg/Na+VIuHto94y9y89WnJ7NePl7Cv9J6cF1eSQZRb4rXMRqts9wxr
WRfngHM0JGV3CRNC7klmrqNxeh/2f2x8nKvUU7eUnz068p2tlYSkLoRcUwyanaVPn1JzvHRRJd/B
6MEbhd7eDYK64Z2cA9qzWAhv/U01XLlSR5iFREhMqt502TzljAQ7MtispCNkDk2vYO/psWm4XutA
/URMDkjlEs1b05il3oTTTFSRopFHXYti40aFPp2GESxHCSGhYv34jKxCj1EBfLa+poph1i1okuZc
MWWyMHMrX1i00GHukyxD4IDEuBRDM+XKBOm8xmjXmk4u/rLxwLdxwXzhOpvSaWv0FJIpfYP3yTxc
Z9EKgTeakfV0VZBYVDUNRE4x5vblERpdwmVpBr/7hk8bXEYg5KZfBO4SirR9OOIDjlvdfgZvByzV
QPbQDJnYHpJphSfBQS/taqKRqNtWbEEDFwXsq1nkWmznmO7I44Hh/+21E0juPqe95KdvGt8uBbWL
t5H6Qyg9Sf3lUC1X7UUrkiAMkFEa/nDRMd6t4QwSfbbUFhtSXdtrNgZG8UZ4+SK7a8cwinxM8UuU
sUJGoDbipiZsh/dE9KAQF4m0tEtos1k35UwKd5XVW1ziloRYDk+g7bmA4rpqfG8N+o+kMChKbUV8
abnplwnW5tSeC0kp8uk88TrWM2IPjqqj6Fivj15WHGJUfcv9Ja+DxSfGQHYmrHl9rvIIHU4qM/0p
n5DHV326nnWjPJQuW1SP7/d1KCOW3hKbploZi52GF45hGK/WHC/9vdQxPzRRaB36S6dKAIWBQ459
83Mdm1/GOtC77ej2xfH8UEhnej87gJwleuPUU/N5O+IIV6X9taKpvlzJmAvIyH+PhKCnBPY6kD0J
lXH5NfTXJMcm0gRDnIaVk0fLpxBIo+FGidUFYpkSnLzyDMVQb2JnKSAs6D6CYOsV6PnrsUJUS7kf
BgHyrgxPvkFCbfQOGVv5aJfaotjwnvhHodD8lDi+8c8OB+pNJgAx2lb/2r2JndilZ9lKIyVVaZXt
kuUBJJfZkYi1GcfUwz8DTjHTlGoef1l0RzhgyxwjHhDRcOW6KjgZ5EugjMQipVxR1zEJaGoE+93+
210KeJR4p7WguWj76/UoEj+VpwC1FU3uo7aEOYg/LvNwhFCJ9AyC0vVUg57vP4w6OIPNcpXGOim6
noaoeFE+UbKixIVTgPPH05dw/3zAAdbTj9ZMvNcEcMKOPjvHmhvLsk2Lf3iCbO8ILsdv0gI4uOeK
07E/2bH3B3I9yZjc8X7nHcbE8ogI0mgX6AJqpAcW4C77WjV3uL9AKOjxemoEli1scA8h1tPDnawc
Ja46eTOm0XFOTbDCrRAFrADRRKnXDNN5SkNcZ58UYUwbujrNpHim81y2m2DCtsLFS0jMtrHGFjwm
OG05m/S7do8J/EkGZ79T3nR+pBuHMm06sgQRZJkd6r8Hj4KB8aEUaRwTteXmmm/w16HA88lb8rPG
admye0VzTIqEUPCPtwBaZazGkghgocF3Doqrp0YI3gC2m9o5fKA9zyRgfSgbJcIND8TeT5v6wr3y
gDC1J7FmakiyBAOYo3iL6DiR6hergxRHB+aetcKCpDbHT8OfI6Zb4V9harLrhDY/GPRtvwt9Cn/5
N3y1pnw3wHloPdKH/bB4OozLhAlyy+HFh2ZSPwGq7EfzjZpctVTZP9nddHo0jjrMB+512Kdgx7gn
4qyqnAYzMCq0ht1XLdkPfugIXYIM76KmlF29PGXCY8Zblv5ZVJwt3NW6nBpUjRBjpmB/44QVfBsM
O6v7PkTrVgFgyngYJUTIk1bRM3ikwmHt0qzukFse2NSW2DbuavqETS3/NOMw8gSa/SmPhS4ix6Rp
LKUrNNZ+n14PT0GBMWn03JfItOHRk2nx+z1xA3OyeeP+YcAJhzAyAPwnyL/E9tvCada7SBrXi4UU
m4mb1m6hpHgCjp9OzccVi6VLksIvyUfWmf/Af2QPue26OKbKiuAz3gAt2nhgDYQ/CHMkK7IDS/lJ
gULQ/BlTD2dgyEWwdDL217MSFkgD3L/YbHnYyqiFJV/LrxrPqeTN0ooiDbUtM77Aql+Xzc2AhK40
67Z+rIFttKjaCqSmzf7drYFCmuK+58Z6jSa2LZy3/X8rJFpEC4G/y9PnZ1pcaOMfPO8RfubwMK9w
HNg8XDUR3FPaNm1I8V9Fv/bZLRQNIwf1Ta43tpNzSP55XexxJ/DhCZX14pnc1k3ZIXH7P1UdspiD
5N3rdfALi/dJ4Zagc4epzYAzIHvbIjdYbBsXP04/idoKWeAZXLGvQNIArspZlTAW8kjK3QeEY8DB
RH193zyaAljWnBHGicmRn/x2UH17Liip7FWzWfth6CSleMlqgnC3q2UrT12R9rMnu7V/p0S41uSi
E9MMcxYJ2RxUyVS9/ZKIr5o1WZ9z3Zj1CZ8KbTsxtoOU56vb5I55hVKpH+0GeHTQD3Mzr6XGiff2
YcZD9ywH5O97a0Uw1ngiz9NToJMDjiAzR3n87mT9bqe2QqeHgPUQKvsWXc/IOQUi0D0MPjBerX6p
ohjWextoSFz4Ul59xz1nkdVAJnmpJO2rGJ7ikVR07S9eLMLvdQF+D0lD9E9JpApt+tuGN+FdOsV1
elK6ozQnVFOjnKN7VOBUqiME2sQuI/gC35r8ucXymtXy6LZzkdfc/slqphZ8F8NEqVcLlRfzJ+7U
3D0r4wlQrzOHuuRPmZVVLPpbMkSfr0Oz0BMti0uejrZLk6zwXoY6+vUjAo1zKWTTJF57j/JXO4Tn
ThiUGC+AgJCcG6EfmYDVaiu3A2CuDXlA7t8gUpsNcwlXHUAkZDl/9Zv1x1chKsJQQBhE6nM6Vcr7
UpNHA/oFwdG9wiHrggwj8qVJqSCELGExYbPfsJci65+hb/AQbEKiTwkAM2sYqeltcr958onxcv1I
244UqI6swv5HWOb3I+Ykkl2mVaWkF/DeK2u/8/S4Rx5fKaic3cTcNgD38IQemX9dv5qpchhBOi8B
cvz+dImYPO27QykLz7EF4jhImBDXik6fWIruSfNOWLgSB9pcZgaWsG7Z/0a6mhmXkzAFdVs2FMdt
XrDGAPkPOOrgBos0pLc02XSZp2CaWWIeXGvItzOwhWireCetxLQzhCLXrJIWpPgH/loDIe/TbGJG
ShDfOyLP+Jsapr0FrPqgImfbtcKuvkKgnBC2XnUMcNJaysxhouTpvg835aTdOkvgRB3ln9lfMd5o
8n9uBOuUJtCrkFxriZTBcai9gZvuJo7gOqGzCfNSzgINdp23yGZcdjJP9AAsH8G6BL0WXQoo3gvX
M7dJN7+6yaEcc9rA9pMDpYreP0ohwT1SmynSW1chm++CxtosLVsIhJXigbWy/2IhJsFZfG5bPqx6
dmmGSc5GGAsao7JM6Thm+xWR4BUuMtn3uzk7GrO1DVfAeTjczrNfa8JpeZoXDCk2WGSUz0Y79RVH
IqSyGAG4w6+RaXKtDJ8L08PWSyzYpNvQbAO5GN4C7DqeF1s8Vn9SFq+C93577HxQxT/VXWfYQHKI
cvNMZ/2JqhHIakn9iOYhpKxyuBj7XJfZa5y9fjGFr0jxtWWH5hE/Xsn98t28QS7ewc80vK2XQU8x
ZAUwZRKdWbRlMOxnJRA7Zx+xYKZJkIXqsdtPHtB42xO48ipge+6BBA8NdjLYwYoqMGifzuVGT/JS
gHGU2qILK19bwOAhWNDMl/zDlYJcl1ZqsddBVISJzOYRMOnlWqn1DXCBvOBQkcKddd6fumIXDhBi
RivYv1CJZx2w3Rjdp7y0UwPl6M1DVPo5vBNu/u7GlzD05mOfg3VdZ104Q6so3IP5rBrVFfRFmIKU
zmrJrpn6BFfvzV5+5tC7YRqI+VHlTn5qwuaqWH+nTvvM6T9EhAkypDyMjHdqK2Zbvdj3pRe3qb1e
6GR2NZVr/8qNXluAiiO62HyhxPqiluHIS1fsoJtk/9sJX5RyhdLc/wZpPQzYzOZ/eSpdGvQLdCVX
twSQ5HqFifeYaUoPzx8dO7uvHQjYtmFSYmvxwkCQs35lN4P/1BA93irkgrTAhNJItjqmk2qe2eLK
Q4rGsNHsMEEKxCntnssWQ5Wwdsz1DwhE5zPpMg9BrYDYpJA1migTHCiSx1EHSQzux6cZkX8cJQGK
VTspRwrpio5R0Ck9mGhUepsvxV1ju34BJMWz2spFCxF9QUdKec0u1EINvddhx6aWWj4+7CW2UoqA
F35LhIqFUy5dxQY7BdnfPBX9dAGwqh54VW3/Cjf2cfeoe1ZYiBANq0gfb4mTKAyQv8dA0aRfyzwT
dqcJ3Y6o4Pd53YzckxKJ3S9SydOZ3nrG50aPJm/vCt5fA0OC+wxCb33+A30ykKu/0Gajkv+JPHMe
nZNIeOE03Y6mpHjT/ZMIGRSy+lJYAS7OFfdA3b3mb3KdTitKcGU10/1UBtuzN6CVtXdE4wD7LhVI
XuTBg8GGbJ2zuJQUYQw00RvJgEOvviMyP0ytCqTAP18a5KKQt7DJcPlVbnpkz/dfa6CWDvX1HDY/
VStqJ6oAQ+Piy2JDQtGrhzAyP1m28t0P4wH1EZRepzQRsBvWvJHWXHAgJITW0g5ecLcDJGU5UESd
yXEoVp/PuhLug6d91x8gqFzVfzq9C7jZ14o5yschDvEmVFcB8B1dq8NRACN1SVpjEmAqlcFskqBY
CvIxPFal7dck6Jfr3Lt8/td+M/FVoIeGckC+3AdKYerIBU0upxP0yxGfEie8kVrLcgHJn/zjeIk6
GWcvTJsUUW1Y4Vb/5fvWO0M1UbxbFRoYgU/28Iu1QRQC5KvAjGOjGbii3JB9JbvICqV+HpMxBhEW
0eavlHLA4z1xKr7Eb4kYkC+SWEXmDERtkB5O4svqtHyenbFGvpCXcmGu2sg7s3QBQje59UEasiSv
wVnoeHQu7b6z6fPBZMqt81n5nhXs/tnMADTza3gWQeRRWUvBmvwAH3rCY4M0YZuYU4c3nZ/UFAl2
PiSPYQfYTZhWzc42jZWiq8sOYNqqZXFCQyetXVKtNrw9oOBKrN3syPBPHLyhhPf7DhlPhfkUeKCg
RZTKXXHuOcw4LCw13hYBUtjb79etXSxP5pI6pB1mwf/PHwZ6tRwV449DFMl5gKoaio5SvvfbziHC
5ZhdddsdZMLfCa0Nx2TZaoRXfXUc3kifSHyR3v7nq5+MWKL7dObqqkl8gJ8TzGJwDsxDKIdfIDV8
3MABqr/DO4mWPlT5jN0x3KXe+9H0R3UwKckc40jBAoBsRqN6Gi/9YjwoI4on7Suhaps5ZAe7ps+B
nWbZJynMTmYseVOkbjOobz+zMQ9i7ELJDm4jxLekmmPz4v4CrTJdMn5Ixs4d7pzOAk3FghQPNv54
n32EaU8S5OHF0ITGoInwzqnwAuwXj9nJ3qzN5GG2EaNfOEiO36Vjc6HW/DxaMjLRWdzyCDYJTI18
ey5kv+xhS+5OcJGOTjTNRmilQ9GwgTqnAGfzliahIQ2LCX3E6JbFe75qI8LOoWNaYRd5y1ZD3eUI
sYqbZqJeZ+enpAcA/k5pmR142C4k+KSufbNMOVeG9I61zJYePk7g9MTowCNOgBsyG8IZn/LYe1IG
DO6mjMMAZ0YA1y7jaRwv5Iz9LtL1sVJ9D/kO5B3dtrzbSeFdQOrdWVusHWLSP7MxC6GABBzPnVND
tthysvxm+CGP7vMVMER/2ZNvy3P+fZ5dGya4xrMIGL9kUpoURJPfem2CrDI8ZkSpz/nmBLLugKNw
KXzLggLxgXxlE4PpXRQLItMYXnmhzJ5WgDFKOske33DulQgAwqupyQ3//jrv8KtRgMPuUbD3Navl
by6AWK7SizESgEYFPmrnqvB23D2a1BylQjRF9528HdiF/S56zMnjPLmlnYcYvjJsODibDKtUFx++
msE6Hw9y6pUfiOAHLG9knJe28Zdj5lEUs7NG2pf1wPj8ZDDvHiWIXnyHCxmai7NXcs6GHCs9Mw5b
1ODC8mJiRyQm4uE4McBLZqWdvk+QCZDrly91J6Rf8ja2g661Fkrc93UA83zmN22EHAFn5RVXI7WB
gefS0RMuKbg5xCh9vHqVH2RmPxO0Xq7T4pkDKV7QjyxV9sp/lOeTpdx8HFyb1FjHHagotpzXP0iH
6BzkrVBtHEkjd6YF7VrVs/MLpQ4B77KcPwhwkBIUAAGpo/al1YrJCnYLCX5qt9FH63/zeRzurhw/
CQ2BeMTTAQc4cIxtMCFWJ7THeG7eaDtPAbXgbU2K4WOzcPZKTgJzwNIhwY0eXlqhk4fF/dJFPFxE
t9TalcIWbHIlPZjxNb1Ii2XUyPz+9h66SZ4o1yAy5YZ7UTjKNcCs0PvoS9xjKZwS3JR+kzLwsG/q
uexugEB9ZO+NBc+AOlPu09aYUKE5Zhn5Mg1il6ERtXftqlfCUWlMEZytkDsFt+rxbSaxz7N1XzNA
f0bjXsvX7CvZ1i1TVIMZtSP09cIDuoO2frafQoqyvFohnnQyX1G61ZhjREW0zBUg6pN1PhWbyRkf
wALPcS05HsVCHzw4MZDkzTZR6YAjIsGZIYrvnW9hPw85CBhgvpIyN6Gk1g4fkHmzmi0/PrdgCLnP
T2dE6N5CZh9zWJHpjCgKnr1rb6GT2hRH+oayzNtbJWd1dG/PqhKQjxTfo9woeE/Jgx5Nur3IqBAa
TrMq6AI4067BCpWtcJY+m2jhfbf3ZfsYB8v0HY62OLfHWQ0dFl7tOIUgmueJkG+dXNi9SyCJvqUC
DNs7JUJLnLVqBFrFgiEtXvRe8DdD33XIsNWe1XC6EweoYbw7cn+ZddWQ3ihZVKIYJoSwFlL5x478
PM42sRFbaisBEQAXraVWkRSCmfq5CS9kAI12iKZCYTxbcwAFrBB/nb0WXWBa0xNkIrd5NVuxT247
gJe6nOMBD4xZ6ZoKUN3kxiFbVdLgPf+Q1Z4Eyx0ozZGX+jhB6lb0D7bipcx6droApKMeAmw9s/TK
OFmRw+p8Stc9qqaHclZwl3rZKfoQnTheIRj5fSSXWnQqIVjcS0cAaxbkyt3COrz+aWKOvtu7FMTD
XRCX7m+lNN9sRLxgr1UqnM1piT0kbo0XgoRgeXniDzPr/ioERdfT6JsDOOcLS+5X7c0M6rS7/f6P
dAYSS9WkQGO1jAjW+WaWLDuywNqXPuwwkhRtwLyOL+WGcAfhN/5V6uVqxkNpOBAVmeyXNnDEe+wD
DdNnm0fTTm0AXHRj//sZEmSjOvr3EsMME4UdY7NJfdKubPf91sd0+fzbdOil3XlTkLajOPfqx09s
1o4O5QkjwVXEMwHAoLqXAb6JNaCY7LuZYKrWk+BUXKzbEEkJbdbptkccgxi+8JxhklLDwV5J6ElV
mvExx8oZ0HfQ+MIIUGITdc0GrnC2fFPHW0k2u1z1q1uMRjwXyp1WqaY/E63OY6zm5JR5yYt+uGTg
7JwIUp4Oh+DGkRkMAjBKL1GX81QEq0Go1eTeVX+T/8JYXyqWZVJuOvUbd+e4m/8YpxQGrAbanL2G
pKIDGN2Oi2t1l1mJrPFvvtsH72Hc6KUyccKhKe0TwIAg/upyPJADepOgrc2+Tm+DIY2uhpH9aQKp
0vcIXwBJ0P69IR6czJU8NwOWJY456txm2EmaB6cbVPYqwQGbxoO+m3oLjHH4/nSfMeYAvVvy0Taw
UbdzIXo5ZcRBCeE4+JSMSv77IVwMCJrZhbxbTiRyyA8Z7TlxfloXfCN1evIib+4Nsmk6rAWdEuf/
0xwVbVoiA+ISWweaM/N5FJt7yFE5sBbsiO3D+Cemf+MSdNypEH4xgtQllJTgtaheFFKzG2xNzPzM
dCwbJO0gYqGQav53QJ+75mXNr8QGahv1fhIn3n+Am2OBUbiY3b4/95dqT3Yb1igC+mmlixzDolDf
S6KthI3aVe+949OoZZD2nI9mq3HneZsstmfjoCoOiXJNhVuhlrySz6KrL37Q04vAiQrIiTCZyRgy
7zB5qGqJgGtQGY1ZoRzJSl3A/r93WIV8srWDmAKJASeMlKxVtsTcywm74M5kPl+f/WjhHJdjuaI1
V69NaUqZE0kHKAdGFll8Sodw6Y6fdKexQio7kXpoe8TBjAw208lpn76Jsx8kmwrrSP1P13CFQXxJ
/mTjZxvBYbpYsHuYcC4z+WkSuqdgvRkoFlK3qS7ayspqHEbXBQ2OJROlxUhttORs5xgicKuGEtuI
NENDt/N0t85Rw6Ev6TuZgS0A4HCcrKYtKrfm/tcRTJ9sTtG7enN+8X6fSo8uhiTLscWKgkepOGcg
64yU8RFsHmO8Cd7l1jGouHbmawdnsnRvUWc8GNugoudZkBoTF473cmmjYKdXQgNt2DZSy2riItaj
ldguY2qjVHOz6jrk1hP7iwgKyip3+801R7XpIFedND2Ci68ZfithnmyPiz5YQrB97b+fxDHDK+qz
UR4OHCzJND9Qm6660xeK7WX3yX9tGOLwHW63Wnttyz1Eo7JlMS1Eql03cIR7o9SYgqrjzZs2v8Jh
YuvrUteNUjrTi73+T9CPYNgQt8wHGxJytV3taKPYRHwITDtOBDNWRI7TULlMfpaGkEfObNUo9tEb
T4XaLPIS2Ga0xbYwYjlvZR6+MThj2mYje3/9nopIgDcuZG/vspcWrFAQn515EwH/rQDIiLiEx2RZ
bMbDPeWsQD3uqKtm/rMbbX3bxmTk8oaX4BF0I7MKIh4YWfuyy5eydQQpqlGUsAd/n9Ugs/lA7iFM
seimg9lUtPTBg1+LAgF9lug285Kp5QpjAobuq8Y1pDkVQTI2ndeax/w/6E+OPom+lnyctU9gMKje
mjN517eUOts56LK1ATKW8/qbwSsSrv0Oi4sK6dI0EqdSTi+4lIoj2o8B3G3wQFqDYvfUwX+Qyugx
tMA+wtzxguwmOmhLwjnT7NVwbsrbu3Gqx/t/Yal59aUNFF/vQabQ2x+e+R6RJ89IUTgFgP7XYhpX
hWZ3by+x1Cdc0pQZDWOVvzOR5Hx529D7/8z94aJXvzv9gtM/912KyUhPxxZ0gSZkcZ1lys2fAlCN
1OwgWYFPDFadeoPKof7mOjyAPwPHSulI/GO6Uuzlh7wBAmrbU9qaVAdTJlISw7KkcEh8D/MSKu4s
BvLM0qzvY14dxkP3V4+pwJ3CuTne578qG3FxSr6fhbq9BMFBIycoEZFfNH8nRCwP2cNRbiugHESu
48LrcdB/IeQx9J8QwQerQI2TRzqVWpS+5D1j9Z/XdBl6+9wp14Hrmc5ogzV8hLDpeQGW4bPMWeQH
X88v13jtnM+8VxKIUB1Ti1VbEkkQX5oYopTYREFzDHtJT9UwebprVCJ6SXcuhpgfM/lSQ89y1sgM
828Gdo8YKZJSIdIdxvvl9vKOAMxxigyZ8ioJt9rmAFpKDhHaqJdttqYZbbKo4zXvrOKO5kx7opwf
HTYAzed1ZTHbLhoBG+6sr/1RncD602DXkgxQBRC5zb92mQroykJ5eZTlnPT79ldN9A3E9lHmfqi2
k38NvuypAfuUVyL7EMkBkQA1vh1n6CrN2GT1QsgP2SYtZewYHPtxN1GjtE1fAininaQ66CA6mPNh
iT5SOtpLu2UaRFcH+JMsjLigutDtP9rUR55Ed+pfBzaH0UM5ixeyuHXTTaq7g4liAFmjpkRoszSI
nAjiFKMJ4PyRfBJKRx65lmk6/cmyBcxdQsmMN1qaXVKfoo5wiH2grduKiZ89rOFCknEotPEFVENK
586aFjTwaVR/+fHlJM8rtJTJas73r1qu78P6fjWYoD4i9JDK67NZnqyDK+b6Cg+eXCOCZbWuhjyn
BL8qobZVGZLnHSi5kK7KpOy8xIwcJD969m9VOD+ssWXzHIQjgIH1vDyetfayldg9OGln4aJBFbFt
xSZOdtes1n/cTMLMgs1hzdiByhetG8g+zDsLEkE61dLJfIwjN8nRJfPvGjt9dSB86Fu8M9Y1AZ8R
S33gKVDGBNKsJE2zT8gxD4Y7QOlh8diKg/lPyAOxMRU91d90LRxTjfzb3uAtqWIohGwUZ4ynFnLQ
ylgOQpbUd5ab5mGxNpHXbzhNoIrOg8mq3+heOZy1pWHYEdRxDknZpaJFrIAH4/IJfKrPtwZDsaU9
gU/tUe2vwdVZlD78hnFSpIprsbXvyd1J0Y+UVz+1NAOdAW7Yl5GvDg/3GGuPwyx91mGN9MXl0eRk
qmhsWoCKw8Aa5fnYMkOmG2fuGfqLqO6OYIB12yyOzhqb79oY/5yz5L4+jSpZ31M0fhwkt2L61km6
r8w4J/6iv8Qhycl2anKnPkCS3kYbamKCu/nDkCdEWipk996zs9iEAu6nY1H1xI0mOu0YDEKebsG3
c7YY2Ps9SVk5cgqqh6ME/3Q2J4zC4lrUKuZgGFMKZZKmpEF5otwL9jwIKV5h/idRzGazPtnf/IUC
hMExXGjqpwUcZpDQliIt97TBlyVcR8yHOf8LbDTwi1JvyiRJTkEJysyNHczv/M4ClLJDq8s04NoQ
/77m86eI+r/19RN3CN1lCdhej6S0SMkER2hJS86stYLrKwToUsj47Co1MCKsBxbtpFABWyxZO4ba
WDFPqwQwDY4ka6fWIZGMnF8gqRpblmy4x9Cws5DhRY2VxIEqMgBnzfLnnXhi6p6ScCyIohl6SZ0o
RqSbfoB2Hg7hWyttNQe8eS1frnCwgVh6g+o1e/F0l/vjBjd59tZ7u4hlmqphzA5AdTHRuQFlnx7y
3VmrNKWVW/Y3Ubs+2pW+hLzfYjSnD/wyA90rKpNwpkATcuOfRjMjkZWuEPXU5gNFZgV3WII5oJ0D
kVWoZQsB/X9pER6XoBxfXHjuskYY9CmVFpn2EI5AbKndQs4LMIOdudqRVCpbC+w5BSGMuLtBFFq2
J7xLVjByRCxGfOgmdeHeZpFs9tq1UcnWEK7OP05UsJH7CGwNz6ldmw7EaB2qu2+DlFXR4XjLjWZ3
u2zC33suX7vs225IedlgpYJGLCGba8pMZohSmuw1zT7CpHh1Am+rOKrvJGk5Kq1Xk4mWgZrm7ChD
ss+n8oF8Tb2VfAtQrL/5uueYJh9e6onfs9NtkoWayoohYSTiHw0GSuYFfZO6KYwRT1hrMqmmDGI2
2RVuS12xaTf7G0MFRotI9nnF0rXGWkIWzSSuu3wDjtYDWLbdMwTteV21KSxh8PENbzWeo9NlieKX
7CiGNyjZPyYlbY0G7tBUZSdpguP6RNEdAzHDGbeOXjUYWQJY7FTZEXkYQkkpL+tB6d6KttbEF2ud
6HUzSkGRQ40EkgCLQcxUYAxhD37QZ39D2xrVaagg4AQcz+SSnzMiOHTcoyZAvTlGgFO6d+cyfIGQ
DFEe5pF2hhsjpFxUfnzF+aHpnlASLJLVWizILN8HH1uNtGjZ2PN0G5JDkz+v99cJ7XIPwev3EkUD
AJQ8r6MsTgyOZ4WIYh2GWSeVXw2wY5h8OqIh6GeUMnYbPEWb4QvKCAiiaGC/JGQa5KUFHCz5I9cc
IB8hmEBCh/CBrBV2AjGVtmaGqtPTA8SKIo5CLWQK8FEyexJES4jJ8v7NIUuQEjTiuVMYcDx5WJci
ctZ0q20LR+1bn9MebLRM5ER5M/UCYjwov7Gf6ux67XriGQUqpSlV+YLPu+NP6MQDl4fKJj8KLy/1
a6OLUY8BJ5MdlyJVXmPO+hp8KB8A946RKp0LFapmhF0g1zuJSUZqVHJoWpnKvpgZX7KBRe3kqa0W
iM/AEjRK9tP4IxhD8eiZf11gdQfBgwXNY7tQ0x7YoaNiy+mNF3twjiVS8+rpxMEkbpx/KN3FXfIQ
Mw6p81QiVf63waLo6uvM0TCKpPw5pETAMamHsIottftqfUblLGj+tyPjCCiow0/mm8wjzDaTG+E9
PVpnLiTcPmd+cAoeNKbcG2HeUa0/gzDgxpJ/vJtHkinDbellnbhnM5bynPW07/8nvc60LtvZgFUm
rStqQEiY4mT3E97qUjC+iY5CWG2K96P9m1AEIYtAWLL6+tI9dqBZXAxp2DUAmLZV3jNdYk3Dq8vS
6QHaH26HgQvTwLb7SJaz3+/2uc2ypXcSqB/QxAhbQx6n8FpBmgjeCHrDjlL7kleDm+MZ1lonSe9W
YDR1MTolYpCGMMco0Zff0cReHg757Ps3xx5/BHVGslPY8xS1b0RROr9218JwIFzemEhzcMJPyMCL
Xq28x6Q//mh+hu6irXRw/9NF62J6bYdZh24yNaOJbEMreIZgp8n38107722ll5F0DZQw5K+kIQa+
cYbmpjKAVY/W4cNAIQM7o7mR1BjFbQEFV/VOin3mYaOj+9OzY8k+FlN5idXf84oVWqTPEd6l9Zi3
HfkWlu8KR75NV97EwClGJciTbpcS59O9XD1ZBk5Y3rOtJlli7/X9a8tAXQe/1yuEJikek1gYGBrd
6M6JkiE6ZPjMrhRNcenQ7qNiVGo5+iEh2kaPfMSsqKLcumA9VxJBGFSMO/eOpgGi40gGMvPk7Sal
M843loxJe7cMgWuNE1FiLGEuRP9fVkKq4FOQR5lIZiekhWeSgauN3mt6LlBVhKgpRoCwXUzi82lv
6E/BGOF+7RbOShpSCNVFKcY1Wxnzd0U7lp5kdAx3LBtB2RXP9iw//UKKccISIfb2WedhZPwiHG8E
Gzr/nqUtKfDCuPt4dKqwdBUWO02Rt/1VQkiLiH8L2JZZVowyh1UwNjGB5EOWWliM9KLG6KgnuIX7
NtI00+XFNQg4WQZnrAmesO5ooWJ5IfJ4tkR9pwj54+EITDWdU2d6cHMr437kR3DC2wwEmBZPjk3T
oKcVPXfBTS+6oUBbwwqChw595Ejkf/XhlPyq6E7bKFpfD/GfC+YkcYvCmqeZrO97HXIu9KU7Kwbq
b9HKjfKR79f7BykT0H5gxx8HRFF2GXg3duLhx3cSuowGXWNAmwVazmY2QTwV6FFrgi0eFNhZjfiW
E81jU2f/jMD2/YjUHxU4erwMSnfwkvSfWvnN8E+aKSn5gvRHZeReRcS1R7+vJwsEGaOyO4M0QmS7
t3uc5iO5WXZRDSgqrgtz6hs7uvIGH0lwQoJLpLnmx3KNyrpE1sHQQFT9vMRSdAvbsIKY4UinxFQZ
lvYZayK/tEJ95tuBJtc9p0xHb5KkyXegy/ujAXECPxUSn57KUyAvKEBk0KOOSMjQfmGZiCQU8jyg
yu/sYg5vhyCwgu5ZASjGxJOPpoJG+g/95fn8Sj+k241gbdhR6Xuceod3DyqW2E81zoC6cGuBjmiD
Pd7qgBI3wXOjNZI5P/mT7nH6iCXkS4jz9o0456ShFPE7kkDOJCCBishY5HKvlPkYFRAwNNoaYozW
CSmkwkXASDjpnnO/7jytGwlF1UxhKVm8vIZCowenoZJQt/fZSTJWVfjhWZ9W4ppELlDOUyrLCqz0
WcVI617rJX4a1pHH/QFfTzEdfb2XKeEKoml7+TXrQ/HABHfg/jVFDprzNAOHywJ94+7FA26c62Qt
WO3u7w6fuHGWNCqRCvDj6ZD87qKiAxFl5rPxEYblo0klr7l0HWjRoak8iGQDcHSSx2sfMNyknWG+
JwoBYiXoZ+nHitIagHGnqy5crKCXenlNzJc2mE80XrbtaY4EVCknYGnyJMD7dBVb1Uw8OsLso0kk
WW90Tb/pKWMl+qOwCpTVjOfUEUDrzh28ON6go+QkWzh/9NEcCHH3omphZQPd3Afe+cD1kTCnfRpK
FJzguiPbxtOrgFiwDzK16ZCDyAI5ZjqEAbr8lCXkh9x9K0q7MZX4WinA8anihgduTEb9oKGDWZKn
3gCFkh+8gvCeqGTG5yL0vb+Z1jkQziHh8nG7Ef4w3RcjQLJ8VuJQK4qrpqV6fT7bEjeu8pGBghe5
6hjsNirZ9QzOB6hUAlDuvTkZ/6thwqjN+mfI9kwwCXgL3JKZoQHhK4IEpfFiKTsL2dhVEO5vk0r+
MiIB2CDopGRfC5jQteDCxOsZ1V+TPzXPOiMKAqMSG92hjCX/vBHcHBX86mbeatf8N+P0ROofZmzw
JTh7ww7TATk+fiCh0s9/hRfslE/MLZXZrHvqmVpxl6qeRVaWvA9+xiV0q/yxpSP0SQAmY5yNXQkG
THrzGFQI787qLMjfXBHAImlwV8PIm4zBgqG4OjiFHY6fKsNwhiuq0UrVYz/7FU8bw+QKzB21MTTO
0kTtFiAWkD/9V57uks74fN47PcyD/SwtTrgeWyCBW2m+lJThaX2uRuN/EfrpX7n0mP+UBnpvsBLf
5XjXIUPzb0Skcquxiu14FzrELTJh2KJwz0ZIJGLUYLMfUHA4EEv+SRAJHE344tDZr4a1u43w7xXt
vZYKaNg7hOqgxY7AhYEsGD3xuUUpo6AsWcMYcbWp0uXHoFv7vQQcqTgaWsIAvO30qExaWjz24OOa
s3eFYRQxE2rf+EQzoe2o4m20A8N/3yjRcORBw5nNWBOLBRVgj+NvQfg6o8W5r4qn3B8XeMQ885M3
e1V98MkjoYOnHGUfZaac0Kcn86AZFsTtpbRPN6NfmDrQ4upsOBjxxTCQED1poob0aIOS4JrNAyTU
isWHjOAw1q0fQXQIAk0AwUHJVCVTW7TyHwTZb8QlBj7Ax1lEv8g6RWOV+A44at9l9Y5l2Gzj2Cmy
Z2h5BDzAFvGByLsvlhPpNqPRi3zVuzIVZWtXcjFaHbuaSNdj6AZHrMHJB9dpyr6hpwZ+yrKx9ciu
NoVwu3iao1fy26XJ74XlYYdFF8+sAGGH/eC7yvOkf1usWUAaHVqPXHdvndTHvOPUF1ngqpuBgVVk
X42vA8Q2f5NAN5vk105qkshjPWoax+Syr5ZAS7JuElW3SeD4Oi1cHM/NWIuBgoW6P4C8BhqyOCcI
2vDzRhul1oa6guLxvwZY/mXvcTl82w5YBm5YNmsEbmGVhmUpgp7ttX5tkg+BJPKPkpbBFPzpXsXA
af/+yrgRHYRt9a24eU8y3GS1On6+bMJqr9h630HEHnYYJefZr032IClMmwXh95fvKTfz6xOb1B5g
2gA5khqq9zaRjM1ofb71Es2Vl6P8fKeH1zy30riP459TFXo6pxmiFtwi/pdv3QoHs5Wuy7G1OVFB
zQQvT1UTSzh69rkVfjDmBF6UTH+HZy0WmybcVG4h33d4iSih07TWmMds0JE3fsMMZwUtzcVij5n1
c6ynlhatSWg/IPp420+sn+JLCNYBhFVuN5Lctn6v0dPW+ksZE4CYhbayuU5EsPg5rtIz4RUuv/Cp
VLct6jPXLHAPpvD6sP9E63X2igb2RGaWk5DN1n31WkQeXMSxIau1G49E7Fn0qpPvFRVMcgSzUU6F
UzSlb14VJrVuPEcsDuORGiQ2QTzZdsG8eHD6Vc3Zw7PIA0V3RX6L8rA4aXCXN7Bi1Dya7JyLHgzw
0ncIlgqfyOI0cHbFoo8sU8Sd59LrnDc32ddxu0v9AkGufC+SMqSCW9AnLN3XN4NHz3TH5hJJkC2F
9EI5RBXtTgZu55zH2e6VYlKEtAX+ZbxbEY3DrC2nY6KoSXcB3APV+FPpZvtzxhgTGFzvosLirlvi
3zd/dQMZblOp5W37RRa0kK2AibTef2CKhnx4bzq/102WKdPzBuOYyMWm3r0SjL4Su06aI4U0HVHN
LhgQw33pnAWmDr8/pdaSYSgx6oM6lqdiVX0qXNOeyh1GL8MQT78pme9+ae6h2I4mggoj3PAOg9h+
vScB7wXJ4CzPzNZQR9aTibAj+ozsT1efg38SzZMFtkA9ID/yZIqZeZxtp1+BJZ+gxzdmTxqFFEFU
cxRC2/SVaxUpjolqqHJG+qbES88lhq2JGV+0w4+RBn5AfZyWSk5ncHJ+jTcyahjIsOjviC8dGPAr
zfmzhG7Krxf0+3UHPKYohIOdbJAbsolqvpD5J7hiYO2KkeVdR6y7tTSwu74Rfgrh/PvBFedPtkRh
hCaZ2V8ROIM8z3lplyqRxqy1BC4+LlRLvcxm+xh6OiindvRLf8fIHmvEwq3EPYWY1JfsMsw2wLh+
1p+x/nZ7wKVSaIk9nJylCcvA5mG6kyWIgy2lgqflYFABCoGPVXTbpOKlXxjEOVjScD0oH/qDSGUM
V3/fBZsJZyYrPh34zCVAu6yfW/SNxRL9vTPCJAQJ1Y9M3lT7N2UOB3DBnLtE2Yr1iDQFAT7uSDb8
qiF5dHTgZJulA7UgZX9hcv2aycJ3fyCj50DRl7TZdaYMOxJLOXNYjXo32+2I7Z8rcXKSY36fTCsG
5XkEepz1P2iRTdo1vgv93fX9keobZDQPgoXgsDqa0DV16WM6L/Wjs5qgaySRS8yp4bqMpEmlOePV
+Z00GiXeebo5XkD6IQmQOVtpwli0kelFSv9uwrAVpGDjJRx7B+pPskSauzrcXhRU+LVSHPegE6Wy
KCSf+R+z2p4B0EtzWD9m4OI3ymJstlyRVDGBMa82fTWhwz7HVMsVB8YFmnmL5HJErByffPs8Lniw
GPbAdfT12GW0EAi4UyFpaVOg8hVWW3UcQFquwDewGNabVaF+PwmxkDZUcGcnKdS8lUVrwhv5YcKA
IcNyxP6KOIB5bpqjWZLWU/ehWQfUxX/5nuquRIUvdI6+baqDtfb/Ec8QdtL7ojnSuzjAoXN8ei5/
dyp9sQ6Cr/WgaCDw3Sfe8k8Adv4wMs/QmfTbO3+LUIE0SXgeEVn0tfD80hpsIgRwyLU6izymFygi
PK2R7yJ4Y4gLzmkWnzog5O2H3DJl20Y0Z1Rk4KJCWdC29VZkinidFgM5u+pRY+1YkcyQJW8V0rsU
tdh4eKvvW19RNPeU0Dn/JBw6nObWQ1kgqqsZuUU4I0sI/Xj5uMOcXH3HyB8t4J42spSBxlYdS31w
kgndGda8yYpAb0aLyMDxm2c3ZCoBy6nIN0Q7JV+9U9QM/+w37fnQcffU+y+RYfZFmjpfoUGTYEBQ
TLIYLNIL83jk9ULXBZ4y+G6kofcxouaAO/VZ1XRNGrnzIS1ds8q571x1Q39PwRKH/fV6oIGPbL2j
E4zBeixCmO1Z2pN06XfPKK+qjEiepL2jYDvji2YGxx+ySnfFwMo2Qyk94uk56OqDHbYJ8TyGCWU3
CXgwgS/2WNqF8qsPH1hZ4b+W0MB6XZBr1/tBTNVbjDQ+Mse1EQUsI4WJI+x9vt0HnkrjlNWmcckR
OYg1fMeg8lyHG0Tfyl6HVCVl1ZbLl6mCHOF/Os79A9ruO5e+y5L6UoGEavnkx4PhyyCuyAGgaSp3
x03yK+/x7DR2Bq97fGXjoXAZmB3psQ13W3NVFEz/AgWx6f4tUB9uEKUKT831RaSeQShiTGn7HzsF
PAEQfRlmt5ckm0bd6sdAzoRaQNxMSSGfJp5if+fxIHsQyzG8qh6YURUPHfQd6c+Q9IXdhxxqWlaX
QHookSB3I6HsVeISXy76S9wVFZ8diFk4Nb+dG8m4qLcrqWkPuVj3Un3rH1s8Dptz7sBAws3hgro4
LVgcgIxKcqJrWDYfHLdvmy1XjmVsmTomXAQtdhrg7jsLMzoG0nqrmLmdLdv+SuY+cHUykwGouLID
HUAAklQdavr/MgwdenQdhOSK4h8VMN5QE2jfzIRF40+XTPmKNmcXiasWNdCScIhKdz+dIco+HR7D
gGt9oHtFQsma/ctKXPisYjfMHQ2YrRQZZlQAHlBXn/7lSBWSr2Kk/X3GHwT6q7Fclb9GKEuhKyHC
jFHaG/XCGrwY0uscy+otQyeay1H/6aVLPyeupTYfZKRI2Ei3uXILNtzLy4src2IMjCGWuGBu63yl
kC8CmafEp/kkxPFzWpmidWdPVV8pM4VowYgr1mksdolb7hKCYUty3bvvj4iMXFLoUeBbYG3nKOXG
b5uPSmHaGR9FmY+4cjQ8M7+Nr4bbx3J0i0I3GfC1qZuXt3kEuluI/TZiXQFyiXnMXfvRAneS+2s/
4yteP6VXuCzLtNBNhtqIoCiVXTKTcD9Aij3bZUFLCw3gn0bQ6HCqMsqm0HOn/V1DqIe+3lCu7W8I
AqIspzUQBcNBqw+v032oMxYbyp9XpytPyqK4/pq8WbFYfLSruiF967wMqTzrk1UkBrz5DcnDUqiu
PIFuYXS72tZlkUbexL7D5ZTVZeQ+2nMI97cKfzC7KweNQyQapIcNElhD0UviCuv9nftSiAMARLKm
/N8DLDCKlXha9UOnF7+tA3NqHvDIyY9aryNayxV6+PZWJVagsfw5JmxAS4YVyK7PwrDsix6dnkyV
+C9KTPMulkJBj42ofN63P7CKj9aDX3MPKbiDv3KWnqA0aI6L5p22JK2QLrDQBwwbV1GwnQn9tM4y
jl8lQx6PWStNtc6x1MW0sve4gSdQAyFXsecIqCjE0AZrejPPXt463b3XK2j+21wQhYsZJJgvS3xk
8cHr07VHGz5uHPovauf4H5N0eNaita8m1RLonsBAaPOa6rP9jTrnY6p2DS398/HR84w/wOxSQzdg
nQARiEwW4/zJvcND2XviJ5s/7OV6G/d+dBcLTuOOzmvcuwuIo5tRgWzy0zYbiPgoo4m37ZmyMANr
CqSaJI0xkJn0JUV0CTdExlaWAKGkycJKGjPUZvVCAQVmi3uZMj0WWgUPaHJfn50d2rTTg+dlK1O3
G4RuGxRpe4fvFa8Vd6DCJmYfu9LD0HYR6MDFOKiL25ehGkhXNJZUSoKgPLF9Zk+FQBg1IBVqRrUd
Xnc8alOH8xHAnykQoYIe5sh/tO2KeMkavVl9bbL7wCu4m6ZgzA+YOx6XaQRxV6AhalvUZNoCOHdw
ADgtYZy6rD6ay6C47Q61IvooGiJoe2YJdezKeUGNImKHOY0QuxNxchriX3ywFEuPCPdRabQBjB2J
H+OD1x4PSE70J7WDGFebQkctaK7OimNz4kIT2uzUK7ES+//5daM2EWyDm0BTdAP/XjIPI8s87cFV
1whhcZnj5da6DckSstmmIKQsmpDiBkWJMmeSRFdNnNLZEbnNiW6atM98pu7jqz5LswIdIRyCLp+h
WFhyGt2ByWzAuuPkvIvUpxl8KCEX2tq+6tlLZoDEhj51ABG3hvI6Plcf6Qt+ISJEfRhvnqIZSHef
72O6X4xr/Uk63OrYEIp5SP4CNxIG6WSF8p58gR77YPDSOQAHNgH8BF8SVsOqnt9Uz2LH1mlM0BOM
tpEIIsgbu1JWBsoC4UUmd+jMJZf4Ek/eC2/eFgbpLzRrx16FCnkVYStd0KxAgHsFiv+VSftKecIu
beUt70g9bqz4L1QLOX4I6iceHJREAOut83TykT8TIL32bbS/CxrnFbJ7X4Wof75JJTWFvbwTgaC2
og3TJF+bWSFWcrzLLhRS6NMub2nfJU5Ab8MHezbzclobr7jgAcZqCj5HBhdcbJ8IUwTx9X903RhW
J2wCHH1TvRN0/OeovQ417IO1oZKpBLREH6uXYXf9XbmGlnD3up3wTrqjdQUOvp/nG5ftHDhTjm0n
kA++oF5btVmfozkVgQLM4EvrZUihB2Zoai823KG7nuCFAancw2YTUtQokbKj78k5cmP9hdxbERQQ
HWMmI/+YUaKESxGf7AWcKw/RxxPiTiQ/GoW5zWFW7Lofy4dcW569K3A8wJJiAcEfl2Hmxb3stmtX
il8fZnJwzVwfVEWGxrXNlw03BpuvFA5Rpa7LADrtIC/aM4ocbJqg+mqWHLYQoxMPQfqvtwstYW1o
16xk7YU73mMSKyGdp3x/Gc5Nm1qqIqAg6iPRRwzWHX27ySaQkG/GWshD/fH5mCiYQ4eWcZlNliVU
eV6RdtfUYZcr092HogLo5H4pUh6ggtRFbUlswNhyRkACXkPQGD7qc+GWk8X3jfQtbDOB8ksDBjrp
7Za/P8fFEuGGw2cDJgEDcvShyecflfxG5PQBXfbHz/M0AKXra1JG7XINB90hH0W4qefNaSnuru8e
D6jZexzsYOY6oRSlFVviEatbDs94v5siJwR0sl+CKnrVW//IAM4S5ByHX+7CG4sMvK4KTgAuDcl2
nhkqVTtYMXbuijqIAw7OeVX21VFedloF/JAi9cvSSO7yn2X/Q+zKTIHW0jRoRkcVTOxIezGTJXC4
Im8tuBYfx4AkL4VU6RDJrYlAyb5DTw7UsGIj7Pjlc89gzsvHuz6XuqtD5m+un/4Gr3t5q3UcyEuQ
UL8QORLe3Hou7yjTDvSg3+6seeDshIYm2us4eBM+QJXMpCBvqVpLgJwa2Nw1XDMpHdfq9cJmWsoI
tl9N21YXpO3C1fqzE2UqGJqYuJlB7fGfx1pt5ZoZkI1HhnYzXRJ084UwdjhCZPDgPO3J1XCU6nph
6+lZUBI2DeCzIlaRL1Bq19G4h4ri5+b8TeMyrAmjGKLVTlxSN0PPMSXnj74N7EsxqWKsJ7/d0YqU
lt4ho2ApsoQEqfNrzuVJQ4Diygq4MvRv9xKCIrGxguU4qYw7w5bIGzuFb9e3bwTvrs+mQwqwc6RG
c9WOnzaDz2ZT82T4MSVUxtqU/Jak9GM9qRduIVbGGuabLaZ6rDasC995L7s8TLXJmZ2MAl/ldmKN
g7RPGM+oC+jFLveoMgNUvbbQlEXWm6x353vN8KpXt2bwucWVP49vaEJZBaRY4EGZXu2S4YoHyWdj
nAF3FaqnuIvtpYOvdI/By6NXeIAPEc5VIbj5fmIiQfk0abFwph0tr6TUdq4R1Y4Y4wjFSUAg2cZ+
OW0MKw0617qk04JxuRKgUr3JppDtwyGFUvCrRR/3O7eNh6r+MechaMRYCijj6sMb1u8BcBofnl69
kq5wqFBRvyjJK3VM4lR/7NQECDi9As2pnLLaO455gJgclJb9SWRa67KIaDHFEI3Xmzb70wcoJX7g
S9auUyKRvglPdBQgyaGFFjRMtanrE02x12rYrGqi5n2rorwBbf0kRZqHhXlZm1olgmi5ID2M/C9d
bePDcEKwhfcySggC6jde55SgAfGqh9gA+Xj+eI5cEs//hgkAlZOaqCg+gXXgpXXZhjcVcj4I79GA
9smf1/51O1jKMJu1xQ6OXR3FwzU4+OpeSHq/KLIu+g+qcaHJ+S2h3oR6jBFe5BJ+XdNI47xX0RDI
8KZj7tdkHolpyJH2OBUwEBxeyqs+GiEt7bFNwvjpVAvGkRdgktp7Ftr7tast6otpR2lnU9s5Dph2
1ZdOYAHLsyXIOpCpf4ZQxImO6urn8JIatFrCz4RgRyTy0aLaWAS5KKHUKzPueLguNInqNR7uTqcL
EkWlM2Y30JqL8KIf02GUo/i5anvptWgZccFmZMCcPgHDYVR3ODxzBf0MYfH09JSIcKRBEcDOQ4f2
qmlavLfw5rUywI858ed8cEzk7M475icMcNZMqxlBjpl48DwipHQYdPrBDcV7gHOmbQzbFgILJ+bf
s0ZfB7ossG+4zuw39mhxcA3PSDvaVW8O9QU/IPU+74pWXbBDXkM0KQHHmX8wTcF8Tfd98xGOgWDr
mMf1ZBBJb7ekOUN8BHCfNEfPVTZGm8AUckl/zOajX6PVl3X4iJMiIfi1gUiRbihB/wwzw4EGnpnL
wKBhqT3FZogZZIFWu+dwyX2t/55R7tMR9XaPv8ZzftDCNCp/IdH5kgxRYuQoTEaSlET1YnfAX+uj
nmLOAMmpX9Q4KLQOFWYIFYzcIU7dloTi/jmcBspiWgJAriVCR87UJ7KGGyU1ObfX8CUEVxCHBHr7
U9ZP/0yFPuq9HPLZQG7hZWyWVecz8d3HAg0mdRPmA7yCjV6SEJkpcAji6LvH6x791wgTqqt4X4Ni
y8ZQFbCjyGtksPEPWOUCsV2Mq4xCWrp+6SlD+wCkwjLmXVXd2QhSS6CJdsXnmjyN4V4quuDdUPBb
rbj7V9C4g0nPcbmxy1+XrpGazqAnM16Wpa6NhyQv+YFAQ5Qj8uz5+A/ca+oSd5TRRoBJ8tz3pFL9
gDHQH7H1wd8d844kf+p4rASefoHSTTfENQ7iSYjicIXoj2y33E4uLRxO0yF+LsF+uhJxrfW7BolM
dUxJb3D2GW9+NYfwZJ1vd4mGmtPrgulAZpfJZ5iYWD+UTVnF2gYRtCM10y/sUrM6W4tcjobyKLyv
Py+PO5cWfSoPTLwWEhmKvAXTfvm7bkjFZ6QWfNGioe9o1jyZLpxkIsjzcz20XQAKlxvwDzSLCUnb
eS7JYITbscfiUKYHsNAQ78ReHWxLgnNuLGirOkHMIZUP8Q8hVDnYyP3qsoVanPXsHL35GersOEpg
ny1t0T8yFe87OIxIjo2dNLH66dLoyCPEdIaSf7smgKRu0ESThILCc5S//iliqQuSKG2PmYmij9se
nTeuSvRoOaNYHxVCNjUpc+sDZc6XjMZ9q+Xc6Q80rClsHk+9IUcQLEpZz8F1hjH7243qzbJzQgeU
7g9HbR/BZ8esKH+q5lddLC4ke95uGyFJoktnUi0EYwlHtX1dX46NKLaHgU3wObQieTYr1byFbP3g
SN1Fe9CGaCxy3//byQQSwZwKO3EszQSKDlMx2451gtcsQ/Tn6qPoM9yq/ENOlMRwpr672H/B61Cq
rzgbTM1wvgnjTilDva9ei7NSYFSJ2W1nHEzxZGkaPbiQTlGT+S3T2L7KyYrClgzeH7H9xVIBE53S
voeSrE1/Hfv9AjE3TvXH1ZatrebvFPTaqWiB6BX5wCpCFsIeqObFswDynw1Gya1bfFrspbeHISiQ
JbjQWewnyPGrvnb1uKJl6NbBBXCEiJdoGNZQIxZQrBLcPSJjtfFK17t4iRHZPnrSwGALw4aGLqC6
vn6bi2nrUsOzV/EzAuXkAwUPyaL5WEUppVfbbl5+f3qffQXuAdkRDmFitQpQjG9AzV8VQ99hF3Wp
JSfPrubqWjW8UNmYwpNcClBe8bBSKQlvmuS74UtNDxxxSo/9TN3DSl4peO88jYYjGZGC1F9UFhVE
JBt+73L6n7bOl5Y4okm3qudyVNgajhOpjVYCkduUeYcUQb29FTeFX6bO1TNDmYxAvlTP8WqSXYb8
R6/UdEvLzKGIZ41HOPEcHMQiSa1+byDRTNCqYL1H3pJTFGxzoHK1LVNWiArtHFAA6cNmfXAG0DN2
FnmSNJdU3vQriq7Jb3pzMBNai1+AvfQUte79+lgGKgE/mpnHIyJTQ6Sh3M5QJjbpQcX+V2oY54UI
t5tRUrbUHINyrblUsYEqq9hrAA12j4moVAe98+slnDUpfrnvlLWJkNvJE290k/RXKvbrTX8Ts+e+
+O9UlSIiO9PUYLAMHDjU6HU+SveDGOhQ1KLWchJ7NN7gFN8DUZpXjJ9cUQq6zDp7MJt7p0ptUVN6
BxDHjvI8roopB5lK1jYzOsvCFELOVNbDzicqDC2FBuM2vWqrxQ2TAPgs/JkvLdJnBKU65bTfXpN0
WVfrQ2psojJGl93XVrUlSG6mN+ZXByOvDvAKm3e4JLEpHZ0+Oy1hl4KCg3akoL5wYff1I9tPSY9o
lyxRDOvC/PVM0/aFcbMMwCHT56dwzLkAXg9B8vN0NO1n85mS3Zt905tV251bxvZO+CQXIwYHJZiT
+Ju+CCH7v6TF8kJp/HclP+WYWtXkOgLkls1Dq9QJ8fwJL/x6iXkuN/MwL53sxyRrCGFo6UbQgWYM
VoFDFY7ACYfxKH7Ah+aBp4E37zGfNkLMRSvpRTFEdkLXxBf3l7HJnLJO+lQNTirBmgpAQzZSdg4w
AVJuhwAeW2OW2SUM/WngUZdH24c7ozISOLpmNdF0gkuIeE97heOQGraBl5S6FliIobx9x5SeJEtp
wVuxv5Lsmct9IdGWkIuZUba86vj8OlCnhf3Evzfsa3WUcbJH4c4FVvLUAEjkoXA5FGvO9JcKK3va
4gw8oX5gXhg6HOP/nU0R6F3a4XHCcWC6NNs3TT4vJuC0b8Ekq99F14GDkwhj263Xb6J4ht1mWtIW
Bwcgw3X6R54IgfzXhh2JFVlXf8ulAvpbFUVhOQcaqLyOtsHt9iXG6xJwO2eeOexJRSWDOGTEDw6K
NAPT3XWdSAC1h5icR/Oe+lmsru91rSY0qsqcKl42eJCMf/rJTyvb/PeJXDEofxsZRtuVmOTSqoBi
P4gE4bVm4DezMEQhWEUMSsfjWm9ohjBt3klYflrLxp5ZxnGTSa4/XBAJnRMy1OhHU/sHLAGsGXAb
jTn7SdwDgVwkncVsoD7LyZ5gorKc5UH7/zcWeS1snJTPARt+SnUjhTeUqKP4RJKstQea6kK4d2YI
/S/ta78TnK0UWbBiABI3cN8SHQ7UgjS6+yurwGvjowF/X3bd4A8JiUBqS9iC6SEXtXCPx++4VFdD
terK40aTmuHPNAME+u17Hj8p+NZmtSzEj+crqklaDNpk+imCBLHImsx/N5uPTUszzHUd6/J+EP0c
mq7J2/7qLXmRtQNXxTFUzPxAvKyCqdBdGAMTXGioT3DoCh808kRyzztT7vNa7dcyB5MwWBB90QWC
NUx3/pSG7nkzmFcgJiTOT2zmWYF4CxuVWxVprrQtuV4xvW3GtnFw5ENSOabCe6Z9T+Tg/R+OBTYt
0zj/Q6aM0xMS2D9DzjjnpiTHY9pTGgy6JiBjcdlDHpqCQcqhEe/iitpaTQQ8G7wPsaGTuxwXHLFN
Wr2cwKNa/VuRV7p0gJuibI5s4nqnXnvF8fzPFBMvCd+SEE3LFvikYApepoKRMti+wQw9wxpVFLZn
ImjYkWhJWp8tw2QRwWAWNroID/elHzQHaReo1MTd0fblRF01rfCJO21n1tNVOJQLTZ2Liz86+kFW
JJcY6Y8SMCPFNmq5KCkoNu7F3+WSpQfYjYkxh2Aqou9AHH/BFzMPE3az4z3mN/XBuV9PeMjLNdoq
L4YhBFzTiXSAn3cD+4haSKTHf9aCzJmuKgFf2CcO1xXRi1Ao8+LPR6KMEA0YefoWXoDW2mw6GEUN
ErlsHkazkHUG9YL/eII2Fa4KNOL9xoQctnV1vwHokMpbRzMl/NZy+vf7b3DdtEXAEg5EUwNFNp9J
18e0ca5CoU/CddacmpgYJ58mjKgOrhaZce6+t2DrwgqN9nFVcWBHvcrrRuheds2HEcON5ew8hCTm
UUfr1UoaAZ4kaxn+ZK21OJEYPhB/IHVnKKhdaSJQxKuX1ulwZ4kLKee9PyajM38+gR7ocVpPw2zS
wPvm/e5lvz6gNb+wCXGYpkplp+Ry4H6pwNUZUdzkdDNAY1a9ZIqeEb51DsX8FtO+TWcmR6zuS0Vu
98zPCrRbCj2j/VtCmb32Q/ELCnY4aIPgYNe8tMNPcUkYBwzy08b3beXn6Iz5PNnV5OCRFE9TcRid
Bi5xh9qLxcbxc2AXDctiBcLP7a6H1NFlggTjngVGWY9Tm1hpaAmww/zGNUd5Oljsi+473QKaunpn
jRMgIuhHpxm9qSW2cT0Ub020Xw9jWAaWQwtyzp4REm39I6XwcTov0MF54ks1Re8lABw8iZ/PmcCS
jctn6CGp9iiJXeZhsabITpHKSiEtlk/sB2If4/XsWPGtab4WQ0ZqeHxnVYaNHvDXkPsF+mvtTqkS
5pEdxBLaKo9CXkAJrD1W0sTtaw19gIJqg4x+VukS2xnXr6adNFA5OaUS9NYntqez9EIcE5ySu+DM
GnNInAKAVwuY7I7Y8YgKaZRP85r4fNNHwXCzTbBpNHICYVGb9J6BUYlPOllwzka9+/fQI8luRsqR
TN/5lRzyWX66JbcQfIhteRRJXbh8mT2K1/rkrTI6tAS/x/KrdmOzo1ZxmVSdbt5J7KpKbnwnIbD4
1opo0uvnZiuvfruuvZRlv0AGQTuZt+51XfhKn4zxkuB7Zc4VFSb/uQ+h7Sp2J5mFLk4I/jNdCZl2
jPvZOaK8/ywCgWSKHBoWEdknlCDl11wgACaLeADJdkaPnbubREpJqYTWoDuuVAEmR7ToLV/0vG6m
WlMRpu53aPH1j8EKMFm0BVIlNBe6Q573zVEXRHq5RAc/WnmO6OnNXjHLoKuETXh3qE2Xk/OHHkZf
E3w01qw1ANVALmEat97DSIib+Pb70XStyx+fE3ChkLCZjaYj4uoH7C/4Xu0zea7m11PdiftzGAu4
DkZTWHPPsAVgBIko7QUzTj/e1xRN2J0kkFYcdDz26KAM/Zf0+iGYpzcUGzZSWAaemJykIJyZ/mua
3XBUbZPg4pwM9yFV4iTlykY92duHWPzboHsDe3ApnM2PQRh8Pndkn6aJB+KHM1y05rFV43TGeWqV
ObWb5dwvSc7UKCacd6/b4hjuwmszuMkHWq8iNdvZ5+TBpWUdjoMhzu5Ek/CI/jshWHRStqnQRv+3
5LlH+yrrttscYtfOk8YXAskb1LsQQApFIzDJ6V+huDvKA8sQ9+QMQGnJG1N+Kb5lNj1oua2ePszx
6MSPEw9FRTgZTr0RmyuiDYBLvZoSA1dZ3UNyXnbR5wZNHaNxRX6cCYC5wb02DHTcjTY3Kq6LGe7Q
zX861SgXxRDrHHOITCvLogaS/59G5qrtaaVni45erEcpSarxKKmO7NF3tXG6liY6DFcmEMNEvpU3
f/OV6QHVhwuST0CJWI+2PW5+Pij3x2B7cwEa3PYCHkuhxxKTtEofVLmYeti6QRjbApH7CCiFAIvZ
Q2t5IsiwpyV/dDwWqcSJsE5X9dssPHsCqx+2aruc3mXRI3T4hXan4JAQrwmIxPjPaUvlHD5YUZps
f4V9wHyxs9cnpqmcqlUpjEMI51r1bb2xZG/xVzruzDjWlc1BcCEC9TYox5h1Ni8AXlHOK/dSY6vf
HYfJRPenLlor7pnCoHesthkaCUohn8zRInTjBPXKOPJL/dEnQzxW9uZYr0/gEIGdtIPEVkGN7FZu
kbU2dqxcu/RJvUAu7opjIa4tI6YyY7r0CWQR5FeAl7p8zfbUpOEN327ZnZWK6FxeG+doT7apq1Lj
4Z0JV1UnOF0mAEtSjyjK1FkHCJlRIIKrKf3/ft3gRg9GJW8cdNvMfDu1DbsdgqmeRpYDbKUWYheT
UJktUx6ppeVhiY4ahQa55j3WAPgCO5XxTDJRZi6X7IpgHJvuEB2pMgT634q6J2kZut8m7Yn+4z2l
LGkDTwnOI93d/KvN7yaAGMjEpmi4+1ohVGACq6XPRZ6/TBjfyC3aZay233gQ4lETYhjB0pxfXhBn
ZW8RROC/fWCT+vOfLRbHfhWG2+aSMIGuS2oH+0xsD+nS+IRPa/qBXNYp3S8LMCzZ9IPIgxnZIyjk
a6UxQ4cdG1/s9Qqgft8Zsf0cyJii0QWWhk9wu6R889/Z18Qxb9fvcPwddAw/PlqPZDRUzYrdVQL1
7GY8dPkvUOg4/hDT9pAdEAL0ynrVy+1kc/lZuq6WnxjDN7cwDgfAboQp4+y85VMXoX56rrm8fAEY
zECCndFZkZuxhEMfJvTzBdKvblgBMPW0YI08KhCXJAAou6MNf8JgqUg8on5I/al+kiKvgdlrC34p
YnzcRbWNu3ZgO3JQ7PajcNh0v0MKiGqHFp/pk+rfxdehVYlRH7yjo1l2FyhBNE6HAf+XRq8FDXxe
hOf+mhvO7P7umBluN7vbnLBeswk5gr0b45ZlUt1p6m8lofJk7x9hQpqXgcF6JkOnGl8GwJvvbHOY
ln076GVUiKbyMD/Cjsdlt3Qa15XJVGxdO9VO91bCNE9WoEFAzocCJt6+SPVmGHav/mcZThSDjarW
1XSqH/YyZRW+E4IZptTwCBK5liyxmlWZjqa7+uf6tvo8+sBN1Q+CoGt+Jvu86xdHNaYpV6yuwFsZ
YnDyhCa7Ccv39qNorhUMXechMsmkyB1veCJC05WfJ+qg4tUq7Vo+xJVPBKmO3NU7LZhntpEc3ics
90rVCf+XkUQ5j7ry4XrZh+keW3mCGz85FYkWbHRUe9UtcVKjzJdWqD5KVvvRImkZZsrc5kZzODvT
xq0qvVljKusUJMlPz8cR9dPeo5muuBXtq/gQuTOg0egNZ4mq8VH4Brl75B4EokRoxrW7MxOjasZq
bt5jwdSFhF49gkDpWCd9PSWwNULkOQvE6XgGgqj+9GTgpME/BwbMEeQUcSo6LkDtDfIYwgJXxbVp
2Y/tGXbxwQ/aj2MOGaTJ7Pux61V1u01F2UxvHXeBoqseiL5EuPSXlEA2anF8I95/l4h31zECGBdM
k3Q2D5dG5P93uBkUyviCpDtx+PfFa0PFUEjlo9fdbGOksTxAJbN9wYMtZjcSmiJwqNuJmFRdshC7
SPS9F5bHBOPKCxEcWfMqrRRiGVVJUc7fgKGTZD5JQWN62tZiCI9xdMSlGiOEN3TbyBWxZp3xl6Nr
9bJOgTLwToX/RFnzHafsJhENhKrn6i0lz/a+gZeCy9kADkzgBTeaQcf2h2RZ/a66FM1F7zRLV0GK
84HP7IVnfcVOey7qlBwtav9cFxHINzdW04NMbruzyW2eYjYJHSOMdV5nv9bhjW8Eg935SNW9zQJi
PNIR3Ry2aH0zotIWxjwUe9z4w7icawvj0AmuQdVM9tcQBPc4HWGVGucH4jY0LWbAQykXXWhwx9sL
GspYZlMILU2IhIuTRLECro5oVIcyxzKXbqXGGlcZV36HcFccxi5agCMs+2Yngo+7YZ7hZjxJygAp
WcRH69BABmtSLL/nruY0FIK4EAd7Pvr3OL2WIr1oTbderUaXfoRVzjihBqwrZGS9fmUqKyDhc5m+
eK0CgLFju/Z3iK2dwMcPGahjfLQ26gYrmxCajtMYib9mpR5v5wbRhn4TWjof6v3lu4dO1KpcE7Zj
Dclq+XWZCGjR/oqbg12XcVxD9Bw4a719K3jTsQy88CQOXw5/qwa0VpzUHbHaZ+19BdC0O7jY4xge
Pz/B/NiCPRB3iWUGkPRJpG1YYpl0nbwBOscvOEn9Eqj5au/h9vNRwV87NQgUM/UMJPnFpnppFp3/
fSvaiGfciQbbtHddv9FNENPTJMWbVdeNbGtiVSHP9RgsPRr64G3SUi5hrNw71OCEhSq3/C405a2n
0BRzzsVporT9IPmwVbd190fL6OvUwi5G6niUz5tgcu+6a08fMb42YqEwRqxSlVRLu6ZSTOJqzzef
niKmxE0TXTw1CGZd4kXWMfqX8pr2DOED05EXWXHEyImJOZNFjg5xUpMOMj/iRbDhCUoSEyzehSRv
twjC5cpR5gSDBDba28DU+dvvYnbYjeIp7pQCF6DO+GIIcdoWggsg1VfUqd5o/+8C7qIF37knPASn
ZkmLLkh0X0PqpVO6YTAX6ZzfCmEF6dT6WlwOqc6An+TbeN7TFuv9LawGW89Hqru99hlBZLaMx5Fq
abwHAGnEeDFXnbOo9X57vv9sNn9OKGtATepXyjafrPPsS2+QmfivNhN+uXBz7h68QOzufg5IZ0YS
h4yQgpi0Bi3nAkTq1q11WYulWmJhsZui5bxytUjd0dcNs6KvGm+72FRabqLfAvktD4lcWmNHoCQl
z8YjhsAu/J+Z1EfIYBXgBU/3Y4L663w5t0JUH+61nUKlHF9T8IRJKI3/aj0dbArm8PXNOGuK1JQr
xH1bdufD9YLaTc+6RjFqO4YN9arxL76/iXSldOM64VYtf/cmkaWgV62XGlrLxd0JlkiyeNC315F0
eQfGDlxwlbY0U+SNB2NEp/0ydkpbChVJhYxIeQyixldLiMyT0LscTlMEQ4aAkQyDWVCZbGf1PsE8
2qrkcj31eGLXEOUTxWS2A77LpBxZXLzLvwnWvhVFkTqPDoryXnTh+AKEvr9pS9+VSv26muKz5qQu
6qc+iAtio/6d9bdOkislLe55TMReZqYvWH7iyOR8USvsu/pCjOwq34tuR1n3YG3zvDFIQs45Vl9/
dWvyZ01wBKq+wF0y85d/q0P7MUjjZM/WH3Jx1qEUPSaGedZM20Z+LMDKuwRU/qRdMwc0HFHD3QzI
D3CxJNVt9N5LMqRVNVwbtADgghpZGZaE5oUA23QnjzLelxkDN02ycivBZweqnGZT/+xF/GAWIxj1
QfpyU36aOQicxUNEkw5WkA5sEYOLR6znAP2gHj020oxv4gMwvn05Sf/xRHLIDpo9QZT2qsfcDLIZ
MZigBSLc3QXmsjkEfwItixWGfWMh+VWGxLDU7ncTSlnBDodEggacrmkJWxdI+bCnvNnSvBa2jO+q
4s0pqfqnMv6D0MS7Cd9r1Y0FtzStVHQp0ScbNotq2zztKusGdFiYIezqWXIQbckHhpZcdwqSi+aA
LgtZgHP7xvq0TJbZsa2CP6BbkQ9v0ASIdOL0nGXuIq2aGbz/FVk4b4KC3b0HB60w2C91zZwhpNBv
0Nopf9L0ruzjj10wsCa3pjpd9ATVBvXdlM8eLxgOZUk/EePVELARzHb84zNi6KPqPDKQNs7Zr0+1
545unCmeSRrztZ8nAHxRwPbvH8KH0VJeKgV7yat0CjloWTefHJknG2xOdSbrz5ha7k6/2Qk1D75b
7HhrqHLVXEnLzu60YsG+r86DNLEQC3Vlp+UWouYBTOIWG2zg4i7FYziHFhHaPAB7QCQr0FWpQI0a
itEMx5ZehsfjrWos1Fk19uanephQJdKociQ+bJLoGgTRspy0OIyiKPizjLyf3JiWBFA+g4Kwhtfw
PtPwQ0LSpSoroTMaJh0/5pkWV7cJV1bBlM49FFD4JGbCo/8rT7E6GuwmzO7dTdRDU8Iq9IhLpLVI
O5v/eqLFd+GwNyzrJcvTJxORyt6aBdT06RG3lDolVfw0nhx4gh5YjcgCySU2kmOrUll3RdKX30gp
YaSygW94ogJ5npRACN0V9/VSGBRcwLYdPlul6O8k5MH1GscKRuWLIwITBPGWdDRQmnu+CxVq5qsb
7KRyBk/caWy9E8tkORCPQtGIn85b7APclh8UcHG3LUQP94+muGw8aPFPbwR4AEIEw34ugqdjiSUq
XyYGOfhN1/Vm9hLLSNd2wof1yxFXNG5904PJjK5z/cWAWadqCITD21XXjmHwHffK37MRLfHszZoL
4mzD6jfqMfd0iw7B/FvtOzD5lBn9sPOwQ1MpptNxXvcmv/Rn1SziKD6hylMHb2fqrc9/Ikea80t6
jx6NsqVA6/HypMKKRFvUVFZ0rhpeLOtRDPQYSthFkaaFV41KmGlsYO6oDw8G9xeEpYRkca1rgHay
yk57VZY+xlGmHNUqYJbar2wVJyCeB3NW0UZNgUvMwPZF7ZnvwSiduzzkSqeNWwv0HMwRhwZvyexD
F8xHRmPwQecDhwLFEGTZUuQDjqRap+gVHIDIeN+UOMN9zFr3qnbynuR/ora/y43iQnYiGwKQiyN7
YrGrgdkdAYhd4gyqIOeeFxMDggP4NTo0DK+yTOAA2r3ieqhNWzgxNrkiYHPQziWjvNnReKzhoQS/
SSYabcRRLZVgZj+naI8wAZW0Ac7TsB6+kNl5DVuUU9ELyOD+qaUoDW/nb/s2ZeEeE7jyjQi8Fsa/
Ak4Ps/9mQ64k2/mIfu+wnDileGezrOWog9svXy4qWs+rupLIlNN1dLZ58XIzcRsZSU8W7IFTtlQo
aDVCB9C/KoXKeuMIuCgHz2kTGyvn59zELse7hchi2NmfWeW6qk1EoLyQhtVgKqg/0ywmYb9yzDsd
qxdHbCKpaaa0tk/+s6SZEDXHdG2OFWfTN6N6jPz1f1ERriRjPX90ZQfs64OIZNPn83cyWd/9asei
JXHiAiteJPem4urAZHdCtgjlQVtrtCyMyRUm4awA0vFqqhwQjjJy51WvdjfiHSjwdiVXuJxRB+JS
NV1EheemlS2yyCqPf0dNfLMIAXyNBbY3jybBrG+4caimaxzyaylbi7wJc/4r2eu2CAvj3ZD8biW/
wZjEs3exmE5iPiAG/hINHoMO6f5avV2D7GwwCJDLQPQz8O+IVKECSv3/xXy0Pne4sH4Szeb9ngT7
qQRK84fwubHvtZKdoN9kcaikx+ah+Dx3eTig29mcfO9+6MuzRpt4aebZlRsSr8DGD3m/YFqRPGM3
3T08MpgsBQBFdI7Jv4vlxxAPKeilgUhAYoEf5SUIqhePAw3rIXduSFGgrJHOPI2Yv/W92cdTBD5G
A+MnzbvQSbwMiFozw2sxhn6lopma9B2Ey1IzgI5v/hw/SnLXEyee8KWHRsMu3gtPEld1+vJ2WAvb
MkJl3Gu0yokKgj2LjnCXlAI5n0/hPWGQj9rJYDz9eDxQ9q8aySPG+9+bCkrpMqoejgN5Ojtdq1+8
irifYd/oyycLbRhxsLSHRlA5ZUZiR9D2lV4c9wtyYQ4KvYDfQvfnUC8UisYnQGG2Zx0gGIByYC0j
gD10hxVuacvhmU8HaU3I1A3Ue8DfGpI8TJBdw8AuR7Pce/ZulkzDxTHnU0QwsOKnyTvk+s5wXx0Y
B7VIRvnx9ymcNBujQR89tcJur7XRpAwNysIHN7xZqQg5M/Gs3jiNyGKeKNJL2KQs82frjJ8Cxc+n
zbhpQRppZKpnpjjJFIuygPO+q1KNyjTivg18NahVQ50A5iJXIuuOOnLLfbes1PYddvGH/b56385S
XykkAT9OnkwnLcNgZ9y6L830BWU60mJbrBpO5S1MjFvJhPvZBWFM+PbsbvXOd0XWd09xIBFMJBr5
qifPdg5G5+n3vExzgD3kOlN66HGbnOqAh2D0QeJafrySxBnOSNdEBE22sVlABK6yd1ZhbXDTux2v
6jrmsdMA7s1KKL0Jsz7XouS0Q/v/PmpZLg4r8eEqRevBbFg4ar2+KlBTKRVjdyrEC1qW2pddm9m4
KzhqnzFyqNSb0+RJmuQ/tv9A3JeTQPVlhU24OVfRP5iir4aAB96F082VHEMVM5udh7hM3p7Df708
Cy5N/clNkHWvDEke1H3rCx0o+iQElu/bVJPkqe7YLK1sypWUEKzIuybOldn1gn4MHgjJu8Vqg2gr
7wxvLdpYPX52x86kGRHvxsjVvqT7d0ZOxz+d0kq99w5nxWK++/dqnEOpOz0hpElhcdZ/ujlfUQpB
bVPk6g+xcxO07rUZ8dgkAjoT7A57Fx2NDyYXS1+RTmscp1fAvnM61P2x9NAMxPkT3l+Wc+4LYJHf
DjCfqlYqnTyW5appjt2ZLnLt5iAHvnWc1vkvMwJspV6PzooyTcNh4cJ79lkLmt7n57aW0t3TBXyj
VLSl75tyDblX+7pLY1dsEtYMaEgboqrUMUifjurUD5eFmBiWeY7FudqYXKYjNoJvfUDuY4ib7srw
S8M24T4fxNqG1OYZ4m8G9H3kGtLcL8EH957BkGIxH/Q7HFPXzGCpkum1GfhJ7N0NzRd8g35fmdYY
BeLb7GWXsMMo8/h8uH0stdCSoet7T2QTuHMnFKCrDjAa8Dc13w1TIie6cKBVBrEmklByBqD1oIsa
2WJj6I9mtIuMWtD8Faajto76atUhddGWUWEqGTMPHYOIvPNXVHb30ID6tSABzlg37TLmN8NCe1IZ
pQfpI8yhA29ZA29Zuyrpsnbe4ie+Tbg/SxH7BoiEtfrC/iPJMEGr4y3RSXtXgzOpNsTKJQhCtCxb
LOYk60Y69QxZfFZhLjtbOI5D1NcZPCQogfmKNK/564Uw3RXyvBhFA0sGz5AEhHqU2nQjp016kMs8
3kXKmbZ3eZ/bq3gleZYd6gXspBjgzysnQc8qaigehfSZcYHQu+r0vg3TQnXIFYnkesBLANU3KwpA
skeTlHtDnz5W/5iLvLYtB41PaIo3XEADPVZvyOOkVurVU7N3PTw3uax/CVY4xuRCF8ml04TQwnhM
BPM8jv2gUmvtTI7DJv8vsoPCZW1I3V2RlMNwNE280ssk/nI4o5AYU9kI75XzagKxDBsfFb/gnO4p
7GFHKLCgIEkjb8hqLR8e1tWdnL3dq2jWt0BgggNoBJ8NMz82vGvG5gWLskpTFnzXjfQ8CAWPBa6A
IMXwOU4vRg2W3ewEqXLPoDuBXKQBSeDuoecPiE6FGssvmorCqnpwgxAueThdOjjUmZAzi/joe0s1
xn+tX8ys5C6Enf8Q/CqUvN3p0XlIot8PeB0ymdpPrNLgWmmQfWbOb7Lzu+gtcgjsrGO/bXF1cl5V
qlCQoZ23v7f1waANMHTrTQbz6RS6DSzux3pxnPLbtEpgDit0JYzyeiPgr9XwqfkEMsI4RQOIZtOa
X1f32k63Veci5v4zJKn/Y5+X/XzGtL43g51jVq2WkSFImePODCbuNc8S2S4Q2/2ghFNGGfAFaTzQ
LeQpw7s/RElPtJgssTwNT206A1ATrNtw2CZdykMA3LXFRohm9Sya3WY5X25yy26gz1SFaebUzWUY
KQMZrcT8c/Fd2928HElk/kRn0SAI06LAAjYi4ofd76YIjUjh1WL+SdyHTVyh/vFS2VSl9yqFPBUB
i846q3VUV74AAy/4+30bOsjNMGwXz/HJ1JwVK76t/Bfax//chWAuTn0KXbfKRPlzcGq0MMfMjw82
++Yc+REjWwFOHBX5xBkzbZ4MHN57SwKJhAWs7PchGTeRYrz9ukPZ4R8At8rcZk9VQziJHA4db4DC
j5FWoBTQD0cq7iaBEBPcxsBOVtK1Rckv1dShMP0QkeU5QwOacjDBNy8cOw2DAtBbqqnxiQ0lUqP1
BqwQiP0Qg8v+c5D+L5GYH14W4cZmitAzvrf9LinGKKlz6w4yi0mpeutDHsoysvMIbdfBb5dPTEtj
QJQxvSPBHyldvp/idjzgkCA0lKzEDxVe346QllIg6EgUvhVrzR6y1IjRp2wQrJuZVVHii2nWRacU
2WoLlqKZ+0VEAE+Ffr9/rsLp3SRo3YedOrVV2BZBuHrFa2LTJhReg5aZV3f0zVN18H3buTExvDqI
fvJfi8Kf8FW+3CKtr4bOdB4fmD49BxzVZrmfVPaDRxPVE/IHXyXFqJHmfm/hcBAJM37yqZXmyGED
A0N610JBazPk3LDrrTKZD5OEvXcCw8s3EjBqwPqg413pURwO+TCw/cue74eGHXUKkM8MygCITcQN
zkc5ukX8f+XJ0JB5Z5cU3at0gIwrF7UPB3F04FEUmXELVi5Dvf+yJv2FrC/jcXSU3dGJ3SygZclb
Zjjeu54oSemK2CGImtzAkYjC62yyPtN7LudPv529G7dOCKL0m7t1hJBCJf2Szysf26/LMj20kwgt
oIbUiOUjqA2Y+KxGhnZYszA1otLX0hHJjnbQsn77QyqE1P5YRT0KvcznXSBx3eKQrU4DhxVRJH1d
/9erWT56GhQJrTnsor3HhVabnMnWRUgkvUnB5LpsKwkrikC3/F4n3/pCa3vKsocfO6aD4Fo8yEzA
h+9nRY3zyB84n7V6OrzBiWm3JREPZ+gTiabHs6TQI/+eYuLES94AaXFVjki2HKBRuuLUSa71/lFR
xEz509gZxVGWxvvcomd4vFSD9eMFgtN83mYoBzSB3U8GtTxxGZ4twMtJ0xIjopwDlgJuFoLS5nD3
y5nGdsQvu+Aex/8Y6xb3edSBfyalP0Qh4VCcTv8DIGZC9ZLj/FhIZ6DRGOY7iQcut80aHpuVaPL6
kXFiJATn6qYiuzUWFc3RLdu/gcE+OFGK6kqytmeAX/WdRihtc9oKnD4xn+zXf8JM0XaS0LNnHyDN
1ATmRznm7bhElwmTHlSBSLpPfgHO8cS4qjcpI47lqbCflxinVvvr2gHZ8K4IvABd1XFwgCnLOek9
yDGYrYxyCfODQjQXGSctDAAL0/aVGbiup15+REs6Sc3E2C/zeBxEhRUqKJuvNiQO/6CQBsxKwHEh
AEMxI1QlmRCfS3XQj7tm5esP5Y29HIsyxCWiA2Kmu3kVu+W/3l/1hIA8kL8UETdL3Lm5YtMXzt2M
KuIq2i8APY4kkT1QnPusdHLaIHFnFrdDbJzDGjagw7TZv9kyd2G4CXC4TXbiPxNLDKbak+oXRGnU
y37IqHau0GK3ItEV3zKXu6Nx3cqHG6LX1xxbTYSoNV4gg1jl8Aokr0qQ35dbTsBXCnnahgmTGTVM
BFvkhwPpgV05SmkRCgwYKoWA4AQiHKpc8NMw6g1lfvNwTwQLB4s4JcVuIIv9nDN1Zo7Fvl5soaLj
tdwOtR0Ge9pPgrZWsMcnLT5E3Ek1jYDksmbmWqHr/iK4y8o3odg9zMtmMHFqq2V3herTFbgKJ0FN
YZ0GXx8L4DVaqFkI0/nGQ9E+sY+1Eya/sMJVAfTuLo3fSmTlDepJophOuOZ1Ooy8wlqnvRFttBBA
guToT3LIDC6yG6bIAa1TxqECl1Q3tTDndkuWf05na9xKBpYKZAtzkzATXHAD647KDxYyQp1h42Di
JYiBnXi+wtNv/fYSy+ajtRcghaHsRp4sRRvwcOGqik7Itc3dbnclHCs8UAOCwlEg7+HlY6Eyw4lP
00g/2gASbiIr+8Usey9u6+zZCpWcquLLzgepZIABxNPP6aqKvrIvZO2VRi2oB8L3eHVo2hhgUv/X
Q/KBm29Z/HK84GzTCyUYLWE2nPVXZyx4B0ZwMjMu2+PXruK6Z6yt81Uhx718nmdu+pIcN480yVBR
aBxZz4ZHy6UzoyV+DArIHCb/PurWgzRFgbNg/DWRFp1HbapE3thL+yJmysk/wojK0s0GS/oIauSk
X+tD/6wraJRYXB5m0YLgJ+t/CHweESNkuVsyewLYok5Zn1ycOeRpoOLDdxoHe6ojhBZWIpNK8pzd
uDQkTQbHxRrNqHhEJfinDIxXVcWZyu/Q3cese3Th5qR2fSHcLDpPj3y8ZDMEp3oWOOo0NetadO12
FNb5GxW/zm1m9Z7tw9epEdc3Uc1l8fLMpJTHMIrwI7WRbui7yh8AQLEL0sPAkx90DaNhDmRwQWGJ
hZJeCv6lteuZtBHcE16tO3vTQ1mTGuKEBSZMEdkzTmAzbmFteMG3+l/yp4EgHZUgLwXIpnsmurcD
PoItOIWs26T5Jjf3yBuwOYYGwPfqczw71za/nJU1XE68mVvgOTwX7us12QR4k03dUGFD8kYiy6Pq
xvbbDb6aXEME4lbrykh2R2mqdA6BAjRpatcVm6akjP+VVsjW4OJk0RdrMtHg+rTctN1MzdGm/A1S
fVwoCVFkiqkY3P6VUGxD2gNMgWOu20GYpsPwowWQrwC+m21iF8Yng1YrjrhMJtr3L/04iPyRTRO8
mEQKAo6VbBK2QeDBtq8j5N5Gy0cm74+lBd9TXxaTShUZjBX9woXA1QCoSn4YV7YvL9A2LFUNq3q+
OVdg6ZtfxgrnS1JFUEYYpp/m4DlypVnTmX3u7zKKVAMStEausZWuD4zvgQ0O+hNOwysT4L77DFqJ
VeiuYKWOsQM5Jdh3vRsI9yQjYjmc2GZiAGii0DtGOdvZvrC5Nr/flrRbu9fxk9eR71pMzh1qf8bC
tWT8/jHX5mSRD28cuLqgKeRTP8AqzXPX24InL/d2aSJgYkPNYTHwNgnhNdwhIDZPKcexMl8IKGB6
IZrVaxpQaIlAyA746N2Rwk24b84mmv+QNIHuAeYLLD5KwZJrDgyd/6utwLrrUpZVgA6SEMKgSi1P
Jp+Oo/A3be3KWwI5/mt2mIuvIlS4IxVBhU7K5yepsKqXc9SxSPOt+fgO6W2xRZr/B59b7MWie9uP
jSwX+mTOVVCEIv4hIXBbJAuTxIRx5xZ8V10XUHlmCynw778GsPn3J11/8qb6/nvCIrf/tQL1ChfS
X/Oh0BYguaa+1PPkzdk9K0vHv5K3VepsV1HJKasyCLQ0AlsrUeJpAvsKzCiWMU7B8qCvDizyTxOc
QkVvGCVFCyGuvUVslXluW8A2o1JJ4G72wk7ycWJNvbviW0KRmcZ86Pf46HVExSbHJoKDsvkjVCak
5iC6kAzdGCzbX77GTOtlDvlGlHyviDrqlwHv17a6TqGncYHkKFlvW3RJuYXYIcW71zqkAhALwg73
k883p36RjwfQdCP46jdcaIbnv71bZ0PiJf1LrHh2eCj7mcsvgeDiSBcGDPqEYdIL7i7Y28UFNb8x
BGBbMwIqshcxz0S/qtl9r1V2yW6740iuYZZfvyuar4HV6xAfaoEcqt2SpIaCR88uXmWP40DKAxfI
O4S8jVCbAvNso94bpw2RbuSdbUiTcA3XBKompJynJERM/Lt/zoT3if9VekoTIzOzeFNTdaLP6XDo
w676GqP+ThZUZvEhqyyrrVu1EC8rHAYtxUkPfkBIXp2+y6yOJSlL9/SO/9cIHScEDCwgfOxlzn7L
R10RutQZpfZaIh3HQGeyalKCMbjqZodRMyyFhSNUoeVC3e5+qk+F/ac27quhnvgsuKaCi+yDo4Pq
pJQs7Ztma0lNcLIgVNUWEkn3vCHvB0zn3ULsfAe4fZ6a16mFZIhjFI1Iu+w3RU9Z7spTjBxGcuIw
mQvVpnFeGya0Gqof2d45453KazeZu2wL1txs16naEON+H4QsarIdYdQox3UVxxkQpXLOQAwKK3Cv
bdWatNT1GlX9vshfx8ZcvD4vwelWnwYaqCrVHjd9yG+SDUXyi0VXviySsSlayj5X9M9V473tnghw
JNFxR8csw4TCRGhGCF+Kz7cCGyAhQdsUs+wkCBh7ru0xxIT8jp2F87/macwyeXF1MdPvhu6nR45Y
D8OZzMhTIY/ExJBRCeiWkAqRijMw6faDe1dsrWvAv5rNfOAODu7YjQ72quVWavsWlg03548ybJ7w
F2asEmiRYmXzks4O288kPJ7MUTcDSu1EAYy/kitsk7Zx+hG6mc1v47hEcCOCc8qytmySP5wiqDSk
mlhcD7FPOZho+tMXEWiHmUm1KZClyNpBsTnEd+23YQZwBFjEUP7Sjdd5OzuKTFOdbjVAhFr0SDD0
4NGurlXca/XWxltx8IdEOYT/Hegovb6nEjxMhd2EOm3ILBixAMb5CUMVoX0UD7mQeC5yXL76nlRh
GZvT0U6TAachHcQnUwR08EsaB4ECEmG0qljbB4cmNxTlo6y4RokVB4dh+oItREziQOAr1GbII15e
woGsGGrA2AZly2wMxg/wVqrYZ4clgicf525jdEu5aSeB/oyfOidOjv873ohntUKKJ2ee2NrBS9Hx
glIxJI0D+pSJYmdZFdBXGNtu8KtWJ2DAypI4s6ykP+GR+JbXaEvFiqRnkP15Yt+H/Mwp+mD5ecmF
SxTLlh+c+9VGdoWM4R4bA4FmybhVgbujR/Hu5yokCUaeMZU32+VSQ9MRQd/YG3tSMbCg1GtcgR5v
DZHYiP2ZvDz2CADwEJP0CMfIy3dGrVGRKF8VZeTGozbchC/BW/5D9/HXYjChaZtP4K5Kj57gvCMb
lRfYAUjJwgDFP8APe9gipGVOwLqh1QBvDZSTylyJh5q+cAwODIHZ1vEBbQsf9jBvjJlgb/21ZDIL
Lyg211XBi//fr13Qf9EM0Fti6S0KRmZaFTLCk2xPvPSU0x4RzdmVG9nrIl99O7FjkY8xXa0RqaTx
yqBImQpTsZhLLDEvzB/RzIZ0KND/2H+R/z96bdXrdwBwTVeHXQdfwlbcQoO7r0vfnz0d8oWTVYH2
scRDdRwRmXZC+gQ9rcVZBKwaaiQ183/1i8w4OU5GmcUByoG6QoA/QHhPt/iD44aYA/8NxlE6KCRE
PIPg49bZFxqenN1Knh4Dy16UKfZJ2T3Z1DadrY0Akvq72rGPWdp23+QJiu7B7ySjgkBUG4g/ruep
vcVbg+U4+j9LkWxZ8mq6dV06TCIwKIardEMgSQeqqxXSSzweroeYNuWTNNh+SV1EVPt4oJJCvvE/
KdDOIc/ci4AaOE4BnOLcDpKK7+t36EPQtlq+OgquTtaiOPuuBjBxqf7V20dJBo+vvj7ZzyrmOLH8
ShQSCEkeo3o8tGOToLzDjPwXfUGx9KTCI8cBfSOlvDNMVLHj20Kl5q8mf0pNIYi2Pm4KdzCNgKbP
ud6B4C1NTaN+6cfpPKxSgFsi/xcSGg5ikOkGUo8rzNewTfbE3hbKYCYccqXgw3kTOaN/+DQa6pRq
09/eRYed2+in0aD5eUHdMp+mf5v93jPBRfsEngZzDRY3nkZe0i6RFcQUgI1aYIrFjDcVne0+RJHT
tfhZBu5N8hdqLcZMdJBZkguPhkF16xbdFAMy68IPgFmll+13s05FTEKYqUC/uQbWAwVHu18lahKM
GVPgvy3nAF6za84tazJ0kZBelrlgdrDLeD0fxt4kzyL6kyOkKYQ3u1nq0oMGMpXc5HiPcNs1YrcH
TG78JOoZ05dWtBcIWJmgq+QTxIxRhStKkO6Bgw/J4QETCQU6JcmR1v22maWvCpVRbkTlMm5aS1nq
yo1UvrYE/H5sTRUP1gsxaA2ljeqgAwGtTRqJ4nu3g8TRt0Ikq0fzs7OHX4g7cH0aS/EGZUEbewNI
aYxziMvX1XzIjrYVjoVErWRqei5VUvDY7hjkv6SDbQ/aU6t0Lc39YiDw7NQmUym9Xh2uoipF8V7U
jtFX+8cbffp0Ia32SO4apfTkoDgkeE6ZWbvk24VNd2ENX2QLbm1GdV9UTRKDL14OCx7W+kbwOltB
wjQNBy11u2Zim5I1ZKAWVSV+HzfYYDbr8zvAP1Zh+rkq7DHjvctyDclHiSJmFs0GPaek68sIp7MB
uU+yAxgFlxBG+RrEU4JtZ6g1R4SuC2LISpXgxDi50s24UlfeQ+vYL2rwb6TNcHS6FSDbbZMblCYi
bZKVlS0FBrpR937bsg3uSBmmE/+1MlTJxm8jb63XqSNgLGUjwc1rM0zxzqGN1PTe11vlwT/Jf+Nt
uT7tOm5PdPawsTE4AzUcOwhVsMayOKBqxvlhwLQsCORSTi/KA19CfzjUIE17yCk9UwKe/SF565i2
mHYbDmtVQRXpBcRoURqxUjKSUmmBOk/rDYXnceFpvqV9zwtBP/SCgoTlIuJmFMQGUCNX94+hf5Sm
l5DTsrQ1S1JMm5MZxJTK0GkdImVu2Sg0NWdOuDpqqgAV53Rx0KBT+x5Ds8oHecrJ+pXC3t9Nde/N
NShX2/OJFwkSZpmcJCIAWF6wW39PiNFveQIrpPOY4mPM4vojlVZcRePchdkg7HGVhWo1Mrmh+j8H
rhWH7VpIuzgI4yY+jRfj5M1Sm2duAyCDPHriMjPW424sKI/frP8F0hJkXoXt9vCWcTOfzCBOrjXF
OnW3SQCK+k+rD4hrO43TaHAEtja8tD2NXPE3wxEhonRvCdhXRJQ9g6dLy1FMm02tx6yqQugdAsEx
NIr/TPnsPpql9TusR65TqpXFfHp08LMOUxXVouZXyIdA1VxxM95/q2fgijeQKy7aqsfkURLoaGu4
WnuURRbNHI/XQUhYzmfyo8Ty6vJ28soBa7wCXxyoNAJmdLYj83yT3D2TwPVZIiuW+N/r31wIvtuX
UJotRvsuKjKeP396ruiJc2vrxTnLZquTdimgGEc/UwZ6WLaTsSOGs8r5WMsJ7zJnekBA5pfpQ0c1
XqIh7JpGZ5C+G+ZKPJ1J8IENt60iv9XSCM3Tnuy64uzoOx+3iBOT2QsBOK17hvibeP++W7k3jYMK
VdIochbxwPe+u/eWC1M+IETf39SFq+nIonCKxRXvSvxwI6h0Oc3gWsov70m1IndckY/Zaha9UrUQ
b66Svo/PQ7AV5opBPGHdZ6Yb9JGH40FfZ4zRjNu8P6ua82UV9J+cu75AQuMMSpEvtYLb3IzoSEub
2yxgQmy8C7Qc0DJ9VtGCETUoaiwItOWGCf6yNj88IOPEbGQuKIWxsmEw2x6qy3X+toiYdIiice2t
T+uWxZmT8/px37jlN1zhjCphKVwG5k4Qk7uu6UnG1gljBG1/Jmu8WrCY7kxOKOIwXSLZ0pzx15Ca
Sk5yzNOm8GKkQE7h3pje/vchUBjgnOXwfINRppId0RaazdqaS5oPW8AiDO+nGV10Fw3+hnWao+VG
cqPvSTk8VDwetO6PiQ5qNIh7wf1T3UgidnxrAcQ8dXZf3PUEffiem6Tx2YwRna570CHTBPpvK5O1
vpwg4ga6Ol8gsXvCxp8tzvQT87gdJ/wN8S0zHA8YOLABFPkMDa0ykv2pmMEpjmF4yCL1euaIa1ij
W/jahn9kz9tGZi/4ygfCSILPTo4ZiD1N4A/vT6QxU+NkqRvFzpRCGAxZG81G96FYp9M0m5/+vBVC
/nMYB5A72Pf6n0ph4DsHSEtVPVYbQh3QbGYRQguea3cVlpkI188SeTaquLO5v3wzI7yz8j7J82pM
RVBIG01VuOLXzFKef8G5ZwX0kUNmpGM1xwhnaJjp6ihk6Nb6p1yJhD1s++alih2NHvqCH3gV6axp
1nLK11uItW0+ySGsEffLSCo/v4+IjytHU/i3jXkIRGjCvvPfWBZNwm7yPN6w16N4YaNQ9j09QzBf
lRc2jyAkCKIDx94i+9E08QbVtbDOrq86Kx61Xwr9KRjj3MpgTyl9qyXaN1DNaTUiGZ+prTtK8ZIM
oUanEolinotj3mXO57RPJKiZ+B8c1fl9a0aEemiTGl7hTCIsiFxJQxEWEVCbosAn/iT1b7f9qJYw
Mt/gGM6yQWDMd5/Wmu3UGxdWDwgjI2xJlzk8xmKjqMOPlJ9oMRWn7Fu7OPjQ5i2pvSwnArfuP7ZO
br72oKcIkgB1jeiX3qlKA/d6W2YfUtWb8EednGGbAynxSJABDo0wmcivOdDYLT39QMVoGvcnb1Fo
faxduEJ6BIbt10Y9PzBZq/YtRIm0VLW2NGz4r0yDNiCGTcPaiemFcuLeHIkcLzz6Tq2FmxXfDAY9
mnLYN5yvrMqLQXjkkaJd4a6JW5bWs6HaSky7SLJlHihrIIlftdfy0aJLUucm1xgDAeM5FPAcFvw2
pNdHSJ5Wxo+a02M2Ho8OUXOFMlyvm5t8D+1BmRb3viCnJEDQQj+f58trIBNDGClTapcJGCBoZn72
re1uFb7aiFVGSsVVWcudCuQECsHGGww7QfrP6TGou5YBtx5cBDLg5BEgp4B3bFD5AISfSt5JM4TG
9ZbeG0vttt1yTX3/rw8lp3LLaRtBG7DvK6aJ6m+9LjAhIR53IMGgKlxyBv3pjqaaxUD91FDM8xdK
gTTVMKXC/YlLqO8Vv1t6E5gnwOSmjwSl2qyYMGd8J2/n4yRRRwgBYnECUw1Kglx2GSFWyev12KwS
TgqsRpwZSLJ2H708hlYbj9FeaOSpqm0AOS5t29pvmZJSIR9F3XxMtY+5a8cz1Lf/DFOWwG/NG869
VA1d1krs5P1kpyoEWvQbws5vX+5GvBgS4UG1s/enslJ7afvuPNTzO+VM5Qicm8jfybXdzHgf8Ivm
LutklezqGnakoXSJ7NJcuBgYr7aBt0+DK0i8nKnc6RuzmhXfTMuxF2O1vSo90fSd2gEOeEXIWBLb
5oYG2luAxmw1olKZ6/N7qjEmt8SEpM5hd1KI6/n7qWo0oKgMA8SU/MuMb65st7aLwDEYupUQa48h
loD9g10w8S5QOWknmrQwuCwHpb8SWJE2HmDjes6+x1P2D18YtVW6QV/9iz0uwy6AINornlPhbnYC
0eEsnW6vJGcHPSBu8P2ETPXJtpHg+tIqELvvNzPZLTK3xiPa9HHAGoINF4kyqdkvnzHQOKyMPo4X
UAb9RhOKIumBPl2kBrnu+SORGZeLWpf+CR6OYn7yEhvoHZ5Dp8+haSdvPYd3D0dNIrQuGW483o8U
Vq+xxT0zmxi/JdlETBqceM/sppCVdwwVC2DVVZfBo/GjdfFn4ZBqr1vcHr60csqJdBkeMsKI9zSS
bNCw4C97Ry4Ypykz0fI4Q35bT98lQ5ewNmtsfWmDR7D7AJIfQQZjG/Teo7tt+bglj9WRuzFqSfO5
NjB8i7tLa9IJmy1D8Rf1hICb4v60rzcsjH50BO38I6tdNwxuPYjnayFBV9iW2oPhktwBIrNBnQ07
xjsPdRyJswE3fiaOHwF5BIFViEbFn+QQfjOq0YzDUx06FTPUhearU5qoVTQzkD8h17lgBOw41yD8
O5fsYL0xV6AQDAidtUxRRunnPqzvlfekhdFqGx4SNjX8GBkeM/wiUonH3/rRBeYUeoF4QepTcX0n
ZqGOwV947LmkjzgJxX32ceg3KcifGUsv8H+NAFEFDUzhjQNuzTNKZuEvfMv4eRIB0r1IyBdBItCi
bOsQyJAqyKNaeacQ0PmE6+mLX+fCermsWAFs+8/HjrOSVNOjaA0N35LY31Tv7sBuTlBPDLj1xUkE
hQ1L3Nh0zcyzO497tU/aMY52xroSmMp8TAjGaaKvSGMSC5gUmNpBq4hi2x1QlCs+t2iyGCt/+cF2
8hMwdU4K/pKtJl1RLtN+7bZaMRxZvgJcyM0KJQTdlaTSvJc7Fgl+NZ0yuhnKydh98Ae1TTj6jAh+
sdQLKhdEa86zZf37IH5BOqKKSH40pVUyv0900MFjXsp9TrhWweezgaA1iTh4SQj1/FrtJ0y3Hidh
EIlnv8jHsYzN2G+M7gOERd40RItrjO2rhBnaZP+csfU5RUBhUvXyk3sDEVFlW8/5A51qLLQ9NiMo
UBWBl0UkSGH877y6TKBdG9RcSNfU5Pv82URjy1uOwZeUUqK5CYBoa+7MO5aKtSX3cZetELZPBLgs
x8C9nTcZPzykYia28PtIvfNPvMrbGeq9IlJC4/2eBx8z1+U/V6iTDvIwtpimno7X0V4RxmqtNWJ7
mBPfy7b6RjIzmxOPOLweE1ovspJOzbKXBQjvWz1WRxTzWN3TemL7PQrW+s8ijdeyHwI1/dFSkf3Z
hWurIbRR9qzi+3JEyQ4orDGY9UXgRePr1OAaO4bTixxwkkV3xj3r+njjMn9V9TjolRNnrGNJwFKr
k2BH/nYgNLhz8W/lVijt/IHYnP2HQzVVw+DcBEjeUL4SnfW9RiciB7fM/KSbiWEdm7F20ltHllCu
7WzcL2ScHVG0cdNSvOyi7l36pRA7LXKTkPzXfTrMs3gB8qtNkCd4eP7RUAGfeDe0Cxo5BuODfuXs
rr8UGY8Hd09le2+T3z1GaOm5y9IHDbFgX5562rUNeatR41Lz1XwU7FSYdgjKCuYP2yUK9zBtnKtx
GteHL2N3AOtkk+VZwk3VF7DBoRn9WsUygl5dPk8y4IOUqHXzpcKvfd7TNfa2qrMfTvkJRZpdH1Ak
vFscp9DfD2eP76Roysehc5xduX3glTpbp0JGZp2WQahaVAP71WQKV3x10RuCPSobwHS+CJsliGnv
gN0ldeKU/NLx4Uzjfv14b7qV25p0ilMzxwg1lB6m7KL1uH4qsGxSsWWLKlIVef7rBoU0O74X5U8z
Ogjz1dTlM1DL6TZyxbRkujXTz5j/ZOk1EzH1jYEA3GXf54UcaRGCIJGJXp5wJv1uegX69SKWKbUb
pYXq+zRWXFa/U/mRWSrYK3gFccN906pQ4anls7LvhyPH3Ol9RvG0dZQGprgZekQmDhSCaH+6XNty
ktBSVtZ4QZyaEA1021i3fw9LbExUJjzf1/5Ccsh/5ZXx+O+0jsVg6T2/Sxoo8eaVMGF8/Fir2Eh3
NDfyifm/ff7XZuricpgryjCd4loIxkhsyvqML+WcvIyyYxYdC3A3WeCOEVyt2yDLiZ84ZbCO0Z2O
l0Kce1s/vSzn7IlwgcSa3BzHQn/oO8PDn/5lw1qNAoNmmzjGl84GjMEpjWKWlXoO0W6G8VxC3lbZ
SW7L50tkMa0csSgwUV6VlI7xabQ9ZEj3x3/A0+4Bp3K9JC0qvAlRGSIL5bt5qY2ikcwokvgXZFcm
RA7D1Z1lYp4OO0e8u3SRCJ9VTAXav+9Cs1jvEk39tS7bDphorQ6iLcHv3/cHpjZebkGWwF9KmPXX
BAzLzmkdEOxUVYe/5WgM9MZlKoHS53d7Iy7/rMYC0wC3dOI/Wo5H0BmlmjZ5O6dKLZ9YbSCB5UE/
0EkkJYz1tOozyXZmDY5922kvQldnvb+xeswjIc/Ivj1ZBUHGa3y6zngb+juDl1QwZsKWkXdcAcAF
aeyHwpGrjNDMPlC5diwGq1A4uEmh+lqtMJ1I09NrJuR6tvGEF2IR8IfimqQqFbG/CLdTD+2CG46Y
BMiS5LMAdQmK/1vwVrysWCOa5HHNZ7XWxYfGh/kSgoqstcL4rj1oi/iyVXGDTyqYuHS2vdqeK1cS
eLqdjzB50eSAVzmkHXImHm6YpSRflYmnuSgSyGpT0BddG/pcaVKsLzhWHU3dgp+HZhCXHcw6+Wo1
D0s3lEz3hn1EvZ/xa1cIi8Odbnb8V32DGAHb8IvFr+efmriS6j++O9XpHKEa8Huu+iwj5ExtQczy
Gx8eyneMVFYWf13XYkZotVGfdUniFfKYQK3c6X2s1HApe+eukpsiwdHyg6I7lhx7Ey1SkTVx8979
/T+s5yPzMP1gTyV5wODU0WBIxt/pfav5efGsxLjREg6czF7hk04LCmKqHWcyHqfE8vZ/LHDkWCn0
V8d0XPaVl4PXW606DaReKUpwN7A1WBHdl9tdibrx8rVKe+Z+4sDLYdUfr96JdB5VdQOmQNT6EZ5i
tGJ5hMxS3xPyZbYWM7Tpu1G1qUciqXNTDmEorrTrjxaI7GMoCBGifaqiDCgEMzvG5JWWa3rc13fU
9ADCrhwyIf0DZms6sbIYiobBXUtNqmpjOaoN0MMRJ17m2RaAwVcjMTWlSCqNI8XM5QFeZ5cdpClm
Cco9M9rtodANyEc9PwW4U9fp+4LZ00YmhrkGl6gMLFRxztaJTgwmkxSP3lB5FH3g/phDH/QK0jOy
O3JfEn9yvQDLwfe0uv8Urjj1ybsu6SxAQOxiEkbTR6oDCq0Sd2yMtxY9WEKhQpqk0kcgzcHBs9jT
sTJpxne19DQO6H5kOP3N2Zy+HS6FnyvB+iQ/gFDta9v9EKLF+pe5yu6PDOF/rcqSW/PQCs51RVCl
3dAs2hqRtn52RzyergqHwGCmrWL3Cu+NOhiucC92AP+PRF6e2xNxXH/QaIEzbhbpS20V6hr72JlC
QpvNBpdVPUqLsaih4pFHxL8rPXcqJGfmEQeAElMe2dlWNcUXe+VOKUrqjMbc3ubucl6VoRtSiq+9
6BseMabflFos0+dzZHddq/IhY2DbgBMVJLare54xj1z9bl4NAPSVJOr7hBb0ofW8kHZbMTtZCvw0
FI7hKTTzP5eFpCFQsonhPMK6zh5zceyRijDn/686q2ehZxpCxOqAyBDMk+mKF6Um99pQ5AwQP0m9
C9jCCQHgmCTCA6NdltwSsxikTKRT/PYV383IqXuYhRtKpKUqk9qYsRSK5+oN1eEo/qrRsBeUbNU3
HOJ2A5p5G4msoOmTam47lGRR/CKPSZXeBU7vKSy9qLc4vcDhfkEA3fDW5GJ6A4bYI3fNkmUW6OXk
Tfanj9xaXJQ5XzAAY4SZRiELo91eCXwgdXjWAzlkUreyKd5qk81mVk97mmRpuQ/FcmGOtGzLy42m
+6WU54lq1JmPxeA+2d2B3EWjvaMcjgchBosvM+wwsRNapDvjSfVIfoiKtKINwNGpnMX+CmdyhY5F
0pVokpCk2OHxWooenX5eqQBsmOHCHLylNcu5/14N56dPo7wn1qwyHIY9bdAttRwk3R9pXJcklVfK
CgT9ZZuQU7OOdMCOsi32BvWw/pDiqi8oJgSrw/4l1O1+gFP0Nt/cx1YqH4HzNW6Xnf8//P0eWVg+
ZWdW2MuIUSUQBXqURnISh0nkPsih9eswd+jw6CTi1ob6lg9sMZBIJOufXvyceSUBwmu0Y12aQK8c
Yct6hU+G9J0hor20oFJrR7eXEYwamC+JCrXA6ntOmLmb1NmltuRp7SORY3NGygED+HhmP9Se6AFn
T45ifrqOoe5k6CR3fvGs1mpgpQAjg5iHNAq1s2MJeNpUpqvciWEoVXQBXBa9MBIrb7grdw73Yqin
J6RoLsUpoJvXOe10ZRGOC9krF8LiMc28M0NcZAA7VRqZMf9upaCjy+4+X+PNY66o/JKTZuTFGrY0
bILYg6OwcPJFJbgG6KDmLk03G2abDcF+yrXL0VflfR4fZdLP7GfwpoedkJqbiXx1e3cN23heoFJ1
zmg1zrOsxgC+Jxu4gVDJhphQjfGkijlOreja/6MgJs2qcolgl/J774lBe502dRUWyT4alR8jIpti
65gSW9r3I3Rst62VbwULbu4LDEmmE2VbbZob0i4PbXfrqB/kiuciK6MYEARAsbnd5RK6st1sy3Qv
JRHVSOuf+FWjdMjs+XMpqP353eceZ3UVpTDidfORrPkrHZqndg5K4C/brKPzx4VLu9Mn7Y0Eawd1
IAozBMbEUKAPob3zG9/71fBBfvCabFYfneB+auumtKCnDGIxX2rlTZnrsm7T7yIzUH51zCs8EdxI
NTLGfjfQw5vh6+BSb7+p/r2MXF8NiyhpwB5yODRtr0eNL++p5+dXEuMAaOM64pJpIYTe9VNx/fct
jjpqxh4Gss+VCYAPPcJvzRISNY/HvUF0tuZ6M1jtRPlcrAu2UmGjPyGwnP+hG212tqTUUijYwFQV
w0EKl55qKSXUz0BcKFdsjiKg/WlLxXQOz/fP67tk2R9aIvd7m4hsR52aKrZZqugbwZxUC2IuEzZ3
4y+KDh0JbL3fJE10VqjOFE8jP0q+QktHg3J9KFdn61uCDAFny62qH7D0G9joKEpRDw0Wcd/E58TX
DDlc9tDruBjd75Bq1hcn24HKFWRPvpy486pOUFc9Yl3ctdfqwC/kCKUZdjrgGdAN370/tklrF0Tt
QKw5jWVSZn5B4Drbi1pKH0YQbZzSNnDZw4P7lfHZ0tw/+9iEdjIbLc4322U8jNsUj2f2v+gKrJ58
+tNdHrNUYux5Itn1cKgkq7x6pzlq3iOdxrx7OUK4O9fhA9mqZEslGcIBAd1T8BFKR+scJqqbbfxS
2aDdnlgRAJr1aOSkFURnmJEMomX3qQOIyzxhd5oMHf+s3GqoYCVFipWOBE9k95/kCOwr5x+gj+dJ
9R4AOjY4bNJhmibcKOAnOo8aQ/1uOGfY5++1KC6Jd5oro4WQ2qmayqRkV6XI86snru1IvQzk2hA+
AuOVGPseW6vYv6nW3+9AgHLtTCArayjNBjalr8v0qW8l89aAkO8anj8j5K8e4tIiV3a0ToEEnL30
GKXuTWKvvC8T5dslJjqzljI17veEFvBoFSfzhxN6mOqTn77ra13h/Csk7x5A3WpfiZNnd3wLKsML
Qm3UrVkABdOZCw05lwyj0Jb6ll//AqN+H6mf9m+r6W42UaeG8JuFzL0WtUHMnhRF1vMgD1emFHa/
vE888D6UMcLcAiUlPdoHSxjswT55yVoiq+EvjTiW0tKGGTD09ou+r0jbKqR6gXRjWmhh1tJ36mzR
aDLRKBe6c87UkAREq05TfgjyatxMI+bb3xQEzR+LVfgCR8qvADMLyRMPsaqlUdGJoZuj7DYaYOKq
WEofYuq7oOPSvhcWF2hnoY+q7qPBqsLw+39ZzIk3H1Yjc7Y2AC5iDFK6U0SURucxhB7yXnGJLB7F
1PzqF5MOzIBHSZIOzCwEYFQyoR+sotuHI+hTBrRwpayMCPYTyg3on5GZcy2XASv1h2wehmAU1Y2b
bOT5u1sHi/x5e/Zi8OxTd+hJ4YxRNsnlDu1BRul5+N1AnW7dfO0DjE2VHgVXLVd9897fK3lz1evM
HuFBpDFIU3zkbXE/c/muIjqZNiWsHt2Z3n4VukdfyrfhPpvS6DRxi4gxU6YOia98JM5vr53UF2/c
/7iOzZLToDGYQRsGwXg+HjkFIq/c7Pl/G5rCYT54hxZ49EQh1Ayt8emLZ+v2zYIrk3/0kSZnE7ju
nMPVa97ZBrHREQ5hYVH0XDCHYL+aDdqqwqU6os8qH6OIaKlC6s0LpwccgCJtbP9WXvYwyHrBfZEX
1HOB6WKdKjuQ1sw7EhiFVjnxxLVs60GCzFmOVPGxcrwa7u3hwQmxLY4XW0uc4PdFG+Ie2/OiX+UB
sBc0hG1/MyuWnxEf+3JiDG4IGINF/wIZ2XlFIog3FigK+OkVf+6RYVbpHbg2XNHdjfhX6SHhW/wc
iqqqnxRRykV5QjME6ryhFcbtg4VrJYb/NHFUnY0O5erjocdW7B5AdUo8UdTPiFXgqGeCkAKkTyjO
sF/qmIwvTz/HCT3kcvd1BUmcTCKi7GaWrhKdQIgdVeoDjVFJH43nxVbSz0aaoswu7dwc2zn9Uvz4
XCVT5sMpVVsMHLP74nvpa+SiogDTCFmK5SoEnsZbEpAU9KYke1s0rt3AaSWAKJsv+w5ngMP+AOR5
U/Q2mo/K8X4v9XYDvp7BCvYBa9KU2OtWvcHqGhjJbOOTpJ+F8rbuw6TIGkRokofyZ7HoH3Erhz6E
Eyaq9mdwM/lVgBZOG4WffdfAvqEPPS4R5WZYo5FJh7a+5UF2Tu4VDJGpYIz2LWis5fH/cIf3/MXV
KkPXx8YyTwnna/PQ1AYgYUyA8mPk1H5q8PADAM2GtAaaUKSThWHg0K+vGmBdftmAyWaYKchzq9wA
H6taZ7VUNSbGsdteDds4Lr+Ha3uqMgiqt0mA9eVXtGSWXgEOOYzdgQdogi5CZa+RPNIDwtg2lmKA
kRYkFSBeVymv+yj2xkabkx9UCJTJRO9XhGgV1aWbDg75BivLOFCOS7erY5jUH1g90gJJYqcc+eJy
Bx4OPwgYJweIuf7lXEczKASnPZs4Kkr8REv3VpoKz+//6VN24udehT8kZGwRhqAZK7aXdStMH92C
Q9gZ7YbRiSOsdlfillJ3xLQhiW2XdEUDqdD9nYOMbkq+9ViUrPd804gKu/G4A2dUqbRN/2OwwJri
LuE7EmLAEIJI024GnhrrW6PGBbM4U765jCrJYSJVDch7yF40M3ovldLOARRhXz8BvMBFPyzXATyc
XFos0yIjGubVv6gHwCJjli+DOu5Kz+7LRmDFHSReKk1ZG5X06YM9bhsA83dd/lkKxKsjtsteqEJH
2i7c1V69WwNdiFzWLiRlNPU7YUih5cE1lMJmZdKt76mR/r2MQqyOhmdfCsJOqjMm6IfDtcrXG3SH
sB2xd/i2QcBOYQGnrdCODdTtKFIUTCTv1NRYEN6rl4Pjxzmok74ny3T+ozRD6cd38c9FQkrPCl7N
Q173gpSXikI1SZJIIM6LfLopz9efpzpYsgB7McDmWw88hw3OS1sQaIDzWg+cfsfk09OanNyR0R4u
xhjXCANWtboc+QAo6Zp66nbAnPCohiSnn09P9g/i1XsGOHJ+mnL68c3nm/PqYTeENGJfzxDUMj1X
1d+EoKtve6F6Z9ZSy6gAKFTyebj0SvOr30O9Hw6HjdO6bYe5ir5yVhIkl+vYzP0MZ0gAmWZBuSFB
K9pNdyRjXn88gwcFBcUp3M45imQYif3kXWq+IkLZEqKcnrVaJLCn9qT/ZPa+edjj3bAqhrFi/Jar
nrtkA53EyLmNQymLzNFvRjo8vNzS6dwZ9puq//jlABPPx04YH2VQJJ6pwisxUUD/I9qNHy/2/v6V
vR+ZTWuvymYoVkCbyfAqha7qmyyndqm+Yaew2QlSrS9QSkfWvXFHqVmiuf80z7v+BEn1oZFBjEBE
m8BVOGAQbGZ71DlYbCZ8czA/LsAnzzJj1sF512U9/vyrbjeUrgC+Im0+Kbci9CXpOONfiWLivYzl
CN+5jE4xuR/DTr2mVD6VL5LhpJxJ2DXb/osyb2N/4RGIcIAIHzva+y7eFxlBLihtkdoVQeYSD24c
nlV7XuJJ4pAuun8I2CDEWYcnLWX988Qxj+kg4sYd5Gs5nECNJ0RTEKa8gKgC/Cxge1Z80qrr4xid
BILHiHr68JfIrq4u/oC+HoSKd3LeRvARGL7+P+2unFqZT4e9tmIaQYg0zql7ciuylFrubowUy3BN
LpUYeKXWVluOmZk8NYhJW3tmCSooivIsj5QIujG8ZoSghAxhKs42GnZsUqc66hf4ZyUPOEfXtb3V
kXoeAeQ8Vhn9dXXT0RutP585A5qDbri5JxkFBWX/AkyWP8qTNfFIyi/sfv53JUsSuzS5oTUbmnKy
e74UIXcWvj2Co3w7wsequVYpv77zQGWNxTvqXbtth4+mwoCMyiLL5ekZAe3MB/qzS9USSoAL9HlE
yfAPkzPR7f++FsG0oOoG9tSSU5r1dN+tVfudacJX1pwEVzl4zVpvHaJVKTO0O2w0NW/qd9opYVX4
PShsxUyN99Nqi/uH6z9aqWHUybf4NRl9gAA/Xr7tIMD87T+xruz5/Xeh28+Wv7paspqCbGME72mp
5YPclJrMFmHBEIZZ/KJlNXEfmcySqhNZBB6hIVqnuQ7+acCi+AKsqf8h4HM122vwr55eoSVA6PbX
hTAJrt9k1i2Gnqgu+4ylR5IqBfS4Gk0U/dtxPBF2nN9IseejEURRbkzsvF8yw7xLEKFAcp864LjE
+XgIy2M3V4IOKkpzD2/FjuLoE3W4WZDrVmOqN8scAnmJgUPQoUQOJMVxioA5FD2hJzWR6etCITK1
rXYxr4++2l2CwgDQqtqWqL8KI7o3W8cE72FQtowz9VI7nXrGqw04QsYANyZKtuxcDgW36EZS+t59
UgZ4DN4M3Xfk28G++r9qvjlZwNRcT0OIjRpV+HKW1UA4aW7lE2LLK9UcuhMc6iPO8zNkrxEMWu9Y
d/7w9DX2evWO+YokL+/C+IhVIa5LddoNdCrFVPgiNi2eM5ZYredmAim/H8Z0GGKlC2CNz/71W6a6
rEW9BVTCPWiqBjHFofb/dZ5AptznyWUvylJPuxLGCfD+yEOG59lJm8fI65usXnLZXg+omdp3g1xk
adKqb5fFiLIQgw7xCOwbvMI7pm4/PH8OExGLLzOSZj2ug82oboMWhbkJjSt7y7BbvMyPvodmaRti
TZE1mRppJkdSqa2ZkEvW5fZZP79r2W0RiynhY4FEjLgJweB8GyCPjCSc3w4BMWGwJuKAg2KTr6k+
j3XdrjLbhJMXNL2aCc2wBcwUO7dq7T9vK75Dx07QRuFm6fnm2B6mPgACkiiUSBTBWVd13wELNgOp
ShDi0FTIXRUpcXaKnKvgc+/YY61NynskpAGVw2r2eFn7qC3gjcBbBoe7oqD9vATyF4u81c+80qa7
GBr38+c8mWyHfptr1xcKIAUoWsTYx9NmPlPNiD9N70nk0MTaOM9Wp4Ox6u9yhSevScQXPPceqf16
JKagXZGmPy+tJcA66gxGUO2iPeJBi74jrdN5tjt2Y5U5PVz/xwI79USeC8ix7C9tCM8il5Skf9B5
gve7Jeqy7E3DXjSSKBaoOBSKU1b+KNTYlKzr7zDjSBF+LGNp71ZN1iOWKNMRIbuiLtOgRaj2nYy9
pbuena1B/QWa242KH8VsL/66f10e7EMUkbhkSC7SyWtQd+rbttRCtNhk+d/9mFCGhFCNRANYaL2b
lnnanyKD63wRD9KXgKxXljaU5PMClQaDkDZdQsHFXlKFDtreDVPxRemIDG6UYO37GQ7y+IqsUuru
gO+SOhXTwSRN3MA03V9zbBVvKx9rXtOk/KpSyL3bJ+nRIXEUuzWsdIA64xjfulLm4TXDTbSP0Wi9
RFat4lLe5YYNSKBUhh65WzCFeFhZNJ/5lqGeLJAJdFuAbseXqcrN/fgYReHn1RNxX/Txtyho31ab
3md4TjfV/UroISwYZTiWo5eHdrVm6TLfwmyCa2mnjpKMHaeNN1hcxzyqWT6Hc/YwGuTwauAB0i5n
RknVNFcHdky9yJjpRbwVepe2ZeeqymKhNmVGn+6RmkLTcSlZVILuF3dsJ3DPPkfA/fkkqtmz7GrP
7kJ8rDQQv3wxvL12wX5nj0N+JIDBy2yFSuQPB95F2QgHEaAk6hPHmFY+ZvVws35he7yJFmepvl8V
Lj2RWDYL5DJrrbKyhAmbwrm2acIVelcydcLoZtRI9hGn9o4f7RcSLqlTwbkIRJxN4fv+peyi3I71
W3BJHChJ9DxgKHPIaTZqvIoTU/tlapeO7yLI8Vk1WyHPQ927ShdXxUkLFKYq1KyMXRcH1XJrMSoX
ekETyJ+CVEpsju79Xh5gOPWUKEyRPI2gLLf1ec+xAoKBmjEq6Dnzk93mzeW2G2J1jWoUv6U4+loz
SUBDMpWVj3k6g6HGQfZfM4dbJcnt5/zdPdO6GvmRnRc+52w9iCNhjFazUnd32Sd+0xXbkegkOLE9
i1ShNs9vrCejG+D07yheaNnL7Mue/FkIkOKGH/3tZzFGI46N2cMUDt8aQJ4c7J7ZTOEd8fMTWSqD
a0zuGMbBug+OgGG7MOxUsd1yhZSB8RdA1GVz4smZdow7nrU1c0a2iF7YBClKMPb3EEIiDXtMbC2p
j4WDeOz3ekczpqab1tSHuZkLbMO/nI1eltCCGjt1aTQVutidLUN3oIAOAmAUlUUGJwBJz8BqZ4Ac
4smkcikCrkMi5NY/0GoS+0/vpV6ZRbU1T1ZdQ9nuG1h7NAxALdw4VocOt4qdRlbDFOg2fcOUt9Dn
PlHk/GzPAn7wcze04OOhva8xOHoY+qIxzYRYG27yzF75WQRJ7MjW6duD06gWVYsVpZcZkBFYS/rO
8S7jf9SNnMZKumYaALW52aV+V9n7h8ceOxAx/wm0DzvjMz2tPw2+8qZGLrKNRuX0iFgDIwhbS7+5
zuVUVL+oguOgpv98YNZDSCPrnjdwqbgef++MPcY/dy7UaIJ5qgUu6aavJhAb3e0nIwhSk8WlUJqV
34iP3jb/c5Vp7mnvAZMPwdjMJvGKsIQ4wbpD2nEr/tA1ukFcZupeScEu/1I23EBOeKg+JIDfCJZ3
odc+DaEFgr3+I+hPuIOcimdmo14ICypu3VDXj5pSteCN7O3shSY0IYp6YMznZ5E29eN/Sj28VxFG
mHYyLZp9FWg+30rM1reOG0wml+wmR1quc7qV4YCIzodanir2atBn8Dih7qs7IyxLqpzsN85ZN2g2
v91UWZJ9Jd2K506bF/Yqw2C06GFKQfIKx5+U649ziAalFhw3yfvrE16r5Lnn2nK5A+VRiahq8ufF
a9nDEkygsDYnH+qeT+2RJogNhF7ANGT1uqYLX9vhljX4YvleRQdNjqhOGul+alKR6FJ+QIPZl2uO
8cPGIcRD7PIVbAFfbth7DVapclefxSWsI1v/mrAaySXqcbnK3MVfuFFEbuEi0TnwFUfO6NhL9Htr
6wp7CyAZu/7hvhdP0UDV632F1jJQJoErvnnMC3ud/OTAwBqLxYy6d4mYyPtLpE1oU0QGn+wgHMYX
A5lSH/SABJYEwXHQwpLDySkXZ/3gzIzdxpzF9atPXuS2SWH/yc6aLWZWknhJYyraPTS/uYXyF8fw
NLGvWPooM2gnrwobvvK67aA3BQkvlHheNSpdTA1syh1BJ0ysHVTX7610MyjGgOouIr69mrqzXTci
OmAWvN78yniW0I2Cpej6QwqYHJB3xdZBHROzHMN/8PdAN5KMskVHiCC9bFboa/zK2v7vJBpkNXji
mU2CS3kmmBHBFFp5j5MJk79xteBwRv8rfF2E3s2KDBjs1IWc8zu1SwFKsTCBQ7avywgypUCp1RwO
sLf4Af7rq8mMCyQb0x0sH+4K/CwaRW+UnRluzWYWIK9UjTvK8yJSR7jJC9J8IzqZiD/T9s5Aa9SO
JSUC9mWCqQ6dJMbMmAocTQCCQl5V8KYSdfM36mfirLF1wXc0UtcgTFal0JTI/TL8b3C9ZfZzWVsr
JuTjXALvReaBlqn9YO1UtU01GCoa/jcPDKLqJIpJVv05J77AgQN+0i7QaUOUX9x0k+cOaZcQBOVF
TneaRDy7LBneOxOntmYvqrSfbL5qBhfLfU7rw2GP9PRUUIAxrwxdrqdViK9M2btX5mhuqRD51D/N
M3tISyXnnlbMRol6o73uUgeQG+LjxqLnKVV3l9isx2u9Z0sY2VeL1/dB4xhQyy1RkjF7mPTKKOAT
462kmUGkcf5bis760vybIGQkFhcgYs6GdNsSC+Wtji9H+uhYdXsm2j9V2pACu3WD73ZCmhyRkIyw
RGUVofbXkWvnj1VgcDtpxT+o2FehnmVi0FGDxh1+tHx+RFqts19tnewPOfIXmRpc+6q9h6yhvLKx
0UTZnf44x3XkHGq10aDO9UsXs47a4xkh07jLZpyF9ACGHVTKqEgHuWO808v1v5OF2Vuaf7ylcSyQ
xZQC2omZAJbO4jJhuWFnKOn/Tyq4iV62N0LdupK1b7mpt2Ed2/anomgNtQnf5SeifdiFmJRSuNnF
02thpbfVrHf2Pi3KoiIg0mpgaYQCVJUaQQQuyZzCIshrmef+jIvT15uXhUphUGuPZb1F8nsDJq5J
N/F9gh+nl1FsnGO9T4RPN3XNWdQu9YyT9jrd4CARu+2aeDA8fX9ioKPTYUY7asew0MIE4dBEQ7RE
cjJIiYcD3o3Ui15QR/ghiTceodbH8AyhJBXtuhIdXYW/j3M9LUt8WLoBDXGhJf2zQtFdQj2a6OC4
SymDjlEdop5qd6zRXpC0K/C6Hw3LKlPGbyIOrYkOfSKw2U4j7K4obcWJH7fmOuI4PhF0SGAJ0HnM
Z7o0GqNg9tqftV9OzdW2hca2TWzYOhoCiwbn/RmNzOuvUvHwMV33xjlZ2KWwICh4jzk4PCD8UWx3
1YugFYNjGvXB4yhMmY45Fo50LvtFCq9I1fGrXrXDgKd6esWZxPssIvS3Jsw9j0K4G28T/xNpfOxb
+Ry3Sfnx+sZQarqPjOu7bbtKhRm2vZchcDuzI8rgXECaVokOSBNWWM8cEGVnmzF21ZjMA/PTWvSj
dEHKLjAawQ0mI23eO+d1LNCUeNLvZaWWF2rSE0w809M0w+dpaLpR5MxK0+1/rr9etYL/QaHdNAzg
iB7N8yzLyZ8KKYWiz4Qw2Ez3taDSWsbtUakCpeeMHCffsqRUAYqrw3TAv+YwZ4Y8nCoYErOTFhpo
j14QC7OWcJklWNX4mXxURFHLMLauFCYTD6CdTDSs6vXm6dq+cglqd7wIpo9gswZsRnGaiVFM02/p
rfvCRhjo+kg8rvMC2OCCQrOfds93YbUCLqsEf7G0anTrY6wmdllpkP7HV0AZ4hrfy8102GdO491K
+tvvDi/cNFtL2diG36u5NfHcXTKpH7tmOMzEUo+tJwCqdzUxaDn00kSoqAIXf0A6L3shsyh7rnA0
zoSoRtqhRXE19hUER6cKGxW5B9mnmTKNOIheAvX+SEY1jQDWQaMKCG49ir5TW3Q+7Q0ioWWMAAw9
MVYzNuuJlF6543hsN0dRro+NHyf3K6JuRbWSNrwa40lkvGnoWrAKnY4qMZgONt4yKtS9VXSgD1e/
mqmuPWOLs9cJ8Jyj29FuGmsms62vx68uFS4KfYALCjCgXjr8kjhigWOuVfmhjuzDH1VwgEkWYd6K
7U83v5STQj7u3eW9Fs0QcuRYyZbz216lnIZOXZLzr7qp/JxKWtzyUkhT6VbIGWoyvTKnBkKPGKe4
jmHdadzcvk5iuSm+DCDJnJszP8ijzZmzSV5ys4yLf8dHUSfQfvW0poMozyehCXUetBQv9krR3LvO
XtSpAXsAOdiXpcGOlVLSJp5OxMwXqE7RnzeJuxfwcZadNs8p/koB8gm18HKitadLAdFB0fo+A/ly
cO1xOIQ/a1AJHN3nr/xSTvcEQe2HOEWiS5bu8T18fnyQ6LHA/MZxYFsAY1wlTfPas59r4G6I62FK
DHNOy5ZhFKowSeCVGJ9fuvzbSW0gxZTqBlc+MzKD+upqNmJEp5MmHc56VLc8aV21IjFII+Nlc7hr
VLEBDxs/tZvF41uOzKp88tojieHjPdzYdK371WFk1INa/18nkzVULUn8uH2bgbCQ88SD09y4jHUL
/ARwePEUstATxw/VlhHbukxchZlUXJN6ibxM3rysbPkS8BMF4WGBuZOyAgIxJi29yIau/gdUoQin
M/jzcEuHMg8oiZZS3BZw/L9FObxr6o0fvlvr4OFVax8v3WJs+47ijfQS7+5BGOaSpufHU7M/G4Z9
1BSZNLwur0HfeZ9vIKboQwqqq7KIthoMI92F8cksbQspM6vJZ0N4/gARWbhlceN1JCENUt0QhVmX
zVJLshpVyDUSEVfpinDYMyER4YklL0bRgG2HsNCJnyv0NqhbzzPOPmSNxYUsxEYuediZ8Xv1sOfh
mrim2Sfa1xx1c8RUheqx91nG2TKtm1UNP/K9IhAAUl2W1rusZY4kw1g0LS36lGpUw5X7jyuLfLRr
HampeOOdfufij/+yEBL5Tzw/NaK3N/fiKSK5oLALkHtrDXeT4XUaXQl/YNaywRr48uQlY97zV7+r
1NZMxZ0xMMrzE5spYSUvwfHvznxkhjtP/DcKAkBYMnCmz1O9k3//PxbvUNRGmQ2zlXkeBKShB6n7
J0z834BL6hkAx/2txSXGBk+cL+nPUQJLcKOUlqZi62kY//TienqycCKOnxLs3H+36kgZM73kiFTm
/izIs4Q7tfGJmFx7ikgKXDUuTrHCiteHVKqAqYs/eJYE5Gox1KCNrWUmFMfte+cbcaqN5yzXjPIy
fjRTJdT8YjNX9CIziUDzsuUD9/U45S+UgYfeii6U4YQN97Hqo6npZ48UxqSEFhQhHfDGum8B5xVC
1iWmWB3B2Ob+sR29f77pPFC6NHBwGp79bTJRDWphMd17UEbsfyKe9X3TlhpZjPKn9ewcmJKFy86X
x+sE//KodXZDmqWV4/73wP4muqd+Q09Q7DzFnErLgGO9kv4eFnzDNXrGOUPelXdAwvn4aTtcgkG2
IFFv/ERtOvF3TOp3ztgaYm7wDqhfD9UiuV3/GNbT/7edQx2liU8LElmSW0ggNnGQ8B7O9CQZ/Mjh
fIrG8rJHNZf1QzLvZEmpLsI2b3WW6yExJfx9Wr19oGDWMdqQSN10u6nv/aAFEbam0VWNXwcvZJLz
Iuulcso6+wptRegehLPRVsEJg34w8334PLGGEf08pHL7OubEDta8HVL1ddGdlHQd5A3itpmVAGNz
YgtZ076m4dR9dzM8BG0553dvjwgrQ8HW3fsavypLxZzrMGawi9zpLSwaSFQzBQR1ud4efZOqiNlA
S4oM0AoFQumkz4KR4Ju3sse7sCV3GiCsQSKuhisqS8vI91MkDXM3c00ZMydsTYYSpPuiX3ddBr0X
UCTRR33SN8TyL5fSamN1t9/lT2kK9lLD7QKNymICBMxpeqnoWiFw4BFpGOfEMc6Q98vosxipv2/L
1H4cmrKxNmUbTdmhG5EGF5n4SmqPOFWsuoHqpE+rp2no8v668ZE3wHC15V0HCndq8VcBYfETzfLh
Tv9exE2eboGO8XLkNsaWmlKrfwz0TIlIwLUxalgR4nFxHpm0WZWGCfgDYQnNZpm6CLuBq9s8w5eq
PxjNA4QD3CLObXbRA7yEnLjwOaWcx0+0zbGSD2BDulLhu8WCbGYo3CR+J3iHSYqWB3c0uAtAy6a4
SaimpCys3sMhNTwZzBA2zB8Jn4pEoP3SquKI5gczhZYR72/iKU6Gj2/gA2WOJ5EtSkOJwVnyZFiQ
uSK8klmV0a/q3hD2YKuOA8wlbAbnQeI0XOCvwXgfZEqd1RTXyNy+FwVhH2+b6kwScNNUEUZpsVLX
sNct/7wXGLYIG5uhNQL68s25tn7N3hcqeRxNVORs0pxKDx2KXtIP0oB9P88uh5kVgPok9NmlnM5M
Tf0DTo9Tzjja0Ax4IUitYfqo99yY2WeHAYqOfJPA3FwRlunwjflmAkAwuHyytE49GmBnQWywXAPh
Z4hrpFfyxIeMOHlIuPyPBcFyo2o6zALu50j1r+y4a7qYO5J90+bJB0NhIzs4/UZzDxtD4n476ddh
0UTHVBxk2LEbOu2xA4yPGdVYSal+jQYXq9I63BPnIBzxd5m98P4/A6UadcTiUzNgQg27sKvd1bU/
T1hY/+tX6XTweR9gGwZmX8iaOn3DzMmCCzX0TKPY28pyj44Hc6dYNMS9zhzSqABnc9uBWrD1dYhA
Vxui0wpzsRg6jvxMQc25rcqQSH47fr2almbMPvhjsLi2GTJ4vSbW1JDJYbrrt2NN/2KWI+Smc/Lb
L7Q4JTYBYpo7a41BW8KdNHFUMqR9eqIguXlr53kLW+RWIOX9Wya7iPzo5FfPpWMmN9r6X/VFicZd
qzRTQv3W0gnzb+DXbSGTKn3fn5nA/nP/GDOJtA9Z5wZcpX/lfZBbl+EBKD+PP70UEBjMoLBYBh6b
jvuetYjtIkOwoyihY/IJVGx2yCa9EoS16WvdvFLVAijmk/a8IZhg0dYnfjz7xMxGctmxYSI3fmta
iICAnggPQWxKiT+AQxldzJlklSvFhRMuBPHYT+jEDtx+vAkitxyOWJGryWTgppYYj3c5OOEmP1T8
rgTgWXmLQC6nhZW28kAOz97AjU3yISzZTBgeR7vbO4jgn4BTkqyZ72JoYJOd9LYSvWO0Y0sm0eKy
OGzuZc2wqZAmqZHoqZ4GkoL081udSCA+FvJY2lxgpwSZngpFVI5XnVbCrBGgHIuhOPG5b6sCNgTn
S8JWjBilgMw1+JMBRvDW1QoOxI9SLxhui/zsH07ltqqlM1/0u3qbe61RoanB9qacxtlzmnKOaPDp
s6xkwKai0GpincbKqy5lK5ppE5s5ews5aCww4/pAaxUKszqJIFSXZA+LhXWS/M7w9cG8GSwaBlIN
RDcwuQQnkx3yHeZU16Cfri4gWCZGqWf9w68+19SD8pB1R28QVloPTMU1XeAI5ew7z3dl12dp+XgM
FNx6fwh4SgRpdNhb9ioGcUr4k4Roe5EyDZ9u/zyEFCM1bzhpCi1qVHyWO0BtyFaH24XPoT/LOljp
s1JZV838r+CCerflhHNUTtqKrbnZBGv9EFCJfw1Sq5Pj2eGVXx9DXPkFx59QwEa1uFs26gwVoYfV
8TowHSqtNTzRJAnU5VZbj9uZBS80J9P7Yo3V8L4bxcQXctjcT3r1V4Lbb9O8RrTPCi6N7cDJXct1
VKE4hJ5+WUVfl6uuM3RA1KI3oFLdPK3s/ZvZkdTxgRv1ZZZ2s3bbNQ7QX95ZsrbnPN1iY58iT4vL
hvRP8faciN+NiWM8XOZqkzYQPRiJtsMaqfQDbbps37GhsFNZ1wJB8wA1r3kEPdPmDh90tKCj/R8u
5qZy41jtEGlwObyt8MSpKkShBY48yoEh3oO7ALytRxFcBbr054QXq+TlB3PF1SB/BBMijST+hKAd
QN8sy9/1oPL1eR4WTihLoLejspV0AodpFwfkz70snvxzSEOJblZ4mJoGgHmXQHXTWdH1IPd8q81G
55n/MVXcNWv8bOkA9xeyK3wR9snEhCI7VDLXCA5Tt8iLr/TuZK5gIvQmQVIq9y5l4epHCF58aM6f
/nu7fzi9p+Eo+8FGTO+JV3fM9/73hupqOvKsI57nOwFCxd/kCw6W9e8TmHizwgBpVl9ru6QWNauZ
AzFyIL1tyl6UhwxozdgE33HGRH0N/UZpeYEtAPKwpeL89UU577VgZJmV62yz6qgpyXWSnAvnTuqT
NG81ehzSTxKSHz9scAfsonEHgcV13jO6W3vTp5KhgPD/H8z454rkXXo9nUQDEmUq79HTgcM3sqXp
+KSDJT+WPTFpR/rnn4g/FhpZAK49aNGILO6LBIRINDXaMkQq1Cv3sA0XRe7PLjrlNoVPEU/tEOV8
oO3BK70h8Tb928FYOdT8yjoB47y0l53e4OGntYTaRaaB9A446JGiqbksSlnQdHxHr32WRywyFCiK
qetErTGlfOTkn2dKd1re/AhrlpsgCzMCta+DV4AKTehPRess9YHxDEASTNG11jxtqwNAS293ElcM
aF5qVb2CogMD93epSPAVDvBXpqABzUwfQkMjBEQ9SNlRd28MI9IfU+ZPHKUqGRcUDxwK4/Ooe5wM
3q1YsNR5Hha3s4e76vgYoovVdB9qJSHrPq0boe69MqZ37fRMch7EEL+56yC1HA0STGfO/WI0hc/C
pbhKkgWSd9P5M2Xu/8AN5ktQnHb8wAxIVQBpZjrxAxenDr/QRHXB/6vq1OhW8MbuQHz5A3YpO4QT
Rxjcn6eiTyscA9fUuVYkyMfNHKVhj06DpSqUMTSCGPKp5V8WKgekvfjgVX6KJsGrtSICt4oeva7H
/nmcgaJW+l1MjXWAV95wNF240/EmRmUvd/aOf7kZ2TqtHpkqPzeY/t1vA5H0cNQ4H8b+QaA8gpqK
DNbqQPh+TvGAaD45PF6+eyunLL3QUH7BOwxlCNWRbyJskq+3KoFAmn+EHPvHLgXQaPFvto4sD02e
lUknuZzBHJJt351xkTRDuCHDAA/bqYFlJq3CPvVPzy4iX+F1OtN4rtaWWndz67tajMWKGxWzfXyg
QTpbc6Y/jUb3MFS8ESl2W0blUn5+nSofRGj4Nq/yaUZAHzO4yByDcK0ZfpoWgjlSXYR+YHP6zAT6
kta77gRE65J1Ybhj3dAWW87+cB7NOqbJ6YKuTUFE6W/J/zaAUScpDwHeRujx9x4voRH2A1biOOyJ
eeiVHN9UqHIf6GaAjdL7AP+G4np2q4D8eQr9Hr+HPiEQFQfdRMWQ/qc4Rpn2PvFWh59arinRjYBB
90vjyQ5i7HO/U3MhQH3zB7oqAYRbsDlsD2CkUU2Klmfg6FDp0TlivDbsSNxD+YLNgWNw7FT3lfYJ
+zu6aWlqL8d2IZEpkxzfPR7MjW4pTvXe13yxWjxqFxpykW+rtUwlAjr32x7v0ChsT7eEnaOD4Key
snUheXOknwyzn46775yPjH6sRBVn3bMEjGFpe9ykj5n327sfiD3WQpbo2Mr+1J+MhyuOUujTwNOX
5uyU9BLlc6r8jjIVku5ExnURIZVJur4063vAu0VEeWV+zeMXC+tbXJV2PT8KI06mf/d+rVZHQm44
Ks2qVtMaPStTUw/45VA+1rLKIh7XkUDmgy69n29MRXu1IXhJVHF7YFKoI2rwMJEF/V0yA94tzbeV
fA3K/t9no9SpRyObAjcD+GOvI6zC+X13zgW4mb0dB8I1WcGLKmnI+nVdqHtN5UKkPMG+s2ILkVMW
yHN3rGi6YXrd6zNdckuoXSdnI4UXlOqMQC3TkVfuiJl1ipyzziH3/RdZBXjBXTW0uTOC8EUYt6NM
5mMK4mzMDrkcxpNJmIAWv1nzhfkTDeNINwTLQhG/Vxqodq4i6qZjU2kbg4Q40Q8clMOzCxEJpa6b
DCGIAbpMB0GGePtfCclLtpQUtgZZyJG8+48GBLhSrT85CZPJX31+sPfNtJ6FMXasuLU8WGfz9jxI
4TfWxyGhDB8PSsoWZYnC2eX+CRQtMvomc/K3eU59Mg0zvOGPSayPMy7eUxZsY6HNAgTGmd3xEDBO
pQcnnW9Ra5Vj94OAhXZZuLKn8s45Cbko7HKQsRAiXrL/HbBzvSfUyXmnuEKpiI4CgOSsYHBaWEtT
h7vb1csPVufTDBtasqy7xjYdEfjm5pjA4AwsTQMeVb04ZAsm24U+SP8EwXLZLL3SRnosho4ZczVL
UCyAhaIaEI51UFai4PDycTgkQ9XxmAOssbu6RzlKr7wv91SBijiNo67xVI4Lh34xqY3bpnqUdOLK
TbILQ0IrHN4q7lDUN841+WoWXdBei/hXHil02b6Ipx+dYpnwUjzJaAsLQrxuIpZVxY6UPoJn9V+m
iCv9aQPAqMOnEeJMIZ9wYm3xmsse07X/ERPktTVpexepfs+kRatRbSIQUS1moCpclWnANjG7TJB1
eNNLUcfXWzmwapqXWBu3AT2Z6Xw8Al16OawNk7vtA/q5unp+GxNub10GGRK91zm6RRaDAd6YwgRR
4ABXBo7DuBEe9yNC07c2Zo647ZvkpwVIQ/w9S+rvI6cHCagClt2UF8Xykx8+luYiGAUqGY5iP/Rq
gRlsgWv5zFqAxBQfioGeAPyJqVW5REono6jJgzNrRIt7/CA5FydkWEZmIaG10tnnIn3+YmdYlmKi
OrMpdZD+NbbwTp0469O3B0dt7tyOeKRf/+z1snvJKJ3Wf0BDsvMnlSJNrKjdPnsDacGypZAEOjxx
4PXhT5eb2hyhxvYCkxINFfYww3RhDA1tbTut4I3HqTgWvW55bj5XLTi0XZi7D4WUnSrGbT6NIEUC
vCmTO5/GIEwBPl3vo4tBStE/AXdLTsqwpKA6HIAfWaRCm3hJ+pS8lC1IiVDVdR63O7vbz7wegivH
iAedvViDEDcc6qFSQgVEwymK3QZAtyUymUsgclKgQEesjp5KB0aCjFfzOhmeQzuovIv4dOJXwd0A
eHiSrbhQvRHZywu82Uo77lPWL88URNV8e9A8z++2eTCFqsavzB1lhn+dQ6HiSprI6cN1mIcoTW25
w01Jix6IP/9dRlYKsUAOw1IGFTxt+211t8Pstu49olYrOnVrent0mLvFt9aM17zsKhNcJjuTW77O
Rh1Zs5ydNAe5t1/4vGA6Wh326/2YTMrxPaFPeg0TdnwM0Zv/6AMSTCOnAogDpYDn33lSWNqlyTtY
h19kQnmdG7b+xpHlFZAc649MWhLk/2JhFE7HAoMnzVhfPNoSjCu/Wq+B5uynnCw/+Zs61nENLNFA
KtQR0nK1QF8XmvMsRDEEUBm+LH14fG2dk07e3PpSItgXbaNkD4v94VwJMfH31tOuNrJcXeLV867Y
l4cgoBcssnnlKFRR82oXLOjtyI/4uytRVx7fvNbrLZDS7GxGpNOeDj8GwjxDkQmaNI0ppxCIKPIr
YXoTaCvC2p1YAUV13UIjuYouAke8O6awWXSzidmOKPbEdSPkdffgs4uW3iP7rAAHrqlDzoUcp6ZQ
xHYMPkWYFN9KfeqVxnPGXDX4M1JOalPy/1qY77/3IFOR6wer91pCEt+P6TqfjiZFT2gRFwBQeDWi
DPKA5uqe66bvjps94CUvofFYLVaXHGbrpGEiU5mofM13e4TdthJBIYQLQ4ulPS0VNBi5ODtiEUXE
akcWquHNO0whSmSnmE49wfB7p3QkVEWFAmO+2QA6uKId/7LhgMYip/C2uOb2P39ZW7DvLDNug0XM
AhrqDQ1WrHWLSJlw0VI424/gqMRjR1A/ofhyGcqtxblZQeMK+DEqLM2mLHtdCU8tGrDgcvQhUZ+0
tEmjEsszu73n/eVSAU1lXf4ro4no5ZlVLm0bwt3oJKit7qeMYrxQOcH1QwMNRVznj4DP3j6k1Mx0
5bOJzqkfSCiMjd+oUdQ1nDWB3aJVctj45Sn+bbshFOosQZnVtDCuNcCPGiIBUclvV85lYHY2D3vH
D7xv3SCG2vLSOAJcxrIUBo1d/hQ3TK/fbYRcKYdJgPSycWkFiTPcCX1VcCssrd8d/MDyL2SeE9gG
mkP0kf9QtgS36xop/riStUGQv9cWzaH14/wueDsAbSS1K0sL+FsQLN6DV6ZznoNF9R726xe8waKN
Lfk0qbCSsJxJrfxyW0xrjZ++PtgKjHcu1APcx1+cX4Szo6jEhTao0XQnHaNcCEC5/D1asyKWin0+
s1oa2P/0JhJ65UWOZyVs+N0Jnx69it3UWxFdxAXA26dw64twmn11k5kZGhGTHPUi9FeKVwWU+bLQ
q9Au/AS6pUSQ/IVO4vgVHmaM5mTdD+RIRN+hTnXKIT6TzxouUhFCjsXlLDj6KbRg56lx+J89o6vP
eoPCrXKbcS4s698ENm/nan7EUYJdptiuv31ElusvuDmcuDQKrtcuRT8YsVtzcYwvLO6IEmdJHZ2s
WKtBUldW42UrLaM03cWO7PzniDI/2NpbNdSXIdkPrT3wFGJsqGQH22FppyrSyQBtFkHiM43G1xVF
77NxXkd9cL0onvb0w92xFxN2/cjTaui1xIOOPzPcE1bo5F+mB5EioGp4BwNB9xaraEvJjo4cLpCH
bjX2YctAl35VKT1XBYk2Ogc0oALKdUfCVTa79Oddre6x12yjD8z6RAlRBYFH5F0cK6nO+06H802c
8eRXqJThEzH/5jrAslcHKgpM0bV6NDTBCurWfft/s5/QpLyxy1Q8tMdla4m7tqQJtFiTg+nlTWyB
/94F6GXUg+LSa5daJNpIDl6yHRLvXy02Ll6CkNRpL1JwwuCUxhPoR28l+foTGMvRtwUSZD6EPYt7
Acrzl1WUikxcPFpbvV7cubLOJaRMj8Rg1QI3OJkWp3eGBylJMs9TvK5aKNBBWDqaD/HgnvT6a5Vv
/6de2PJXvKMYte7YoM2DV21eBAgbbdj1iJxcDjy2l2oSDkRTHiH12/w0L/QIL/BMuSOdqkP45+0j
UgFCbzvDXBQB6eOXVlXvnJs6gHced64Ir0byIa5p2FyxR7JiVhq2izdTkFxSCVliTtI89WJt7JGP
Jntep9FByhntHokEAnwWAgH6Ut2a40DjzExvoBNVnu6yDos74dUBpQkRNE9TfqJgCmPuZSt2V2lv
/HjV9HpUuJ6e/4Zz8sYoDWq3h1KnxbZvEpG9SqqLQsoJ9ZVHs4C6KcnjMlzlrV/KuOce5dyUQbOu
8EhYX+jcw8CzMXYtF5SDK0DRdHQFfWHU7rf6qwsmPx147K3oqtF0Rx4cd10EnV+yC+eAwHnPumee
Q3Vo8/b6H9J42ByamIqslisU8UbxjKxXGi3ftDq6FoK14cyK81nM1pVpOrqgA9RQlpL3EuXgVyN9
cjMJKqkAI5My82DolEDNHbncPozCXAyzkx1aK0p4/8bnb1O1zv6taX6JPSi5Xzcyl07Y7H61o+9V
wQOcvlpuqHRTJi5lu2zmxPyhogwO85csjBHezV83jixXs9vEEzD1Y2z+QXTbWlkUmkCcjjeOp7Vl
tAggi6ETPEckkQ8buqse6q30KQvjnR4oT8+4+nqfgwe5dFwzHRe+l0DFP1+GlC7/qDkB7nIpHnrd
qhVqkeLV65o6EK0VLyK+hP4ltdScwQRZeBdzS1mb9dDzqpPHSnDANdzmOoaqRl0dDRObW/D9d6sc
750tV+r9NG/uLav5sL+FMbLMIj0Lkbe2GMzUNQctA60pABMgMPIunfQWyQVjgL7aXWoP0NhCNro8
8aaQxWWl87m1Ay04khD0b9HnV6v1sbRQqud7zvhPA01uC4AR/VtpJhrmeTg/3dWrRnl1TJRTXB73
sCYd7VN01EOp1j46nVVs3ViPEl667Vq4dN1UEjiDh+yo3ReA8o1kyGYEFOXxSL315QBL7wx0efGT
FjLKV+M5nwA/eAKIfpuaDGYEtgwaak/JXbVPKJ3VIAtfyo/XcDFry0+C9am2smlEOGjKHjnXtVM8
F+BvftEenwns+bB8sgjfqYQfjOPx6/5DRQq0StR4D1PzV9QgSIu/BWiSSsmxGWwk8q/en8vZUg8s
mdaGQ1/DzCt4aTTUQCAA9TtB1IvP6fbUvL9bSlYLHh18dxRha34Wl6cu77XiBILS9/3atJAxm+5i
CgvLin6q8OfjiYT619e3EyNWTzFS0trjQ6pewDCpHbiyppJFIbNEFJvktBwoVzGP7TjaBakgGYce
Q+X7NKZ0TQGTXabxiJxYSeetmCGTDWlDrPfv1fAstHKy+qYfayQU14WBSsdhk+LDUkPlIjFSdKPR
24mHfB6ip8tx/+nTtq9ibSllE3bmSRK/6U35dgQYtUiVUFnV8s3guiFtwS05R254Q4aXnfX8jd2s
DXbdN4LCcRrIQ0UoKdyHoCMMBjLpLwTPnbEc8PqhFwZD6Rva39Vvgg9ug05I8wbyKuT8wgmG0t1j
ivmSlje0zIaNpe6UQ5Ayls4kh/4BPO7c7Vs+YkHPdFzgJBe1zo0HIXeSc9S2dsJqHfYsNg+3W6s2
5MMgtLVXX1GRWU7sCd/AXrrJiGVPWVCgmpzl3y3TzYP/sPLVFXETvmaeCPW7Ti98Opkw0zNcViKC
FnxKciEMWrUi1UWnKAB/FdEZwCICTFhdjU1+pl167wgD4GiRocbJ+91XzrIFPDnN5EVsoTyDhl6y
JAFm1736YEw6VvgUzk0X5KvAUOwqUxHQRd0agIgAvp90oMYB79g87G6/AmKNFXCYuk99iu2mXy0x
nYsWLgiMcUkyKOKaLUaC67wEfVBEIXFh9Ee9d60Z4Ioi8IEnOsD741gOEGHVBZ8GciPczLKfJDQB
0Jx6GKAa/uTB0mQWS/kxRKCIEBMnL18QZQxE9YgYasvrsx98dwunmnBEfXM7K4MkaMiIgd+jwizk
4SjiWKMWsh1pY6aXPghRzWhwBVjZdrV/HO/L/abIHFsaUpqPqBx6hYCgEU60/IwkUSbNAEoi3aaH
z6l2CbUlPSnvfPlRyRJYeGV9PdVL21fhgna3TKpv68IX+BIKk8BRdURyOUuott+XHoQOw5o8vhR8
9x90QQr9GkduaNM1zBOzwmD+j/PkeJnbay1e77ckSo998/5oYXITK0T6lF7VG0Yd8IFbjIlnuhWo
6sKAI+hXTO1VXeik0Gk+cdwnK7I3L6WV6zKxSWin5DRPYqqCgaA5ZonLPcPG9c5YwjlI2g3ByuCQ
ZbG2YtmorU7AakfVovGq5IhJSiKHLZdMh6C6wEB+U1uR84qduOOmPAXvV2KWXDV/rhTbPyOYM2S2
uiiiYBjKoKkPtwSXg95h/4KDarGyPHQdbW1/yWUffU4Uulla5O6VdDPlaiHOtWdEkuJxaQdlTLaW
PT3SP1zQTRs+e/DlB+Il0a3gg5N695Lu1HhzJ/gf5Qiu/wqShYK7lmqbuJq1Ut/fncZyUJoyFM/S
c91lhmHS8kuHgNMfaDQ6Z0O/lWsqc0GUPM+0JxGSM5J6OSlkfdGPLsmso0fml30mEXte7JEsaVhm
0XBvDMNVs3CbY67J8+7q/yRc/UmHxVxNpQrZ6T9TauVfZUn108AdWQbVxgUPIVK9hsz0/iEDxaDo
gfk9hIJok/vTZyMHLdGKg/yZGHTdQrrmSW7fvtHf3LqI3hnPtcHIv8yPf2gZXsm2V+WvTwdTE/8j
WLWBb3qtxh7ByFa+2N58Ss0VKZ9QA77hiDIqjrS82/Z0kYIG7UKBx2hm5kAAqbhm2+QG9DpkIEib
Dfdefxg/RmoFUtwiyVU567g1GzinPHXoVcSRYstv7hH+2DKlQOcLYo2Vk7DaXaL1cYenwYR0oVj1
Fa86b+3CLvWPCVopsFvMNtc5ufNrbg4lYd0Bl8UWnZyeq8Kd/1cnbwX8dvpC+H2DnCIh3GsC2Nrx
o6jUloJ+Jh1Zcoy3yxF54+l0LfSL6ENWHq2BVKlrLkFFNitwzXpUiEBrdkJ5VLwxTsD5H6zJCj9x
BWsm34TmraRVtZG6eUZvKH34oufkhvFMALennrw9LT38dNKL6V7u9xmk20fg2YMNU9PEQa5urkGK
IpgeYfEZm8IUR1BaCP1tfq6CabI3fHeob3+IuYywcRQZlHVI4PhJROu+9FK763YprVElPZoA6PGm
Z++T5HuGGqg74z803mIFEeBTs+niV5jgL7bJcGIwJrCUZ0Xph9K3dxQHvp244wHiqfXGfBpk54uy
aSNphHPaptcLVHgKLfM3W9Y+Ae3KHXz+0VU6Q7uVzR3VvsPbFW2UBcfanpCRlnJbwWeKua13fjhG
ajNOiRLs4VGjwIXYdQLZ7Vnk6wDDHz+MbyQVD+Y1euGZmscWhhhgmB2mHjttOVGu2z4UeHWwLb5F
9JkcDZPTzsFDg8zTQLuKmpZ8L77sDo6MhlvAw7kUAnQVs5z9xkLDfLKC7I+1+LWAId1z/wtDJaX8
6AEUW/x4DVlwR/LBZxW1z/0VzGPBXerEHtgvfixClbw06dFqA5usKVuWEsFPLzgEr+rxCiDnQDqa
5E7JFqKxhcsDJwlvM9MH3qQVZ4f1ouHqTHKlyrjSYAXjsSV5NraapTW08jGsoudkqDYMA7xQrXG7
fpZf5JqwDpqECVHYWsVa7gJzgGvwkzMA+U8Fb/En4PMF87xQtG7PeBja1kwpxMClCF98FORiIQtN
njdFQkajq8PSQp9HbmEJ7y0fGe/Ryoyogxz8C7Rc82SC/u4i/rbZvVZ6NhMcy1MNRj//SDVwnlZz
Qx+66daKrowPK3Ze2PyZV3DnqBMX7Mkjin+GLO6pcpKu/WsmIw1y/ze/eE1bk4JgTSHpSJvuXd97
0f+Yk4Jqoerh6o248DJQE1kSOhHN5CZn7NlesqIJSmzHkm3W8numjaF1jIj7L5t/XPxjeM0wixrg
hwySvPgRBz/+kWMkTY8W2UJlO8lU7xBAHnG4lK09t/kwLhx5GgME6iL34kfNxI/X/zjXvXxOzEls
uB1W6VNyzKlxzmp/IV8mP4qntU/jcy+cUX38jbzXfHeFy2gWrnoM+kNs2eIEtr9d59vAA1Nnj5kd
/6oaENsfgUVRg0h0s0SQ0ir0ZfDlnhFAyvvBqUEijIxvzoqADQXp8fIa++r43BWwiBQzL5XtZuCA
2JK8LyRfLpblJsG8w5TYnK9y/dqZgdtRYeIXYvNx6u7nTIQU+5dnuofwvkQidGbfRASEteRtwaS2
Ay7cA6Sb1HOSxmKH/oDSR0Bp8cMCY4v4WV/O71K0SUZr5QdSOnK6jWLlD9b1GfQ+X1LyUfH8fuGd
Ox3px3Xs4r0xv0NQOAOLFZTe8KEnJN2ODKJZt87bBUG0mv72+FZpMh4ZXR1wVJNIJkEZNXwlbcY/
Jx//2ksFAujkJviCMlXAYrhmyPEz8GnALAAT/YSS+fzp+XVlEbkZuETLXo04ZvVUX4OQf2z8h1eX
IKJ9y//xHW6BmndCRu2Bz2zqDIWeB6x8NhJxoPGT64hlAsq3/y7b++avWL7hpiHwuivHcenNsqMu
9YY8vWErV0uHz3ddSrzPRMhVR2gwHSZkAkMKezNAi0uyLvMASTmfy90PaS36EKltrJvHoE9+Md7e
4eXRez6pVqA4+nG2H8a5DavnM+gc6cYfbtgwxKiN/dpbFJ+dwCtGIZNre6Gf0tdd6dDutGaMEClB
eEB/6c5rV+wh1iCTCDoRhidXBQeCqW77L41yyk/5SKEDyoaCOrVDyDX3bcU0sCe9yXYHXKlfzHib
IG25r3RK436W8+9bhKZy+GIUTS+6MjYhZjmZtDQKZff/x7e5bC+VwjN5XHJaKI73LM8hHVewGgpk
uz4hosqFxLccWzgev6rx5XH4kj/tZCv6MIx6IGgJSaOSintI7gWhLfnLNO/L71uPXWvDpmfbKPA0
ecuo4eW/arhP3vn5XHkYcYeK9Wsn5ANhfF+JWg751aX5rqECSt8YCh8yLnisBmRWBor5ImaZAdTi
eNGYK5n1q8O17dYmh24/i+S0YBNlDOQC2E+JryBAkhqW/WqaxQl6+yPM+qqdHvCoGFIR3jtdtcS+
J87Npm/gnN5jq04l1rMbS0LgEWqm0TyvI4UuCjtSe6ObYbIut3lSqXVRq5qrUsHimAVXu9b/63KW
AbUMzcD/DE0FdWfJNKc18iVD7/bxAXtzj5GjZUewU2IHyKq/+Q0BbhcWg1qPvbVGa/Jpwr1hM3SK
AHbnssrJBRQ8mItVtr5rIhMye0LbSBVZ68EckPfjkcako/idYHn5WeuLJcwCymy8aimTuc1RJwV2
qCC+A3c3MFL3Wcjlmozuko7i2YbdFl7btDjvTAS7ZIsZv+b3CyzhkrAOdAULh0/CFOgNsStrBJg8
vnv47PsCyD2PtRmDPgbsJq7JNEcWYiP3tD4dnkxhpitbN2sj9v+6Dv0N+PNmSNYjvbWi8XfbK7Gc
1qTmvPerHLSE+cUiJYWFMazxVINujuilfgSthJ3fywU2HcEiROamh6MJBbfA9irtiMiYtzr6PyoQ
4SUOdfVmHWu58/BvPqCTReZP+HrsKu+8XJ3+Kg7hRIojfu3AY5vwFm7w02p/ok21FaYW0txcaKmK
neJokYiP1fzRRCkMSgMR3y3yxnuuJu0T+EAWsq3WYTmrVi5f9Hc4C2JARgmdhd6vb8dKGUcWm9/L
wQ416BcH4g2buytQ8vAxGTRctQEjl8gbClBn700Kzp1W0Qnynuuj3Q9q5oVh40SR/tMTgUNPeBut
8P+j5OM4jYnWs5slakEVw8plj9arVADBKQn5HTwZyOdqvkC3PAQqb92p4HY1xUl5EU5d++2StpJE
/5merr1J4Nr2+8g7auu+jmpA5a3gp8zQ5i0uw5GqFmRX/CRh1M4ykbVQaFVW6Eac1/2j+o/pIcOP
4lZRdyKp1DqsBUiuYk1XQlWhDv80Ejb4SFreV996Kpu03DYB0pzH65Ks2NsUKmQBRHdQXaXG1igf
br3wFdhtyR/yGBgwfRvSbn0d9/yBTFUdj/Gnsan64FedG5cJm8G/7MJL9Ea+L3u8miR0hyvxi8y7
zyoJ3Ml7eei+b5frGRXRB045l3VhIllE5mq7AVNC9UUZ8EjKaPMxETHpIsO05wy/eqB0UNd+vGv/
0cPITdGvvhIOySCOdPmPu+O+3xG5gscin3lxXVlLo21Pt0/aC9dM76BhfBt3HpRzGjFFFrHwj42M
F7YwV5YHLqaSIapcQN3xchKiB6M0+dDH/YsxBNCu70N+hws5s4bCat3gQjluHSORMyKUxW7tuefQ
cY+cFWwuOfz0tbWPxZ7SbVdpEPDj88mLZmeArB+ajE53pzlNo6I6JQFhns89Uf3de0g05AWduAuk
qLUL4yF5uPk1um+5mEGxsxGAVhzVSFhhCYJ9NbkUoot39EplYd2EMF+vUshLXukq199CWYq2BoOx
iS3Er5flziPHcLRRpd6br30chBavVgxx8I2RZ3WL6wcQaVuqImA9QJQyOKJFlRz+dsx5/u4a1mPg
LzPTx3kCQ1YQB/DpK7sSuhirUKuCnws7mmcBAHiRbEvOsOosHuHJLa8q90iGktIJdl19GPF0nHzl
Wcc6f5wdxLf2Ik4UUokrZEcTWjHGTN1Z/sKF6uqP6oL7Ai5g97skvoUv2cGsWYiIdvkgkDNEtK46
v97mR1+0vhJvjveMvFxYh8EmJi2e8HMmc1eUDUBcD9CeVX15rhjz8aN4/w0FFrc5g6d3+2DjIE3V
c9mZttCNassyhKw1KOPmZp8PgkKxhrUPM8xTjO4mIh1qspDurhjysf9lDa3WmIaIOIGELALSxHnq
OH217kGGUaW3VKqCX2qvNVgaiJECX7yuwWsOO03SJ3O+cP9KKQOMVci/cFG3g9ygEypRyINi32uG
jqgqFH42yf0tYE1fkpnEd1wLkEBYYxdsjz7stq9FFv16H+5XkNTeQAnd0pnOYf5PUrSqT1ADP9M0
B8mheTYff+ioetZOzsMw8a7A1drJswzbPfSnC87597C+dSJgvqQn/VF6/zbkFIm4hgO0GUeuivTJ
s8uR30C6LLRn/SCgRMNlhcFMyqbvSR+3OJxXXdn+qXUMs8EG5xn7X8O0W+5Yb0xB/ZMnqWbKJgag
sYD6paDTXKVWwcHGS+I9OTUx4RhV4ei6jZe3z6Prc4i9MIAMzFRVRjt2dgsGMc0YqVGzSqF/zPC4
2ugHPcxtefhNUbyS6wPQCl20y8A3C9aItAlnYwYXyrQQnhLNMmoSOXhvG6uWj8muNSKhCKVTDwDp
FLeDGNx+ErRZLzrmf1J8Jv62pK/oGtL7B24550KubIz9F1zJ1F9lAiuiF24gY6kR9LLhFgubKVCS
EeQJJdZlNXPXGTl//Y09J0BexZtE+mlU9H++jKhZvwsDbwSUrTAAWi8UwqjAO8CLLnGQJbkBhsPP
ftLsAoVRPMuJGcsCUGLM0zpY0QGOISGYhQidMuokM3uzpLj6kW4v8g7EC8jdN4ntaTbz85ijkU6F
Zd4BFiM93Z7/lSGfFKhB1yGYSldaeYp3o+G93xhzCM2Q4rwrRd/KyAE3WpFo0T6uHO6A6YM1c8m/
BeeH1IRehR6CN8f0Ueso7gPlVsPhTFbc22x59/G9jdy+aL2QDbTn59F5p9BVed8wSZEDduo1NR0j
Mwd6LibOeyQLgUpsNcfWKbAKSHClCVWTjdZqUAt4RkmaIzd9n7oijaTWdVQ+ojNKddMiXXr0bUk/
mPgcyerd1zQuqrLXlMzHM6Niv9iDnBeCEhIjGOGOZNTxzN3slfqcz+NOF9u5lHQaPYPlILKMOYmt
0p9xVx7dKZKgXNP4R6PG/cdfhMOiaBKiy3RISYkA5bxt2KgJi8f++yztx3x5f5+yZW+Bg3Tod8FA
oEK39FWMTNMwuZCZI6zrmmuYBb59E0k3dgJqTohpkfQ07/4T7LJNgRRXRhLRW9M3S/TKJ4gnuj9Z
awBzJyhi+Vtswj5ELgBEvj0O+2kiq2GSciekO+NOKH4T6U9NYJiVKmh3YRHeUXegnCDFp/u10Tt2
3hoLdjRonAupNPpCP0IYzo18MxQ+wG+V5yUXHJKvL5eCQ9k+4qu4du+VbPradGkCf5Ky8ou6g9QO
YXomY8HbOzP+Szn8Mu+bM4YlDsrOO+DmMzNGKX/21CowGmYRW8VttX+5FJJJaD5thbiyaU5Gbdxu
ZBZXHymVE12AstxGR9A9uEhfJEa/Gt41Ejhc1zxudPtvjdf4zl4bQbV2H5hke3pTcZpczJ1pUmZs
s3ZHgqATHg89nVgSsd84ZCjCoNI/IznO35qxYL1SCq4fxObsQ6rerdI6pY152UxkrfidqaXJp83e
jdMadVJpNF2reoQeZcXGltE5yigTkPhZhxdqZQSyVOFJslG+vfEHiT7CgvxuPHdobyTCp7WtV1Ah
Q0BqEL/SLGhqn9BeTlTJO2WRZYRu6Bvq2HTyodguMIc+GqA1oSvyQPeKI3foYSGtWa/hxNru6uoH
/bZaEyKYlwpjCYo7Klj0xMV2ZBAwYLYEtkls+GfGW2KgsFPaQb0Abp+okO86kaohbj6XE76JYcIO
f5YavKkR7SlazQslp28XSylEAkegklHVzfpNeUHyRyRMUhBUCyr4CguLF2OOfbO/wPEQeBNPtBfa
NveXqvWSScMLL4OJIr3MzD1YpUQ2vwpf3sbS9bbQQH7EEoqKqPRFSzaI5yn9pNrVgZPALLmOQ7hw
LuMJVraxswzPnfB0bKPe4BqVFdDIH/vghFwsKPAj3qxNThZ+bybqTYg3C/A8yqXP+EHjuz1h0yHo
OX4aTJifYc36CsukX9UQOn6LGy5mWYDBqVAmbBJxZ3OcHPrVu2dPVmUaJmYRrx3cbYtSGU+d5h5d
W1ZgO4Dr7nqbYlMDrgyCUmcETMkxRamr2D15ae021hk5TJkhnEduz7Ov4ipbPtkvHk2dxbZTp6JP
6w8jpFQ+jmcJaXsEA3GT1Pwx0y2pho0fIiqch0s+0gpcU/1a6MQpVFDy9/I52SXrXXyHLVx97u5w
h/72BOqJskF+zZ0LRUO1Y9+e3x6Aa5k0StmEn5BHm43V4gmf4kdkFWFsNvgAQbrFyRsDTTv74zRA
ID4QdjsXX97YT6JfbMHk732eRUwqqacjJ9aoolwyIWB7XOw+eLH4+oD1efhhwNIXe3wyNZtdSA/9
58lSgRqOOgptSJzasB/oEjoBjyGlkfjcZIEr2Kv45t/KohLBEP/oeMTOtXXtzuYukVHVaZGCnTzr
+B+AAbLN3uj3t2FuBdy11pCd8dyquDeEt8cKMKFH9WUXp7ISu45kY/5S1gaDbLya+MrYzQ8Y2piX
8GtPIfGyRUaeA4OkuyWMqCWtIWaECTZATRwhqnH+YjDs5yUGLCqt9wlB2SSLi6pxiS5pFCjfq5oI
FEqC5qzf87UaXDZLoCdhuulTGcwAriMptaHv7czkLtLPt4zOIGjU3SfsMOGnnsdUKJkFcpeipmNO
p78RK1q1QOmg0vkl2xJyqBrUjQr+jtW3jHk+89r1yn/H7moIA1a5v4h+zrliN5DJZSpnZpp0aPAr
n1/y9jow5aNnMaEIqPy0pg9ank0wlCN3bS5TTKlulJ4OKZLVPRvuq+czim0Q4M0izpWE+ZcD7A2s
8aFErFBVKpFGplr8Te8Sr2xORtRAKnMIN7ZTkIQ6/927yHwArzxc2xdiR/Nke7LTAfBecDO79TLw
hXQg5PYEfUMZC90RVd3xlQYIHqV9ZPfiGBRmgGQ/AiiRn+/IPdxg+48wl5XC2IrxI0BCFiMLFXnq
IqHj+LXpFspenhPs3SoeNOrMSsqP1DjUmI6bqqwCXu5Ei/7y8yHkHuUqbDph+QSc7F+LzuKak7wF
TH+gu13rxujDyS2s8ubAe2DB44+SjCmeDg/w9HkGk9WfQ9AhUvFqtceuIJR+P9f7ESp2viNYa7ts
33iP4E5TXaQrVvQE/H3/LzVCKKHzl3gu03djGXNFXK/SNBntS169OUxfusZLMIPJXm0fI7z8KcnZ
SgyfXSxbrqkuuJSrwO1cJjlNU0Enj+7CDgwr4kwxYuMg+YXVSBCifpyDYjUXfHzzfE1QDkWAqWZO
lCqVMQDuW7W2XDfrEVH/fdbVI2TGwJQNyaJ85ifLM4yb+D6WOYbHSaThmV+afZIdy0LtBOlZ1RZP
+x2F0F7mUFf87y4VdVmBB8O5mHM8JSG7CAVj7CvIbgVySAvTMpxBA5Yxrk74xsgUUbp3yutXvot5
a079F8LYOSLMkdc2Xy3yjemQyYNrJvOAR/mN+GVFhBlqPsuaQq8POxKPFUnUxi6I2JvbYuhJ6ebr
Gg8dmGm47njZZ7BRYVbYBDpEeBmqIuTafx4wc3UT3cImw4jwsdogxwokgSfCVz40zrG/5OvUUB/W
FiujcaP2Jw2LhxLKqFd/Vj02V79i94rdsBcp2E8s0xhVjMwj2ha7WOAFLkPqEiHzP/7NKods53z8
A2BnsJTi/o8HTKf/USns58oghriYncHFtZVP5wS+Y7f2wn8R0UcU5ychBXE3IIzSScwtFrzyBPfO
KsHVKgLr3NMGvRMUAc5We0xVS06x9QneQiO1gZIsWOVeggCEFtTkuGEZFlClSSRZQOsyUFTJ49Tm
OHwjDlRJIns9hkBFmu2Iet0/QyFtGWsTvP+NQj7ZK6k+81TH44qT63x2Plwy4QviccZRUwJvdY4T
LjlcK2pYxjPKV37tMF0Z9/Q6DZ6LNkcG6w8sLe2RZK7jmC2YxBuMHLEUpT8MEVfp0n5cdhp4CaF3
Nmo5lzPgSLLYjhUDNE6l1RYkIFFCw2jQ7TEdIpsJn4AfNUvvTsERGW5LGhinNXX+YEdBUxSP7kRw
roj9eKxMpnouHWFWaV+PE6b29nPmBqqx5q5Up02vbXULdaRZeniYWIqLdzr0HXOwT9SeOYsr1BsP
zistrByFFZF+cw/taPHzypwRJ8jMdGmPVY3IT8dR8fXEMiolZnbOIOxTmq2LT4TZhr8jx5c7s+14
fZzm7Xh1hQc812USUnzkhTDcytmvoOonXUojJZVxqaC8DfT6KmC+rsHzbe2FfoX5/vfCVpC/CXtk
Grp+jih4lkwsgA9vy30uoBQgZ3zHgVCaGL2h/GLTsG0Menf644Qy34EPcYNXR4Am782L3TI7mTqF
3fOKPihHjViWHdfXOeThCFdyYo/pQGVNu9PVCiVxqRvH/4U8Cp8T35kvHUA8VDc+h/gU5rkX9vb0
NqDACHA3QGKymymED2UqusFlTxD8gmWSkQRdvpkvggSZkz09ahlq8zMYdqzCI7rU1WvIgaGacjpF
2kyQURFDtfPn3abozuMjWxaeIyC7ISIxyFuNKP4xDu81kT57ESEW/CPgkmXPfVbMCDznTSz8DvyM
t5YAPwQYeKmTYt8fguuyK7Be+PXtz1SjVofimKbcZXkfy83fkX+amWWdNVdKbdA5tOi3TtmnTZSr
aURs0vb4i9bhA37PeGDXehPWTvAXjn0TEdHAptPr6KNbnU6WYqHkLu/iu3OhrS8b9S8HDPvAMiXm
bcmzlH7G1KoZJCf4+VC6xAJoxNqpuv9RGVOpaEwb6stZg0aciFx66wuMNCQvelqptFB4Lqb2hiaV
I1U2wtI7cOV53vnV54ahoahuY1RgcEcH7LfN4Vk55IHfiwH63c1It6NHrgws0jowkivWrw4VJaO8
vz0Y/apirQ5QM1vDGZcbEAj+OE8Sx5z3J6mZSk31QURddCX2CVBj43I1iXCkDsagGHCIhdD7xlv5
hNZHlZrXVy/VnU0tN03fApRT/zEshRo5Uxtf024H6LgMZnXd9zbOXPqUQgWw0vz5Z8LYoeajVItg
+M3xeth+s2NbU9SsjAxLoq7dbZCJ6FBKHvXdYl4odhKPw5LE9iRQr4JBUElzNV0fCkgo+lnMzrmV
Cs5/NnokWjxdR7as3iKPji9E1yg/acEruwCQ9LfZVQBY7ZxpBkTIt0dW/6EkvhChadejpa9Ii16C
lRjgX1vtSQ13t00T2xtls7POUwu8NbZ8QJHz1ZVcbVz6lvHzP6+yQkjCiT2Tdmz9oy9D9SONjScX
6jIfjUV83UVaPc+EXa62KGNIA3ZrvioUDwDrNmnRo2w56wj+YVg6PFW+phmvI0TwxpL1HCiGkZdB
gLd+kTWHHqxRohScY3BTaOHIHWWa+izy0pu6RL09VU1NKYoZYejUJdh5WP3Es+ocmlcurdVxaHmv
2pKLkiZ45FllFse+aosmbuszBSx7vkg4jGyTnT3SWrlW6bPPJZzu3B6Pst6OCG2hxAs/fSmx541/
pImf2kMuMC/GuLXwB8lDtuOKbf7H74Gxrw6eUvshIHnFkWSgpy4jTMLWa/YM1Wy9aRK+Z+TJMsfb
k+2LrrAd/LSx+1C2VTNQgDPsb439TFhoUO9YSZ9OXVDsOdpaNBd6zZGGh4Rnslb3zGos0Jigi34U
HiGnTnXQA1/576fAciIzVEv2d7V1BC68kuIPiLTzt3ueEXcIlmAy2mJ0vXwCFh1+lq+ASGvtAFT+
FgDUAxcRfmkUDNr82MAMeTMzBT1VMeXhcb1kG1jm5XDAfObuxxMB6gCp3OF7PXD650RXlg0VoNfa
VTBo3wryXPMieueaMoCkixbm3czdzXv174OTz0c6Dn2WswkpLBZtexZjzT//Z7SW37sWZvAAhQPS
Ze4cWjRk+KO77mZ7jiqtonOjl7YpH4zH/guaaJjSujY/beUv0lpSdex1xhcPsoXuShQ/tZj2wAHL
VBIVuQUu3wN29lL4fwjZXIGh/G3TFDvQgLEfUuu67nuxf6HChBx/4d8IWmS+RB8/zrJuy/aTWKcR
nLsAdBK6T6U0dMaxFwyFzRaq6vnTpQi7DOruvs+ubALNuDnf7vPEQev2qC2vn/qJ2Hfde/Q4DV0B
C2O/7nMFDcoIOzdHudWyPYnT6PZ2aXHJhGSnzeXnZS6NZF1r67MSa+5o9TPmssWkhqjGsLBwumbo
inniVC2Dgqb11uU3cdd3p9hvudCFiMlUi9A72FU/fcoH4DMFBbe4N8M5fXtekr8NSGjFeeptKsuZ
e34MwckxnE2kwDkV7iQp3p4GYimBqrzaayXlWiwRrwRP5l25oxeiCw9LJPFW8wPdg1fGl/l54NsZ
JSvb7wUT02UrtlXoSGj15DCkHvnE5uv8J+BX9TXV5+4fWWM46Oe1fO/swNmcEpkWrixXel/91PVo
uN0mr3zAuXw2lVKHafTqw8+NGhAAEXwLgRSt+UwW5RQ/HrbHSnhA6hjeaDRvlNIuQUYMAcJAa63K
YqWYltYQhto4CuHnWr8OiTRBhxkmrL3k0FFFUeEMFEpZqC7EcHtU3A86jzdHBhtUsMmNvXJ3ybyU
EF6LYVvC2GwqI/5Aop3OrFapm9tcJo6zzy9ZlvUFxYJRqkoRKd1hrF8VUsr8pysRc9Tg63sCsjUD
cvTkYfC4LiFePVUteKO6TGU+dc8NsmwEJHnGLqGX7OElBztGljAFr4QTzeioB1ONr2iDMkoQzurX
lCFyHFflLBI96ASN8b36UEeocRZ0WG+4tFg9I+PpoC40jPcpnO+N/cmGSl0rczERi8HlRX4QF/0F
b+77PC4xkyEn8plG7NYJ96sAq3RplI6D2OEIukbvbIwlaIiWUY+xkJQg3NmYaI3eB0v+2XQR8x3J
zUm01PMYVOD3qVmu3MzUi73/gJAbHRLXsnPrxbbuiZ68x1iCBvpkksXOMs25kJW97OtTYEIZS4Wu
SpB2jbrxYmjUfnJ6Mhw8kQaUYlCzsFDorYat7C1Hzfk5ZxM96W/ApLmg4Pf+J9cBh7HiAl1s0Kxo
KBRdo6+3JlkYb1e5PaQlBdrLmRCB19IHWAv1FlvgLf8DaeSCDLC2/xEtDA8mZLFjNIgwcC9ctxfp
cCjk3MFavLlUkLg4MBGxFqHKxFLON0YTX67/c1otacTbhksztlgeVqxNgo7VwOpv2ZiYzUzZHELI
lPgimKchmeqNIGfWzcBYuSWscEm8YWr26qiyXg6B0iBlVRpnYQuXUGhyNPVpejHs01RwpgX1yZs0
W5XOQLxDU87nx3mZTjydyTaAJ69WlsRnneJjs4/ihZsMNdBS0wnKH1gRhEsznHXiVPEfGN0voV4s
nd3qoBvPOn5m7prc/el309gPjhVmWM6zFKJDQ4FzeslO80q2BXxR8jv4KI7ULMFeUEUzmnCJJM3D
EproeWPErwrR954LpGitiXvb9Fmau/PBrS3rX8pLwzK8t6kOgAoSPM01zT3W1HaBnjtqd5IjybHe
I8XNseEtcEHAgYOsqhdR/SLMwiI0lTEmaonrFLvja/DdcZNwgYTjeHO8NPe570fv5g26ehH2G7cj
ht2okAiZaU08Ex9SOifwNTRqhry5cabQ5F+PLckEz5q+bKvRuvekGqJhe4f2gNNMO+rV2UMcWup4
xYG95OtCG9ABKimeWZYENWfheviNzWmDM9x/Pf6xYhO1/ZZXH8D4pOVczWyaVRsCbZ74TrjRzW4p
TgC3bHn0rOHBNqq4dzBsmigwhuzHkWud2H532wL76yQ7S04cE7gSsiUK4uQCbmr7ASAEajscBojW
lhljlnyxxnjyR22fuv4/Jb3Cm74ln+0872itOAoeNs3nhDX62D44k11DbsMEfkZ4O+ntYxqYR6wB
8j/CJ1qoTb1nOkWRb8daPWiCcE2tdB8PagYs0gkO3rl9Vn9ubRMZo1ACFQllAw+OyjAWZVHnz2k6
wcpi/inWwiXC+tnSGYB1TYLIyjQ8DOAWC4Prs2gqgSUBrkbmbZMRTJGB/LZaSMUGM+M2N16Dy9w6
X5F1Aw3L3GOwPLmZDK4mRJIBplUpVjnwEYL1XjZlnsRl71KvvS3iZBU3W1EzqdZUhBM8pISwWwOR
aOxxKghVN41uxPWNZOpU1inr7kxF9S9EFnCqlcNOku2+514Nd5cdmThhs3SQiFn8hNDnzCutIUJW
lFSuhF2esbG8w3CxS4+epf04yurDhqcI9Per5mpASXXCd/5PHAuNJ33RQsiRPeqHP9nwDI8wbbUf
K3CLFnIDYrtuvYYVmUJ6qz6HPp2G2i+xB8AT0AtIEcNSfTl2fCxcRnspb18TQ6WmTEtocDApQd1x
uj8WiRJQtQKyBNvXzVxJsfX3mb7HG1pR2u3Zrr7jWqfeBb9N2O1ZnQpXIMAVgjT3CZxEIkZo6ZCz
C/NRBW9UvdWb49YhvOA320paxKSBzW7HmKRQd5lOFPXNI3VYIipDRZbKGM+bh2BwJSEIGqCwPprT
5pCFcKCWXhYrltq0+VE+IQJAKvRJio13wSfrhVdI+mMTH+PGGacPJ3vVozU7RG1Wo59r6Rc2Ue+F
fzaKuKKAiVMnuZOnS0CoxSOP4gu6dDcd4yRYZ3Yr+OnBhVa0H5LlTxG3Dc1oubWv+bbcB0RrzvUN
znVRy1UljjNPHwuKhLwhpP+JbTDGxV0FhCxExRIEYK69ahe1g/9ASgFIfdlfiiVvCkSznKh0WiJx
PouJodT0X9IH3CzVu7WWL41/W91gCnFfV5ZoEL1T11MTl7OvaGCbrSVsCWY3X/FPwG8kWjnN2MTl
9df3/Ghjx2K7SL/TqdUp30PSWREt41uSQnCm62OQtGwcUJ+aq699lb+dghih7YKRi+eB+sxVTA2N
v3Q6Ft2PCktVDL0Mhv95Jxz+6is4NYuddZzBrpvXvRZgEjyyjsMix2L7jmHkeadxVBAw8U5hRR85
FyjLx0JO1C1i92pgfFJd0hpQepRlh80FNUyXJfa9ZBxfAJSfck0gckRF7DBoboty8HGT21Dz6Ppg
d+Rmis/DSO+YiqKyBLKbEp1tglUXaf+xLqDcgEgQGUvwuyS5T6viwmEOOgEb3f1dr7voR5ZCIJW6
5FtqRWShGwVDhUxT5WCTRvESCteWKBYl53Hu3iF3YzVWMXrrIXdr2n9rr3Njl9lz2pOAQRQi7x22
hBtuWUGZbIdOKyWwBMag4YUX2AbIXul4dCpdRC51lap1SCyv262YH/YUDw15y3XjYjNfrhzNHyQF
GN6ORjMpm7EPbnlxza/xgYV2r9347AAoec/vRGKI+7jwDOdAjgni/BrZBbyhGDZfGZNYCgLK5kCR
bBf7zTyZySt7m/ll/BwneFX4HIhDf6FP+aKHJcICyCub3yTGE8CP7my36lR/efQ5koty7A7Cdk55
OJ6lv1IyWhWMV34oSmbw8VA//q8uNUPEpEcJGdZiSv7O4Au7af/Fc57ugcdrQ1BqojDfjCubzyBi
yFf1QiPSm+Gv+DyvYfBbycjbMu3Q7BdGwT8ddYXA8nzPvxIsSKGTHxw1M+G2UUr4lOUcRuqm2plF
TvQ96DVWWGXsNTKp6N5V3YiCLVNC/zErcriA2DlVOAWJykdyBrcpis+YDJt+Ih5Wbo4NTQxsin8d
3bu2Cv/25+IrWc/M35+0zhOAj2KfCY9ZOUHycVwrIFhu7LHpiS4e2z6WR7IbPJtywDrEQhStOPqS
pelDBDA49dKwZGqIWb2gsiEnMStv5enACsO6VU9jUnCqf7SaadmWNA5mbHxTM3Uv2oPLYsrdgkV0
AoX96ndc4VUaKVMbwbYW5OGy7g37FjyeU0Zj9jrEDy9vV7FMQS3fi8eKTQM2OqDs5riMho+ky3Hn
WlJgZ8X1oxRkLegwyJRceYrIZkD8NBGq7TSNC12zwTDc7lQn2TjPnmEn3ODhNf3Xxg+AFwFjGvzP
9MQEd6o6NJ1AEO0tPmCzgUyFZ8Ep0Llo+SSAzHFN1I6BRcDkWU/+OOJPskNgBjCZkVKgxeE9Ltub
3qwuCCHFGYthQyxOjlme4AyHfUZeHjun9hGHamVue6Y2hSQlMhGhDMxWkegG3JqUvZMqXUMbT2vs
Ca9QyAbxVc9dICrDutYSP/kiVqQfjSvwp3ZE5GQOeGcMCoV2MTsmBPpmiN6TXRzzwp/MmwBC4tGL
Z1pqIHlRQnxGZ4u0mF8pZBq4UgE7vvrIJV5Bdlm9B69LApOzM2jKQK/CRXHhbLLxA77cTrX+kgae
q3b8hoHgmSNeAtihlV1GumIPJFAT2K/mRRLKeiKXLGJxHrOTD19Kc4msWm8uAJvuUcRz6Q4vssV/
X4G7kIIczVMhfzQKUcMrAku4aJTtQDbeVxI6TOZAz+qO6YuBLBsezzpUR64kLTZ5dyFjr5NT5H2F
cODJ/x7BRhTh+zfB5Z/vWDhk7z6dOlmrWlsFrP9+l/fXi/g1ohiuRkfvrF+4aV1zs53OzOuCXswg
BSJ4pzemv7gZS01MHQPjJnrRDGy6MbrpLRtOvNFTxf4Ol+gFPzUH8jV/14CngYmaY5qqhMamCHrf
DLx2yYdf2UASeaqQ/iQOmmTPa8jZULHSFZ63g4CoomD1ehYqEPJyQczJxqT1GhFNwuqNeLEPac7v
DWwEBui/Z7oXk8fJIUdF6fl5l9Zm/jQwTi6UJQqHIFJLwX6SEBD6uVS5sMLTLlKj9KQzOcU3sUrE
HaqTy72aa8+1B2PQDvyechAy4DUDrLGkceoRoCAlpxc6vmcJRfkbQNhUr3Xnm/riigOlS9gbhL9J
5w5oc+/meXSTk87/+gBWAW+id4ndyH4EpSiVsY9q3bjmXspE/XMYqRTCNpQfANaoM5zpnL8+JpRq
A5Xk33MbPii/mD+TsSC8gWztXws7n5mLwIfBjw7vS1NVdo+hpQ7zLgQeGMIBS2wRi0lEtzB4b20W
Ls9X3csb/WvM5EScuxMyFZeKDhgz9l6qaOtYEqOrSeWl/6CLQ+gDwtRi0n78j38UEh6kOIzsxntW
ZdEIYlnIJ75quC8U8fJX1mI2YnxNGDT8CEzO8Hp4HP0o9X+T/ahmBPUEcKCkXleo8cc9XtHLrXCs
DwyMkrsQtPiiWQEKPPe7NXpwM4tR8Xy/iByS96xmwV2Lq2sQxRypoBwR+XD3siIJ+ZhfOlKyGhUm
RRPBQy7QWieAMFQydZELPhdHUH81zXVayhXSlcg7MMMGYJ+IOx4UekpP5z1cIxZLaoMlvp+woQ8+
XPHU1igehYarKP598ZNPbYuwdY8vABMmKyDfFpSGBSJQBBCGjy8CkvFUT4U74YvMBH99ZmJ1JS0T
+5siVnXJgk3DeGDVBYXCBfKXKPsMv/OF9VxZAnIwHosroP2z1fjwmO9TJk4hhT8x2PPko7JOWcjP
K8KIbHqU217+E5AtHewGGpo7v3BQ6VLUugAbYkzd/RLLatUj0tZtNVaicJ5wxhvehJ2n7feBG+cs
iJzHhbjMQgS/9zWEq3535FvwONmxdHeiYaehnRXQ7OguhEDZo9szKB6ILuK5UzlSRuxKYgME7ec7
TZdLzi9mQC+cMHqrCSbfYS4OCeN5bGpQFIT25t1nIazfpXJ1X8FGYKRdTDsr081HTqyAWl670oXv
nVsgw6PYIw5vzdSixUYooG16MugfpN0iINvr+ueEWGMqah1k4Xh6DZb+bLkC/w8Vs2xvV9wqTGLT
bX2z7/ftXwcQhKF6gZvzGJECIt9gnKJtOiNlY1QcwsbXsb6Gr3sGmY1NSRjjuF5X7htQdbFn1pXy
FqyCXN0IY8Q/AoVPN8N+w/3WMosSaEjkIXHZZk1kORcL7Mo/n7m8sI9F3pMaPkkqiH/ZgMRxFFbI
nW+sIezIWCEM9qY1GGRmbm07eher9dkt+NHZnjKsKW+2/CA6zWBI3GK9DRloBjrzxoz6PUp5WpOy
ORYMtuQcmkNaCoXlj7ZMf8ys3EdfRsxQ4awJ3L65pYDEkYj+jwlSijWO36pBAni9avlAbztea+0e
GAZlwTlmzaU4YixY+XwOgPMIXGlvHZ9q8Edes5QkfPTGt6BQadYMuYAacHosKkDnc2LxHuBYveAh
izWSCJNgABinX0m9gKw2L6EoHDXWjPlr4gy20r2N07Y7oudKLfH/eGYWMIdf6ZhpHcgT+oSVXAhL
iTbyN474eniQXGX3WiL2RP/YKd42eOJJM+4fvuQQgwhgiWcHdAdGaAGi/adHoGAgCa8IuXXLaR6S
Pt2WyY+bF1HhsbEf9VuDHV35aMowIsRTXWL7vU3NkKysazCHSzEMkBNICPcPuR4TfYzCvfqtuCIv
nI9lQlYgVbnYIJsbx5ZTuXI/kiG/UEaLbY9pUEaoqzjl3v3VIoAnwO+PcAcyXu7USIrrkkyUn0JJ
3eO5Q74j79NldmyDQXlU20/3MslZZvzZlpQQMJ3U00NWGzECpqfvrJmhCMhiELOgNju3b4Vi/Hjz
rIQOurYOimsWUeZsaZDFIFYjMpoAh1UpxCzyKdZBy4upFpI4oU/Ea6ymzsoEWlYVoLk6SBLP+FkR
5eHBQtIgefsh0clDgOVcK06tYg5Yj18x/HC7mnQQyMT3UmkwFOdd7a1ABZKt1EE6KXp0hUFRDz8k
cwxilTMxcdlDYE8ACCq6TtEcFaaVRoaG/TwggL5oN4GWnzjMmeC6xbtnCBDiL0IOpVbxzqFWr6X4
NeVmqXPFfTgUkN3fICkvd5cM1pZ/qLMaU2fJ8Bo7r/afLtfR0vVjMjACvazw2UFpGX35GbOVL53S
NdyjvRJFJfQKAfw0hM+zPYoEU2+YmGvzsxVk7HvHjic0a1a2opy1d731xbW7mLFR4W/Yr3PKAel9
1OPq+ixvevH/xuKsBVVZpQ/JKNrbxYxb32guDAlu3NI/PoJ8xal6oVB+QKumc03MYn2ZYf5NAn7B
3gGyvMUoCvu9tbUueYaHzaHt3YaL/VMtI6FT5UZKisJighsoFE0jJIzUvK1t9YVVr7w9upjeXon7
CcKXRArXQ3QObIGpMoSXVmUA/oPxppUtM9n+Hjr64Vze5/RlBezDC9xfpIfSHWV2KPiYWtwvwxXd
bA1fJFtLvSxhHOMprGQOuaedFBL+VBKShGkNm7COvEpIp4Pfm9IbejuLN0gv7iftzP4RXcG8IPKb
UNCVEQNM8RRaHmNRIKdPyZMfGG2oPOhzGVypQXsANXrJJ2IUhKFL5xmOlRvG24jW4I0Y8UvncW65
RUDVxg/k3enXruhF5uYSew7LNP05doi8+ldo5OrplzDQHMuEYPK0h/AmZzMlVZoM5wGPspw+UXhw
7xvQXDeN6IDkgb7tll6NSiEMN+fNSQFgA8/oE5MvEz7iVJe++ePb8VuXRKoCPxRMkaArsoIz+hGz
P3oXPQ1qA74iPByV+U2zCcJbnpaojk8uc+0O06flQh6W9k1JO1YE0MG/9M63kHnqeROYpt2+z9MT
gpMSsZ8v4JDzMfyrLgbqoo3HptZkIYXo2e7b8hNI7ugxnTO5ZW1Qh/Zp0gJKQUWez3TwWfV+q3C0
WlGLKOeKMlkjIR8TFHPKRUatPxWyYhd1qmSswFs0HZbbK7hw8KCBKA17iSg6VH4adl7XNfsNkBer
79xuLiEFLc3LhSKrqiTjgylZVQsxbYvoaxEMyhyruAmXfSc1FRlZQ4mT1ekZiNYKLDSJmhFYMBRT
jbN0k2OYOfeR46hAZRuCJ0XqmLk803rMDr30DD51Yvf+bOE1m12RuPkcCN0jLdKPR0WmeXUAJ3og
juxRTIqQ/bpMcqgi4qClawinrHmDdipqfHS3sfeGpMTIXpCvNs/kigDU5GHKEYAkSI5p8yfbUYaQ
A05bw8iY1fFjywihlm/11mI7UAqnTkIKHF1JibZpC+7E5fORgAtL24ugPXawA4IdKr2Jf7lQtlrC
ocvEw/rW0A9q4Pyef5uab116HYqrOEdcvAF+TKmGrxuKVMn8C5GBkD/JjDnPiILUoztTJCKistDO
Q2+tSLxFdYAsGzQKmorhOyqNOMr8jiGSGVLRXpk0ZRgs6WUbtiUUi3EYpHLL9kYWG+fAT4s6WPFt
zVA/oGJgsyjiUlwGfw28iOj0VMkKKoaZqeMlkjKJwLfe+xbYmTD5dxsO608H0Z+D59/wwNtB4ERz
Y1he0y3Mp0JQxirtyu2w4BuobWaUNtM+4VnAh8s/RxOyfOED4npjtFSYZJbtZor+ENofBVHPSc2p
PLH5wc36EChPYIw02PaniztgKPF8NN5+Zi7Y7om5yxyL59rMOT5baabynytySd6evjSI2W9xFYic
+bSTAV3wNJ2wYFhDDPWlRtvOausycHsae5Q/ZrBUTIjJX97e1tMC7Pnmf1m0FiujaO9HYNJTWXMZ
9NZzto5ypiZzse2SUeHpH27xkBeCX8w/VxibH609koM05V98BFl89sZNCTXNSnuTW8i/yKTGPwTA
iMTyHZOY8s9ajoaFfpaRFrHEkgp7Ce/2G9fgXqjgd9RlWCktR7C+AC/VBiBWpdNKySNTDUit0Igk
qqGRPaccjjc9RY9z/KlqxowGfUl7QblUv8izauBDODHpQTV1E4Pt00TJOG8uLMQsvXrDMBL8H2RO
W8CLPVRhNtkQQsvcrEhirAso8s7CykKiv08QV2vuKrH9sKjlXw2bU1QEHNYS0Hfv0oAai6sxpuHk
cZP46JUKwDYeXzWSZL6GlXHCGjatEOWcBXH0CgNPr8QYtFmmdURruIaRfjmJ2MYPWn8GrbRtARHo
AjUTSW3EfRpxq8zkS1zlX4/bGnqgARoBHHhvcJOxlXrbDv4NMZflwgI3dNW+ONfw3xqLiHeWHpt5
40XOIkjNxwpRBwoicfTJm3nD/XHT/JIP96aktbmkkuc2Tj2Sl+FIhObPWklHVh6W/9Egsft8OzCY
12J7EG24uMDCSRFAqvMMAo4ehtxaRQpBMYDsxlUkbb8cpArjNhiywdnEyyKK50d55vduAVigUz3l
CgxMxZiyUWURO3Mz1L6QHwmRIF5yY1tdBLsvHHrFF7fQ+phcowSnzKlBOlK5qMla5d469iiofFc4
znbpM4dmtp3SrchLFIU4ejyxzZIzUvG3k3u39IfCNQwYoQ3kq4n8FPTv6ZpkIOTkEUcLosfXTB3Z
qd8X4z4nV9VJKoACzhsWTwuf2Zxz3hQECTly00q/7sCEDSbAauErsnBnYwauf+6e0SEQolRcnii7
XYXVfXVxhVxshIB8MlVLmCeQmsJj1+jJgeOVGOsCd+VeZRTLIMPgaSZUIMuglOaOUGYUNpKy1KHh
oOnrQyoiFpIp6kRVgx7Of7ani1R3pxtizAHHDjLKnTs++tRfN26OrvQcAt9Tw9aMw7shcTI9MY1/
SrXQ3tdr/kf1uMEfsU+im8/x14UFx3b+2+m0wm3gf0bK6aUmKdzHqpJ3C2zn8s1qRLiELXC0xutM
ZOuBrDqoeQeBySSW1+dP6BdziMBiWVseEJ6XXb83hoYPOUc6qI++n0gTThu8GW/X8VpDSNrs8ZxT
DsQmhfP903IIuuwfzc3sNGmmIDNcX/2TnSWwN5Hi1I98iIzuPsi2dq6QO28gO5HJ2s2wIiz4UDGn
BPoNNcl6SOb3LSiXr5nG7VrwR72xOHwmctZ6OPEJwsII/da/duS8eP3OL3pwvbN0EenzHTp8ywfZ
3IfUIWRTf9BLGruXEnelG/B8HaiWYluHM/wOgpwDi7ebdNdjV/ebqMFQe2sAy9Rq0ja+d/gXqDGu
foac1FqVBHRuKFb/Rgtx1rnUZbo5/o10jBVw6EhQ7AnG7Wx8kdwjKhSitILcUc34zvE5O+JgGAxK
o1qbfQBFt5SuUsiIl2w2qaIA9hkhzNkaS+vnHIMiAbZB0XPf2o/I/eZLzl+ygG7FrbcgwCi6YMoU
mjCl9LcHt8KgCW+hKzfAMCNU4zAEg2MnW3IY4wLYK+qbSHiYUCluPpdd1MhFw1cEfPdHgZCm8sxs
x/LMCqfW9ZA4/XF043zTXXTftPiwnrq6p65CRH+AftfE4XK/FCNmXm/ls7KXnTg/+lNHa6tHo2tX
26+NZsY7ERM5rUPELCXhnEIHBRJJXNSneL6g76dFyDMIlQCY7fz3VZRHU2Ixm4+cezY5rvzW5CRM
sXe2SpXbvE6uPJ1SR4gnEjmy+nvJGE9zTnGmzHCeOkduazx1iADxN1GUOBqkUOgxWlKQ5YXqa2wa
Twrmmo6V/TP/ePCfqFTgFmZhRXqwPpzvlgmKVJqqyVV3u6YJw6/bm/t7vOdJEG4qkk0KAeqAGOvS
2hvWsKRI9FLm4EMWmgaayD79EvcQkoGx3AwSyfXN+W7tJhlrqOuauFA8Q6FgxwjYO9hiFw4J3i4X
i2VNEoThPZ+u3HUWFTvbSDw++E2rA0Uj8WdR+6XMtzC4+mjDVtiorNfCHQhbfUBhNTv2anf8nCtE
7dFAHVyom2PoE4CWR7/ZkIryiUwhUhduI4s0eW0hV2xdzqwEJd+JDAOd2aOp9ftZa3ga94YHDd1i
uq9JDD/9BDujRqN1pAAqaY1TiuO9aqeHtIKYvXmkTKCBLKkVx5ZSS8ni2vSR1LTHtF2Pe0yK0YBt
nN9OvR67GD4Hb/c4a159Oj0X9Hr5b70YQPcOLg9182/UXEm5d8q4UCFxsOTk3RciOhf4kAst0Cx9
Yp0JpXFz5f8+acvXMlAhC6T0Vjc5XA1UjeTplUDZ3msceD92CnjuyRBRNildfr75im8VOxBnPIu0
wW5k7Oold7DiD+Bc0tPDubAsKytRXOXi46cMFnttWbY4WUKPoHEk6VwcxrFIVxQ9R07VLlttH8YN
DFMMrySy6XyhNKdZ+61QY/ss1b+rGpJXYsykrTpioONTCn7oYX7yN9rdPP+/JNvojZmTWI1KBWqj
kve1iNZiUTwVYbp0wOxQ+HqehtSywEV/J7HGUQVYJNTmiG9qt59jInMf9vb2uYfZkH7AWNIG+9UL
e4TPxrbRxRU/5DXpjFfdJiZIBr0XNwqw8cCGDBIh+tVOzm3Ud0sHpmYZxf59zjPBXTo/bs2JATEn
7uoHqd57eN9B5vYJDjtaAMIfzfQst5MVD0y/pqnCl2hkPTpZcv3rVdZ5N2QNXoEqIxQbD9FnRjCf
endk8F2OzymrLbVRaX5U5OMcEo0dk98sI4gw00j5neXWijYMsMXGVkvnPThF39++ZvLkZXNEu0za
jkmwizdsJgLPoxcMk8ZY4nhCp+5mqPjjPZum0shQeTmJTnzwdNHcprvTerfIeOLe1hPEpnkmEAxQ
9zkk7a7YW3PwXhQBdNG8yJmHA8E5vdCyiJII8QtgYvlFVYoti9q8jwLFImbvbvcvuvlTBoM5DcSh
gfpH+6tz7oXTKysd7r/Zn1BIOAqvCbhbm3sltcSLfOCvMlFEpAjGXkKOceHAqBZ60AY6GofTpKGQ
imb5zVoHFjegUriktHYI9pob/z66r4BRT29u+rRw3jgCyu4RS4oOvKRK7qQW+EgPw5f8uL1sqW6z
Af0VtYN3Aaa5vkaDYEJQsWB3EGVrnsWW4aB0gboRrqzHN5TRvjVaMsI09xvM2LR4pYqqOcz85ld1
DpxrahF6rWNfqW0YLLDKLYwQfocjHEWRjUEK376esP/+m3vbDg4KuuiDuXb8ZUMDiyJt5K3HATyB
K9UAUhqbGwJzMNBgsaQr6c+WgL2VaW6ToYl92eYAay84YpwYGiDM4M1k+RkacvLtw/1tFyi9+gFt
MMXeJ2vhCjiLSFm98N/37dn2f8TDt4nfRah3DtItbGE/dpKd9jBUugNfSXU+AXRH4k5MHcDH5fnX
KfNNsP3EWHZZN/i9GLIObycmh/IBb7oB8zR3xQKj4ZDCAtJ/Mls5+S/C8r4Z9dgAb8YjkHP6VKDa
b3oITiSWRX8ByzmS4lzsC7mUl3+5U3HcL3jimG1YLxZc0NPKxVAVJqh1G3NvZSYa3JoOhtwCG1Rs
Rr4SflH8VSZnJOoVHPJdrakivzpPzyhIVNbi1bcaJslT80tem4gW3p91Df1CUmtPubAlMrJFtZNq
64aVMRWdwszwMgkNdCiF3l+LGQv8aDzr+MvfdETw2AdRpVbXNLfGCoaRVKG247txqWeBjNFBE2pD
nKd94XKkOW+otD07+316moLUvVIw4DGaqdllwAdfgfGmhSkw4WHPZGEwVNFHK81tFIoPEcE3QmxK
4etNTpkGjQocnMQlcKusbqBtqkSvxa18vu8wu5X5xyuYKwkLZ2NeGTBDVZ1aqifGSj+Zo5CYZWEr
hzv7ymfGt5/V7Hzro/0mQRj4bAs14mSuX1qAyaX4KxemcQJ7Ov16p/sYLNcW5e2RPVkgW85S+S7U
Q8oRTc7Jp48HuIn1OhFre+hAMx8SJH4O51g7h5K6wLHo49DroYX5WxmevZfFM5EKOAfstSNLY3v1
JN0wAIxxxZiojYH2GiPVXs5Vwr06Af2YXqBh7fiLla38nwxoZgjt6EdGEXXljpvWcsAj5R1WWwti
lOmLPajoJfUOGAQx23fOeiRFi+ad8jcypTnFH2bl6ZchXuWM99PMUGYf5NDEd43eV4NIXjNzwxyM
7vWihJCrYPTWRty2ONQIMDp+Mm8RV48pFYkpSSJvIMOQoLQqITo6MEKYenlKcu55062faOIgDB/x
pcFcEzD36c0ijuF9DDSQ7jDDg9I53N2aBAB89AYRgJQ9pNaOZPGnGFoKZqHbqgPL7xhXpSr9Nq2h
od74jeJK9hhGppyJFIJ5SQZmQxUwfwR/DxJEySEWdueboUPzYjEavtBQ4CkH3G2bCipRYZMLo03T
xrvki/SRCLT7mdrovOTO9wS4YRkZuSAyMWf5yWeGmUo0t/4sdjgZ7NCrwQpIbYIiJOzJORWX3W+J
LKuZwMlNcOBTkOwYDwBP1sk8QOVG4HtTKiYoz0Cg6qLd+fUeC9Z7EY4yKHiu7GIIjHtsOgIXrdof
Y6w1p+VxXDyBnuGNzD4UarEFqXImCksFhiw4a6LK+SzZmac2cuTExsDlFoCbb9katIKWlBnSZd4V
5+By6fpVrrNW4MULkw9uy9aXZQ1TfSAeAMz6zbVp3rFJgGxwGe+YIlABA4s1Xus8Bn+qZC04gVXr
jBRzA9CdCc4uwGz84/YAfGXk3eI/9s2FVILS0shTgeF4MKj5dDSxLwnSQ0tJl0tLInU++lzPjmGP
v5KdOTmKCz2xYdUxP7KVGAIG7EsxfLViDTL1A4hS3OPKqLeMIosasaCPaJRQHQeyX4Qj+q8utLMC
En6RvC9mxFKfBYwbWhA3rXF8EVPo5TjOkaC+X3yb9Mx7oEzjldEcmRfcIwXYG7ZBqffTkU+2AVY/
nVcizdbDrdbXnEquuSKLWK5oOoUeFdAmWTjgmPMKOn3toVlJfpx8NrmyzdBNtBljmyclwOYY2qQc
iPpMss7CrF5bAMDwacIw6Hsqrd9z4dbI40jpveFRGkaHzwsSKa0Qzo4/OOJEvkG52eMs7tiItVDm
myj/8oVpzQjqMOwPE/LxeMe3lwx/rETdGMQvK93Y5x51w9Y6PvN18PDhUBz4zfH/gGSFj6J4EuZ/
8RvOZvdRHczwumSrmHqNaYpnlET43xRUSP3sA5kZTZFCWj8vuPTiXkDqc4RZRv2ti91JfHqcssGm
WiEi8og40gXVDRPCDHST68I7qzc7+5evQLm3MpSZ+UWRb3Dp3yYYpyvbzpThMPDHutNK4QlRRQih
D3nXswj9wpQwHKwbTl+9OmKTpMUr8OP7ey/xY8DG/X1zrIgXx+WuFlaVEM0bJFuY1aaIxVwNd54F
wJCdK8UbeSMKT1fvJvHA/hLK7lDheNIKOPX1vBHSRkxSdgoliYjXz1TEg+rBdLUQaIKfGL0wnwaM
ifP/VNlGfJKii1PLJr+jx6Saqza7ZSniEwOa2LURE+J/VfPrgTEvNd86RzLG1nhYs3RZcZQYhJID
1z+fvgh9mBYWE9thIk1nawYzjBzeHx3vnm8aYtv9X9oL7rHrq2L0pKFPD2VKwk8I0acZJechPIkv
IuYiQzwIglwxFK8SFaaTu+0uWIrGNXgdEA3j2Z+YILVLUchHawndDTxnQooSymtit8nJBV8Y2Bzb
nTca6FQNprsnJR1vG5pvLbxVTMgLbBH7kXBNIzfocF5nC1nrvi4St8IWc5s8E3m5p3BdWfVdguhm
wKJgQu9diknPBenEchbNQs8oYe1YK5ti0eX9sRfHip63ucgsPrthKy/NLtQkM2wxq+qtivUbMnGd
0Kz0WSLeYVi9T9oyMAx4rqKTXiaz7NJyrVXlnnjEY4FXQ7uegVy/Ajpgx1aSHlK4Ea6VrHCeWlBY
Ky5qJyC153EeliWr2KON5hsOil+HLxiH7Wnx0jNoV+4h4QsT5OlEJb9l1vDeWYFpvCV7A5fBtIgx
a4gjo1X0qGVAD1MW4Uj+FNwrcFB9VLEYZrwP5ZUu4jTagM21Gb9DlqmJZWYzBPDDmuhASsC0nCVz
1Ksy1tKuKQRGE9XtCrKtYZedjSVAtvXWSkDTU0D9C0MI6S6cMVbGBGPnwzt7JKDnMNznPTPhjw5O
L/3qw0DEfayD25mBvnNJqVRr5DItwN8mMfx1q3dPNywcRy1doiit7YoxgFiJiiE4/VW+HH11tYlP
LvSQk6d9VJQO1d3Ao6Qwio9ZDcW+FBOk5NzpC8cHM+KwTY5/LAi9XmiaVQlrh2XMsTkqbFEfRiDR
6aHXYqbgocvbJ6txwEYbzLMBtA+mXaVmtEFWdFUvXoSCsvcjdlSXdCemutsPyP9xmSWGLmxP0Z6A
jUc3Jmnzb8eMnUooAE8GO93gH9nwabzapVEsqyEG2uC/QxupWFZVkUYPL8dXoW3WJbE5TJYUb5x4
owkaUb3/VJMlA569HzAK4MIF+f2s4i9f8W7dceK7zBl7Fg+gWV9vyrBSUBGuJ3Mfk1WiLklL5Cib
Dbe8eNruC8y3hkODA2LZVetCQZjZ0fNuKupfoKqoSenTs30rwvnt/aYHNdFi+/l/eWK8S8G7vkyS
zPLyk1exITBhckY5R1TnBIqevDP+MPiH42Ls0d3fgeHDdYO/r3S2LjzmTqMwUxdTUBW+GxtgiCed
Bh155ALXKUmDCYGxYRWC4mSJ76Dsj78LZ9RdAodMoDZkWGJcrtmF/Xs1Hg/427P8cft2ReLW5oAG
SJm/oWwzvdPQpE2cl9JhvT4dY+p41dkQ/4afSBF0WKwuOINnAfqTYqGTw7LDfMUfMOBDaUro9Z+7
Wq4E3tCeu0Ty3JW0Q2BC3oFcAcE39731inmqPZzciDvFz9ChNVfsK/SItHmdiOMPSXLOFhEX84be
DXJ39vf7niEquqprWUSsHHhFCKh07RYcvyr7Y2wV2c1pCrnEE9+YVqChkFRKi1x0gsS9QvWbd3NS
2Eh8uJyUitUrYx0zSeETyFOj0/iv74ww+uqFtORwNlmIxRdcCuJkdyiye1WXClmrp+PX0tKEVihr
xnmNrRLIFmelJ0Bg+uh1JwaW9MhlG6DJZ4YFeI3lr7VbCi+ewBphzDCIBwtnVo+YtvbLYd6ExU0c
2KDlxFPtesmfSacVIfCmp6CNGXbgYCrloA7IYz/eM81KSg0Ww58Sd2qTbDsvz5EN1E0gigi+p7g/
q3WfKjAq/j3/Wac2m9+VImawYbtJpcet19UyXsrC32zrwqr2Us/H2XQNsFcqzt5HeoxKVoARjzxE
wbnWT1NL3QqfF/TGsFfC0vWJKOlAI383dqXbr4saqzzJYs7EZsA/MGUNO957plodVZX1yTsgucNC
hLaGYRE8g6ozKy2Bts1yuKGrTh32PpbkulYc0GOv0Hmp9HcmysQEHXYDsg3Lazi0bRT+jJIHDYZq
DRR8nI6b0i4b2HovU3KrOG3GRSpjdK1NttX4UJD2IfVQRJpdfCRjyyodvJoOxLJ1R/faF43Vj+/4
FAWaWn3f9UjjU9jpVOvJ5BOIojl3C13ewUmWQD+zzGRQ9JR+2OvOhfZ7RHi3RuHt1Zyz3SFWCYO7
MhmhLoiCU6rdApNnxTKCAFTWQBCceiwJDJnVE/E7a5RYMS320U+OsqD0gfhFjgTX5+qJgA1bPeDR
Dakb3qSoKPXR+TTwQXW7DF5JKWhZRujdpbNTUdDTa95cerDtmgU3SV/m3Oh4lkKS1km1QVpYhSiO
/WzaLv3LDm3auJjcv3P5n1pc/IhKImnNVQtCKzx1AUMLBQ9N8aAWe9ctaBuTQTSI3F4PV9zzGE/l
kNdxP9tm7+V9EHxKTXj52mo6LLKHiPd05sE+N8PowFZUHqxLzJyWTJnRDABXdL5lVZBQj+SARd/x
W5wtXf0cEFiLpY6BgnXKATHOB7yRbF+t5WFLDXcpDxudmKsDQmWcWt3Qmwuw3ZVtTzr4BzQH+Esh
8aNNwRGzE+wK9ZMMcleJPY+PoWSS4a9kXwrxQAECgqRCO2w6aRWY1FDZych/HLco0E1lL004Laj2
0d6znKMnd4pAOvi3CjTLWfndsu45CI9icNmpDFG8hhhLxuLCzwkME44ja2fmTt1reQPGI+CPNzRA
IAY+ttmxh0WZs8BE7ngedoCqYbX4Wcw7N5fHrsWBN25un0Asl9Wj/3UvtAzL9ob0EbJ79Uu28B2O
LXCdqszW4oSodrrCT+76ZFutn6yNa30czJAwRJ6iCTAdbNfwxtX7n0ZjKl6LP5f3vgDH40RstEPv
dfR6ycO5tWwv9lF6IKJx/2ZtTZTQjky9fm/ceO7pVOojlThAGxwxDcVySoM1Q0jrCcRjT9prJHB8
ceqpJKxmbw01ODFFy2T+G72D90nc6oznWYHP4/g24cJDJhYjjgIMv/6FjEVmSfnLypOxuFYpJ54j
JwIGas+VokGdyx3jNUtkkS0gikjc8eNGD+4ZGdBh0+eqeapx/aU2DOYoZ92EQAw+SQILOuYHVQ76
nMyq9WVugp+hI97WckbjgS7vMfUTKzs4KtF39r+WgVhYb10Gt4dE1sVykFjhzC/87obWLUT9eW7V
4SP0AhXbPYeHctLElcqza4cFle0vDwqCxHORLn3/bKJpdQrii+RJnN7POKRucgv+4zuCc9I4G1ZH
SFcZ13RlYv37lAETz9To81iv/dRizk/jAcPUZzKoi9c/UQktBVRhXldbIFxPBQMyw0kpQ2SJ7GnM
0m/vnX3h2xnKy2GttbT1ebQlA22X7bIxobrl/jOvaTzAj7gSD7VaCtkoSnUADGbmuDxwaCcXO/e1
XmET8yk1/NpHMYqXIHrS+Y8BLFFKnHKuUGBJCLIj5DSwt1zXXYw7D4ICvhKeZvGaC4YB32yfagTa
VhmZv96AZXVpZygjiYWd/wIIepHVYe5SNYKYQ66w/ww7ortHhK6y6EzLLebFG3fKxwnUjaB61HjA
rMkz59yaRVLeulN4MNd021MtsHadiPySiN/7paLNtkdPwLWJ+h1Sgwchsj/WDXij103YcPcNzxzx
aVmjhaFT9BInak0zKeh1h31cUF/nkAU2+tj3kB4AUwPH3a+DQpqASh79CoA2WCfioKpIf1ku4Pg+
2bx+lW4CIFuYwu7+2eUYIcAxKMZfUqYDsPHPLvdjaW31plarxaaSyGkk46lgV/+8GLmNmlWO/V1q
pj2P5DKdz7Aa3iOi2+6q+clenVPGwgfkHXBE1cUlTtCmsliTPp3oyoi73yxs5aG5bmJ4zcPfQG3D
jwwZu+ezI5QBkZTx5gnWabIhYVoi+WMg4mfacFIsdozVc4VuigEoJf6/pHW1g/1hlrCk3gETG78Q
kh7ccyDn79DAPSC7LHXA8/mB43WW3xpGoDLh0yVog7o8b7KwUs2gux3mplJH2tsg99egS7HBwSKK
u6mv4E4NNxPAiSgIrq+NtFRa2A3qo6qlMW8s6GGb9cT56Y02HM/OEF+9g6R4GNh1mjsIaoQdIX+I
Q+cyMqGULvYbpo9oew0QFBJuFSFRKqWA2nLG5RUDokn/JTV9Ct6S56a+YQSZhPUd5AQhST70toLh
Q7hCqQgeHzOcsgb/i8YfUsrj/+ojTagDfxOXk5JABN3lnsC1DKpVrk5qtBcx1MjUCCnG+gejhzjq
VbTltnWg5++6X3DCtZ5sDCeF2xZqYBHYco0LS2bxUUXtE3KNMyGOvz4J29JmkYHKNCm5xZJtzZvV
jlMM3CE02tdOYkLoazXK8GeDrs29zMffTmUDcNOzehdW8ul5OjeX6Yhwuf11+zBbV+HpYM3hkY1S
uhtGcPNRz0BodfmWvObhvoWwq8xG8STnY/9HTzz0/NDyW2xxUVl6CMZBSIXsgUaNQMItxCWoxW+l
0/FuszMOyqld7kseKCT1kIR7uDzb8DmsTUM/7kV8SKlxJVfYV5qyhHphuZMw2PJLmbJ8nux55IYz
qgOiekmS2KP+FwvgUkjEYKbKAFO0o35O0ba2m0MHQnaK8jOwd9c468zSyoyqMjmHB+LDU/43uT2u
1IbALYl9toVu/XXewe0waBsiK3CHNhA7jiAE0FgM7grkB+o9qcaqA5ufcHpR7vDQ/jy1fPeYFNIC
ToH1/2GW5BLeIMIEbaiNq+AHG+PXGtL1LLMIQIpCoGhvnpPsPzsn567kSPrITI/PhYhFXalkdHI5
e0uH3+tbNXH+m57qkxCAY+rZdrfS+9GhwCYtovGLFZbsvAWWdwSCPtlzqtu+Ea9oC4+Fzbo0opb/
oLGPnYfUjgmpnCd2xgo4nWk/nNN/tcOuM9XNxj9gthUI8pmOiUs7cZo4sV7MBfY9GcTAv/SDEczX
CFcM+L8cfqwgEkEXlNtJvSJKM3o8s48JinD5JturjMcFQOvNq4d02GobxTVNqLkkf1FDjI3jh381
Rd66OuWl/Xg1xhFW/dBIHlneiV+ix9l8kMvj0B+gRQsP8I8MS0IeUaC1RBhDYAZpwM6gFUA9N5PK
MblEsg+svFjYLMIhzwtEI+4S6S9EiDAxJhbxDSsBcymsV7bKdYyIB9chEw4JaRg3dryCETzS4YsC
VH1qI2E5MDiJpGpGA9CtxHV5MGwmwhrCYH6N5P6lirs01gY8O0MyJFdZ3P+ZFL7pOrjCHCuXH/Eq
3c9EGMnnjRAPLeXmAtne5v/UEYUO7X2VVcRht5xYGepkBwER4TvzTuYG65ah7UdmXWL9/jlzVBRt
Nse7I9OezX6ugFpc3yXdXTVE3oODUNN43ixAXcRQlfODCOlzxblJeCk9ZeCtM6t+r0DYC3YapSYs
FmbogxOKRFWGldtQxoKaPKSErmBppWjOaZRONDRdIH2x09Kb85byEgIVjHhrcWFMqEqmn/ExRDRN
rLEyzYqVH1U8HDUOGNDsFRVopByXf2u+Tcu9+wblcy/ocnuS8IqJysBbrFVNm9Lm9bew9MCeo2Tv
WJq+dzMhQ+5PQl9nEqsY3nx3TfiTC5KS7ov7UipzkaWYiGyS1NZJxgY08abStE/FprpQ79B7KmgB
6b6w1D8kjN+ph0E+pQi+GfqgAQaCEq+81eR/UZywQIFjYwKVv5PjSTX36S+2vnuEzB8/e2GBudt3
wyq4TX11wRTlcJA5DAfJJMbJm7kIkKnBDlrqXFWzN/HXtBygqoi25L4SLPLOaffMiWFrxVXsawfQ
c1BH/y6n5+6QcbhG/C+83s1/WFhHe0W6k+x/rEbM+qNjb8iR08dmEpUAFx/Mka3pqenW4YBuIbhU
uoftAi5B5muTU4ZFwU4pvrXtTr+4d5aURLrtB5/QZr2Gzhd/ehUBvnotPji7X73sc8SxAyyk7r5T
BhxcvxZ9FEjzV/FoZZ8iM2p8qPV+FSpJ38LIoscw/z40qw9Bx4y+k04ed3XR/qgx+R0PkpWKX7FO
XgUw7x3IwF4Uz+++pL4/a+H4VKz/nG0bOKPwVquYjiL+CHY9LmVSUc5OiER5w6nDn++h5yiSqrzF
AZ3fBFLr3ErbU9vL5L/RgJ0mTyP6Y/prnkod9IeCWCM0MLl/Zni/3wONghfCS4k82BWswL6P4lLt
pydLh7OqhjxnzxUSH4iJQEaZrOYIJIZomIgzzkaIkqxDvVB6mXfETR1rq8HL9Jn0Waep0E2eLUnw
/UMTp6IYBZA/fqS0QGrJmU+8Ehe0gJsnAyJMU3zFeLnR1ktX2aBqM91vVIX1RSCTcs8FlPJlM2Ub
qGdxxpYaRaEIZSt8xINgnBJnhrRaV710vqtXqb5hzwN0x7h43tCjIFn+mRYqXX4CezvoLB5X8z0T
MZk56oIvXSsJUXpEJ0U1d796vceJGnr6daZJcm+IzTQ5QUwvgWHdWiQfhs63/rpqdKVQs359gn5C
yreirZzKs7YiIxr/J5C2hm6zP61IUaO4zO+wbIZ6J5h3rMwddFC2YCmMkN9h6jkElCpWHz7OImCO
tcOQbLc32qSpDY2PW6uv60Nyug5tIEyIbDzE/Fa6VU9p4OXcPBhFp9QX4AXekhqPpTQ5KtS3W74Y
ku5KqdbeOy+7SqUPi4dtGaUFrqo15C6lqBabG0v0wHJfoBvJcLIqxx/XdsJgCNPFKjeJaEuviprC
SWj6ZN0SAdaWO0SWvqdfwzY3DgiJ1O0EXuOdYhJslxPLCP7uqNVRREEoanv2OIldapOMQjSjHgWT
FK6S4cMUTZoaOpqP8fNm3B2ZQUiyB8s26c1GsG1llJZjL3BmlIKTIzwzVX8HIDFkpTLW21UX2rfJ
MHCoxYNshYeenjfQs5UNy3z4CjwyzzJbHfmvkbbHBaojaaP1zgXhlnnmVZm2lGXJiZbsmjAC9aLJ
YZaTjHGT8s8tGHydqe1LpjoypcdogzXg7QFZZKi1SkdqIvAeHuNVqlIZoXRY25qJUtVoG/fx1edo
45zY9qAtn7r5K7OSX9Y77+UNIfDpWS9LsdFmeL1hmvOQf4lArsyl5WL8KhS/dbn1PU79wBB6sybB
1piw+qSh22eLxzxbSTgz+ELMlEU6inEBe8vL/NX08u0ggvtJlfUk7bNJfbWtotNkDDBdZN6FXpJp
GTal9B/VUhNm+oa6C81qJx780nER7BePdZfhtk+SS+tlsrfavaa3J1/F05AZWVH+wtwxIjBcdm+f
wViua0PmQNSogUuOaFaasyHlBmwebHjgY+EIMI2yYKiNZFZKE2ISGjnNVtx34JtR/4r5fKJAlkoA
/Cn7hof4mMwiY2qMtef+iXBOm/ZmGKoQ9qwZPLE0CR/jlhgj0L0ik8A/LUa2nfa5BINYQXAAdr4Z
nPdoaW8Oq6XNDWxb882RORPNKbM3M6wrP7QhJlqhSv/dG7rYazC8XxjeK72omVMU9vKaJuvVV/Mv
YoZ5voYaSh+mfPPAqn+VXRLFHtInm7qRDxEzvajBY8qxLqLSRobV4d39mYpzJ7T0q/ZDxT+bTZUQ
sx5xRk8WcFcDfNH/xTYDX144jJ2WlrpdRiDWZC832/m0z/Gai0rZvGB5+45ey/LhkGJ2IMSVbKG3
2dVWOe+CBigRougvnNPh5BzOrr3dFk65VD07fdYKLACIeJOfBn6NazLQczTLM3V6HlgrYcuF0T5U
x1RKSgq3sX3qiYdx0PJB4ljC3XLO85tW4w7hzwMMUz4Ids3wCvd1WxKLDU7nOGczVqZ4pCTHbKrX
y7JNU/iRxeAqDe0GlZ4HkGwGz5fF/MavW/gQUlzG9kLNMoKxtAUNky3gyxC7lfOQjW1t/JslJdsS
OwGMIFBY1kWtE5MNitL63SqrgxJKf4WlNvxBHdKXe/UMRR+vseomtMg9cBuO3x9rAlcviX77Ulwc
k1OybgDoBQEZpntQBiskQsHlLMOQf8oawnjndjC2bE6fwnywFvwPfmK1HM8Xk5Vhyg2ba9RF0k8+
aUPpqy06pwjvtImxHnzdKnSSA4bqdwLDoUUq/Khr6q8QedujVjlrz7m+6zZWc4vd4yMObt1X3rap
LIOW9BzKw/OCRhx/dNbIFA4reTI/ZWaaFeu1UAJc/clyz+YvI4uQ8Pco5FPfOI9bA05xvjDHbfXj
O1L5Rq9p3tFJ/WsinD5PU+I2Y6/u67HFRu9DbyOik+PJDCJ5JQ8FJcovjWcL4DD6EbL/TcOm58NK
oIGWlS8uSxw+47fPnLUp9f2EGApF5Mw9QBLFn6q64fJQAakBZzTsFD22KovkMS+6eTARFPnhcLy9
s7MU6bqhGMKUabsvZqLE4BN844frqOa/HkpQP7vyVkRoVtgAu3SCf57qLEvJ29Yst99M5WIHUpzw
0QgW/Th8GQnMUXEEvu8QeP1qlE/QZOrvAQIhKtaPLGUfHE01GW35Y273duiSc8lpIcW5pG3zdVI+
EMMNrApepxCflcTSedil3p74V6DKTu3P+BwSzKWFsyULk/6KlFhBbs7X/jl5QnAuQtrzF1PyHokv
2j8THiyB/Yl6sVoj1YhzsSxk5YIyfYVgOiKDxBpI5JRtSK8O9qUkrDGaQ6UkG53SlfNA2PvyM+Sl
LqwRdVkpAkQQQJd4rqA/ymNcd5rGvJdllK1xxyhqSlb/Sy4UjxiEgiAMgO4RZanT7+vZg15Uf5tO
2Q8fhFL7hcTTUIQp98E5pt0LHxeXMVQ98siclkXZcTt5AMW+4Gf/uLryO52bmQsD8feRXSZGvW+m
MRdd2esA8zYSEf7iyhNEFdQa+pBYmfQuZOPwC9XVUcatLt5fSadAOYcA/MDRApaKdWz0SZsv+bAh
1E6/YjzNohCGdvym3QxJtpDDlz0R6+Q2OGIAftSdT8xuW8kpkBbjR10urOSlfM3w85hDnpbyk3yO
Rt7xEHuamMDpkSERT3+s1vKnuBl36E/PakEUA9Muy5rQMC0RGG40nOWJVF6GolpPYuMCCYjMoERS
Fl4If+UrMUMuINatMi0e2/BpbsbrSL3hBx7QMTS2ZzBcfVgmT/GmtZlmgrZ3Qy1Q3fEiWViH1J2X
acRP0ICRfEyNShBCxs4+K0HAGZ+xrPzKwDZQBdNKw3nFdB6n/VlwbQ9ffZAoqdj2A7UIJM+HD0PV
JlcpuPyzxGWWJoawzDHLFrUV2soao1CQF5ZFaU/hyiQc4gAs+tKKq/+H7rToBeMhzcChisTVf0gm
bmCJUumck4H3m9zNLeTGhxFpLXI+s0qrVl8NNFS7riRGTMLTPMTCJ4hgwhwsPJdQwY5KrIcqlpDd
5FqoLxJKCTCBaz1yuXoJOOYW3iUkKPtkUyAvZtDS6sg9W8brXbx7jOuQ3jVMWXqUtm38w5XnlJ16
kPrVSqRxE1udK4qltJfouM81iWYyo0rTV0em2d4ETuYBA7wnU7S+aq5dnNhcPQ/M1FrmOAac7tzr
ilmSsCbhfSrUG08azkEJs0dTg/p5FjNpLrWeSdXnqo91RpYJzVFolXXzQGE5ck9H6hfE7E+7XqAc
mhrnBK4aILJ4D6U7CB4wrtU8SDDXZ2xhugtKbLlNJVSmrMbYfAEc0vcNcWrrwweO47n0uPYHxUUN
pzUwXzFb5Q8FvHUu+Z2zhhG1YlIednpAFzPrUSFFOJMKgAOwaEre1RVenH4UymXXXbaNcHPjq/CD
vExI5xCIUtWKOFlVvQOmNLPZ/0vwqW0oXxTHCfP48BalRLOHINGa3mi/qa/G5Sdz4/ttVOXBqOl0
MW37RPchVRC1Dj/269VpVyFDRLPQeayIhZnKi0WlIHE1MpAkGzEhWHiDK74WyxyhEi0HnQgqUl1l
3hNOgSf+A6ehM31EunRJlQCv2c1Pf0RBU6ilumeQxmLC6HUmdcRC6ocAtW9gb/aAWVn9KLVhL0Me
7Fq1BcUhSQUIrvG6efqtYIvlrT/ZfPgwUvXASWdrQfX+9gNVT+JwmpRRk3vgoS87iLwwVW0eLili
oRfhlrqBpDaA/hRC+ctMNw9QIteX3M7UvIZsz9ZhczL5w6uwkDSFI6Z1YZmOiar/uMAmdSzMpegl
78431F/aNKDj4qwdK7r+vw5BrFlZsJG7a8f7EXFEhYTRYDlcbBt4dPTntYhDJah2VEqclb4O9WS4
TlCmwZJAfeez1Ca5/CDSqS9/2nvs3dWqp0FZIU2IDQBCcRNPrdRAgYntEWhFvKrhALFx40mTlTWd
5tt05ipdYZ7HsM9D75ppzZH5zzvo26L2Sm5DUZZhXw6asnrdQkFN3mVSkvroxpYdsRvLDSPmCvtH
WJSQ9QK3SVWB0yqg2NJ4apSn4+Cg7+SVjFdVb/NNd6cC5jsRzuBJeR3PuPdbUmilUpKe+wGaUz3k
JJ63ZTm6iTAsDlbgEsuf2K2QLJfA66X86T5Om6fZQ8jc4gw61Hv9Mdc1w4nFVCOIsqGEqwq4yuNx
Izm9C9PAe2hChCrwJx6VPwvRD6oXLwLZzd+z1x4nsnF5O/MQfSVCJJByWRx/DnPOeDKhsS+qLGxt
Cjf8NcEbRgFby2yQGNaSSuzZC+pxx0j7rtkDOXIgbUrc8o7IGjMtwVcrPeHxkLbFT2RVU3mjAWrQ
rhfqXx2dV8pXkMglIvDnSDPv/9+srfW+xRDAN9FxB3tWEwhNATUgayuBnsmP1pnW1cWh7fZt/BT6
49rORN8W6PZ30InN/cM6V0Dw6vLDSHV1TH8+LU94wXSMQaXsKpRVKnDLru8MQytvD4TB6m/4eLHW
128vkKKQ/8ZASI401gaJiOR5tObi1w15qdT/cKhpPXDLtoIfjfjZvhUMOShLSMbqvFbSZqLYBMkZ
UqmAwmDq/5ufZRCNUeq+zf5CvM5dCTiSWK2SZaoF9FJrt1NwP4oxL4+gus9SDnx65T6OO1ikLIYA
SYudM4twGUj+c3euo00d1iZMvJf1snHQ6LvX+W/RGCNC7CXWbuD/KtmDZX4en5eLA36XicRNp5W9
c5jqSSbeyVvJwli9OtKaQw2lhQyEWnVS5pwupJvoh3gbj7jV+pYipF+iPBi/8Nv3YUsiFx0mqR+Z
+DuXQhg7CebU6CDezBjNwbarO/1LTn3MqgxKEkqEzB6MbbE3lCkPppNfBKGVvIpRkwzieeTQZdmx
d79l1WxIHwlTQX/ZGcvXKmA0HrgWCjx69y/hKGD/VgnFI3JyzMDpcx0VI45v6JiBt8ObS6Cu5Jsr
kgWPqGotMFTTKLHYAg+9qO5g+FluN9LFVVKHUm8qfrAqQ72RCb/RCoYvaYjCn2cUq8Inhi9lRg/n
Dg/gH3aXcjdn1sRAV43K2MQmUeeXkkcXXgcBtyAbHh8fJXSlgfBE1G0POrWpyjMv8V8KuDG6NyBn
FTShqoI+PwO0w29BgVmvAOzpAKj2KX+MztCzFtSbjw6QLsrkB3aE6ckxlmwYpd/Mfm0RMqD9ISjr
sBsHDH7fNj0ZX8o6S8x2wARpNhMTnUjq8+SeTt/2dMtWTRCTuHtce+Mbli++bnYtfQu3/aizaSvK
SZGKc5Lz3o9xfSZiy6O0Lxmi2lZjRdcTdYX8GOgRddqNAss92q4K4Ht4ammeq6XSvRoXJnXnOQ8r
NEj5rhxWXxeU+pOnf7jbKDRoEEA3LNhX4PQtzKryrtY7kSM6xvxsN72kChF0niCXwOl4/QWDg+3l
I+2MrxX/dBwTBptMjOAKkd9K9fPWc6OU6f5d98R2l+/kmVInOMYAietfwkJ5TO9V0Bux/ITf5ram
jzSzXi48eDqM0+gj3NGXo/hmlubDhuqrI9p074X0dIxA4ybjfxofpDyqv3Rh8/bZrsdkbvKvGNIE
5xzCiK9D+EElhdEKLKcTFrUe7CjkgGVd5nQXrDlHZGpNS3sfiJJpClshHileB8GbiFliAkO6puFY
7UAk4/CTG6F7GXAfuYgthdJ8cMdZ5ZLSVPUKYMLcsuMqI9mzAT0pT8AlihaZPXGGggd5FyVyLr6Z
/aB5kRTbAJjXwbWmXwIQGpl1ejFiW32df7cjkFiQ7n0D403K5Y0OPi1gQmX+GsFlnTorVocCGjRr
1L/QJ7sUBNaRINBoevQEgJm0+9cmlwLh/mgMMoG6AjOQMo2HKWHHI6P3exrbkb8gvRUwL5Zm8OW0
FPCFapnyTggiwxYcrLrW/zKNU5nOj+xruLk5eaWiR4ziqQCpTdhczW6e0QXo1GOpog26X9XC3twV
fm6guPzsb06dhBMl1uC5AEyOpUc2jBOongM20RJ693Jb72wsE5H2E4xXr2BGw07s55+BNVa+qNNV
A5kagQQKrR9q8UlpGDXdg5YCKryYUubdMNnN8w06hQPnLKb3diBWvcaGOVMR+O8mkBIpZPR5Ud7d
8HH7aLPa2grIHeB763q27jUXx4e/7EUThGZLDvKO+HVwl84rsEceaEnTZreypa2b3ox+DCbIhl1X
nEkUxcYErYltVj1fDkW/xiMticNMnMF9bCIwx4h+7of+XvBDHWCpeprc+7V9REqOgnEmIjdVvV27
MFPnFt9YYxbFF8YzDw99eSiRL5slYCzQ/ufpz/o2QGipsbg8iOxOc8I4DI6soDrXqOqOvItMgiyb
J+hizTV3B/sLSmJri7HKlqpUhybUJMfjII1Mfjkxh/mj5g+2Zp8Yzud8BQ31jR69xYV9Lwzt0JA4
dmu70TYEk/iCNsIgNCN+NpskX9sDQZ/CdqzO5VwB6HC+q7gT8fLZRqBOQUHzWTqH/jtPJNYBppDB
VgJrbeTFMZNNtpVMvoAN8hof5obs4aPUlNWuBgPi+Ui5h536ECsRkZDQNzWwlqGiYXMsJrit8EKF
zDE6ZIySX4mAPiONuKEiDMqrxemqCO99A2xUzIBAob3hhRngeDSzJTvd96mnBIhW6Kn+uOS59Akg
4BOqHGEw8RtSqzd7Se1zLnAESKW7QllXDCWqyJQClYHb0HVpdnT0j3utfjjaPl93QkuPTenX3AxI
XR+MNqZ5P/EixkFvO7qN9KTJeBC5CRWJLG1ESCJwHuj71JoMRtf6EvsJyhDJlRyCvgw0WAD7FVrQ
5eQZEqM/qo2JFqjTO5fx15LWYsLlqfvTGwmzs5YTXy+Y5uX74cUNzW5hR7S7Q/PHNPQPLkdVOlm1
QCwKkfkKu8K/Thd1Sh3/0/tWtYQrmAY+prtiiDzmig3ER2syK3slzN1BHsf7qQ0kUyE4j2/La7uX
u2635OMzaIcEa9CElUrvSH284lAVbQI9sswtGI9ZB5S5zpEP6T6Q9qP9vDI3/4KX7LZEdyGjqAxM
GqVm2YieobZrTZOQGlUWHkoU55TTzhN/qvOMq54BVFRDYGbLDYUhpovQ92WkDmssffYbBnbqs8ch
wiWP6tIBeg6jqK9jOtj94iwSmrySpioQPPW7CTAaZzqS7Q9dab/4PD5ADEteKRJOgIWgwLqu2jiT
gSua6jE8b9DAmJIlocJL2I8NTZmtY5r2fqSaI1xjURs1rJ1VAbLv7zWYCJfu8UGB/9X/al7emCcD
E2xWzXJ1iOaOUdGNGAMVDmerF1z3bc2TsIf8gRjNU3AsBUhglW05NMLZCV68bVymUnoIQmCZ/nYN
E0I14SqvxkPysHbjYGxk3S6Bozxgnea38SPIPAkyYpLw/FTYx0NGFmNXBBhTJWMvMxzSYi8kN4o7
tlgpCOyIm+7qYddP2mIIVyK7LrjoyqVbBY+aYg8B0zl5YJ1HEpzDakRfupcwnjIM9gDABdQJKJcs
pQl05kI5SsJx7I0XiuWa61V+zAsj2RQ7cB1Lw1aIkSU6fLM5aS0BlBHWpwB8Sun7qJm2ZDzKuTXf
d3Vffgmlp+yf4dX/+0YqGiNS/v/0gwMLTSDLFlp4QgBeCMBrt11XtlPfUAYzjwX9CGCpBfRln8K/
yKzJr360HebpOphBt8HiQ59pNlHXD75aNGQbf2ORq6ZpKS0wgKyJoKV7Nli2KP8i74abPcEudoUy
Trq0DVTq51XLoy/Q0a3M7CoZz25Pm4Yo9UT1smpmr/q07r1ioHhy36TlSaio88UFQQjFAY1BApb6
wmahapW08sTnQP+wh/fZx2I1e6uGHF2q+cNlYD5PrKovPKSgPCDyaH4lama/pflxFfCZCkERyzjD
gboY6nh/wjnnxfYKMjis1GwGImtmEzx0BSiO5I+aRlNrrHMnSJo/7XsdXEOLL2EUgCO/wDOWWJiq
rhlgrXFfW1w84xGvahVBecwuuqZNSsWg4GsnqNSaTBPNvv7h8DNlaiKEkS7+AFs9g/lDyoovJxkM
T3bPlsNmLLPGgDcunxwq+9urQRaZn8kpsSWTh0+i3Ss+xZzOsZCuSLjpdz8UjO5oliDi1x9J1ACO
wkMWoE4sCUSJQH5yPoe3dmPTGaAglZuBAMrRDfY7OI3TID2ipAwHwhqZZRr0B/1NU6PCYkCAOWsN
EcSBqf7c3jtvK3dnIVSNqRXgqa9bI30+VLgpfjT15yNMMC0sfxHWrvcPeOtXtj3ECXVJyxhmOZrV
cSg3G3YYcEbZECgOynjrri+NyzuJ452cQDU9WdqFWqtyCqYar4eHh1pd2O5e11FRx0XRME92LS0r
NQhaCQaCuq0Fe4zXBOWw0o6yGwIAHdxsS5lxAwdNvMAAhl5NkwnbOzOhHEiIjXuMxXcObrxM5RMY
BYyqzd2v9vcLMlYb8CwjpfTQNtpMkGt7KO8kwfxYzsPp6OGXMgkotHUGDq7ikhJbT/iqIF/wdij3
WPagibldKNbs7UFSka53QCMu2AkNkgLgRMUh/pwp8Cs5GOkvAK958dz0JytL34SlBmNx073YYYYU
xVmudUXNPaS1ZD9sJpx8+9Beg2d1PxgjYpwLtCF+mxvfxP+xd4qS+DP1KgXcAYGJ+bB2IQ8vRaSn
8pggaG0Qj7UMP6tmZDNVoLmYlWZFhE3GwGUVgwbS0CwuesugLbGWMnQkG19p7xBqkks0OtNrbPLa
ye5fayLlSftYHxov2ofNUlqDHEUq1k8sK0RIaCO9yFZ0/Pz/3gQftRb0RMQ+CU1I3TBDhcnu/twM
SxcIywVCazvVL7XY2V7gJKn86mlNNkCcvzYf5DbVyS4meuzedAZ4K9zHm7h47vP7e9n1YPBJnxQH
Bd4Ya+p5OrC1yNPI6FmBnDst6fvBSs4PHe9G4fjXUTyO8xcSqmGF9qbPMZImJHwgXS62wijiGdhl
eux5KZOClep7zsGiGOp499O6Gmt9zWTsPbSioFSySWfmLTDWurecZ1opJcLEe8YGSlaPXzfK71s8
yTf0rgiemGQNc+LR3E0ie+yXYaG5bZpPydI2DlV8ER1FSB+3Oxm9eGxC0L//J16Jsv2fZvn1yeYO
jZrZfPQyMDZSLigxz9iC6oixidjEsgBBkFxHSDMBmgxnpgixh/7U9mjD1K0t3eF3A+bcGd3pJvcw
Nbm9Oc5egCkkqFjiDipt8Ji1dbxuwRapYSoKFqPRCm6wejE20D3P87W2k+bNwe5I/4NWBDIOvgne
GaZSIVstyi0zDFfbWQvcH5jq8fj4usPuaeexDOOlWaW8rNnM0GDjZbKJ3Fl7g9mw7cLW9OrYOJbV
iny/H7bf8Q2srvoX1xdNCfKsxXUFv5LKPEUjIPw415uh/0tWHjxyaZXutNp/wPUyX/Z4sFaWAASb
WSoveU/D+PRATXzST+dAdxDXnCHxOF0vQrZYihNpuFxgaQurdCxxOrFOMY7MrQKhHh7RZDejc67o
7lXGoK3alyrRdIQvMOvMfARkgsYt3CwK0X986O5PxaGPF0L/csbsS/rp6wd5/y0vPPzNQHFvB4W5
Je1SpDFhHBwjIMwp71eziIVy2nU8v6SK+c/LMy2AwDw53S8NV3hMUL82EotS6gecIPONLaUmgZ1r
laGE78A1p5ipBkQaHaM/JGywyLhy6shE06HO845HqkunSVAZZtPYQAay64+a0jM1Ia09bZrYCSyO
LJMIEfyqQVzyDVMOp1nkprPirnyMf0C6A2tPt73CdfJy7CWU1AzLz2ZzAFfGh/CDzT36dqIeLcd/
pv5zT6He3ZH7tuT66OeQkjEEg/i30e2J/n/N93yiRUwl9LVNl9nzzMtiAl5Z9+KdVsHvGZX3h93+
HF/qxtC6cIeHLCYteVxVEREIbPxR1yMY5DQFWvpvV6ouQvGTMtjxxIO9Ztf0hwU9fevddA53c7ns
+hjWjClAcNIQQz5LW0mJzkdbWTEQi/ottDL6whPpUtSVjtMSag4BWv8hAlep8ZDVAwhwl3+buPy+
RAU4gkAo4usVEwhHYM7JxBd1VUwpUvaQhqLsc8OxWmuwwkdbcOrG05aBxeNj3MlhKg2g0xxooH0P
3pu14RCnPDirMw1IvhwApRiZ0yQhdGPu0TrnuNr22qCPvnjz3PE+HfqmIXVcQX38+GZg7GYr5jgB
4mYSb8WbPeOKcUQG81JIDqkb0Tbib+z8/k6r3EHUF/v8hNDj/p2C2ST/e3FkuM6+A8pUEUXS0URp
bAuCLZaQp4IY8dl/icrDeGkf/pzEUh5TRt6H99Ljxl3m66rWLHS9aSod5T8YJb+CIg10eQi49TQt
BO2evT9nt9AZb2tzsdQUgw5168K9VFftwHrs7E1huimS9eRYScgiGA0l2wDjBxxLTnfl6uynr9rm
qY0oQhbBaymyH/adgcwftb36d4/jZzLW6rFpAjHpnGHl6rKJL19UcTAtJ8y9Prr1Qn8RPUTYssc5
AhmPf4uf3W20LdoJ2q7bjF+ZVW+4Pa7aYI+SYYtuOuxMMjBZz5sCB+KesJ/u+eoAz5NQZvvk9WPh
qean8QL9/pg5/v9BPP8XHh7nL55Q6oKTXNOtJtn//Kdkn1EKOmalxZf5os1sODv6yO9izOYQbErv
MSxFHr41PyFQmg0tifxXvCjdBGLIys+PqKAzRsdx3KGUfYcAlsShY1tvC1PrBosj9V365svM103s
xch7Fd9IwGOdLAgdB0rb6/nKZkP7BmwGgmbz8nQjMFpHmwLirDYzpmFzS1LzI59E25tXgxtPYqyD
Eyi2fg6zGF4VbNik6KbQ/cw1qS7rIedcu3pvjqlu9KwMKu8s8dGcoDvrO9Ii0Fp6+kiSg8bxAUW0
7deBUBcrIY9dmw+JOz71+EalsztLaRTC+Lqk4W1yKwBnHsQMDphK/vqIlZ/NfTN6l3bzZoOwLdIN
if+t2d18tRQzrQ4emasLOePZbyIU2zVk/vOKgQzL9sMZsfOuOUFkDLJq0IPLl1W4LIJd9exc8Rlz
4aicOiXNIjeKUfgQtTAjmG+wT86FA5s+lX/BIkkgng6GdulyUrLDQ0Cibf10X8oG3eIASFhyE31Q
ndUhjC6QF6jDqmeVxpn7MjgN5f7npnlLghI307aXIlesMcsO7hcDg3KlUqz30QdQUzBgYzmBY2f2
n3XqYdiyvHu9I2ihNi7djqgi5kr6aXx17plu9+JPo3PQCNUzsd/O60i2qv9kpnzGHHAWfly3DcKJ
S+7C5pvMZ/iWsW6Hv9cBFL4ryq1WnpRWNGHQqbLYBaWv6iuo8Kb8lclNzM7zCWhbDKe80esTjuQC
BmqytXL7EBW2W1hae5CNNh8bgZOguKHNEwbAU+sjnQLFBOuCwIDIRyuKFweIMw4oN2r89oe2lpGd
PgUDwEPK14aveDrSRE86WcQMcxhtpAOTs5pasi67iUA0mvZPB9kJRuO7wWeImE+hCCFwSyYwEt0V
YKEzklXIVbNlTQGzO+KplF7Vp3dh97VJKNYQicqv8bMNg0414KU4FAVaPe3fwLwxRVNDjBMAfesa
EN0TwzdBM8rjLvpUhVjX7eNiCZalEVqrNDH/mi+ZFUhM1LXXm7aUhYSEylxNZvRMxBp2wVLh4Pwc
+6SwPwKTNAQhGPpEG8ZJ9YTIKaCH1LWvHssA7GEQdtKr1e3nQLPxGmqQJZETcH6uvrDDajj8pHYH
rD43HwwiMndeVWDschCZ8JcZe5FwFFUBTCU0yy/mVQJHxoJLzqyc9RHm1DIPHJDiR7Ex7SpluS87
+X2O+RqzOlUHNWLrUUrOiorPn8i/g5R3RISD4WtbR8les8fXL14adr956opgFSl42NCWyt3uiozI
cQAhW5xXz4DnUeRb0axz5M4I/06LpOukRsAFWUQMluBgDpAEnbt1jd4pMPcHVsqAy48BHaNTbR9j
ExDmk+BCeAjgf1XcYwY6iZi9r7B77nO8EMsraRIIUtx26aqmhqTNvamAZa5zr607zY+wvFRI3Wty
Q0zYf0b9xQYiqPfGulOxvGwKyExaPuXx0fQobGKrLiEjm228Eas9AjTrJMCw3Ow2s7hQZ8o0kUO/
MSYoum4pYi7doWETUPYasT4QuK8eF8dETTIqLYv5xV7dkLQ+Bj0z/3lxgT6ZidrTHlCg98CX/Z/W
yj99TPCogbif1vVBbU22hbV+iemvq0/Aqpo6HG+unZ7yLNw4Pp8hWJnU/0qTbBVsFNr/5m+3PQu5
rsA0TpCquvPb0Gu/4qtoiLORYQfE2kmPa5WMXqA50CjIsbk2ckbzdqKA7i2OBF/QtkzKtWIra67F
g69c0qdYX5WzvlfNUmZ17ifl26U12I9127b18A8Sp/w3Xii8oEPIXDfO7mAr8VBlz5YxDosW6FWo
TdgvqgKA/W/7V0xc+XYAAhNF1H1BVK/FIleCWTFQRa7amFc8LcBDZDiXntdHxShpS/EWilDkQM1C
xjB0AD2U5/0JYnjAE1UP2BwOUXBZDi7dpQX0sxfFIV7BZ9shEr1FrR7YZ37lib51LZ8hfSVZBgYg
37zl+CnshjjJK/x/BKj6aoft4V4VrnpOXbxT5IMu/GTp5agF4rz6CTh6SLCLa3ddQMZ9T8ohZrGj
8psy0N7OSmvGOpZz+m55GQG6QA9qMIf3SwmVrBpdNRINNKlAK2J0/wgXnJFHGpJmXKRQuAB7TBP6
6vaIf3jowDI9YHRhNWB5Rdk6iQHTWEWtMrLp+zhZntW+tzjRbwb4OgBghVw7rtNyuizfsOugUOvv
hY5irnc/nVxrhBwJ/4dMAgDeLfM+9v8Oj9+9uzhBgAGAinSWGRED23naX0RQxBVsFqR89jPdKeFp
TEXO1lE7Jo3rzZVr8TuzrM29yE2OB7FY1ntjhYKftc96bzS7xBPWkTjr+7k0Dk8zkj44n+O5b5bN
dYhlhoohzwmV6tOjYc6DR7WMj8pAdWa8rBqAGqD0dqw/JnH2AzMrTvuv0HQIijhTCM3hUgPvFfVW
s4B9FXjnk8eJiXqg2Q1hIa96ppgDDY/Cy9CchXQE7WlUkKpsZGwRBJvehcUGLH3cfFeUs1ICnLFt
xrlxYrHQi7ILcpmPZJCN2L5rfnJO5++M1BY4fpkc4fWjqfL9kGlYmtZrMjqAiel49Ho3qXBA56LZ
hVhdmchPUz3cPcxzFq1bI6y3jfM1L2Z2TCB9nfvT3EeTMk85WSM84LtBQitG6Hb2pvexZdccmbn0
NHayXCsDaEVkdtX9NrX2cfLW84q9Z2H+BM5c15CJowAjD+o81iI+1+XMCT79dLY05Q10cj6B3RiT
hNUCssbdyLvWIRw9Q/bAEdQXI0dgXBoSEGhlqx/VqnUSHA3z5+CGzYdpeDvu9eY4DPXVOC/cpYFV
/NNzsrXrejIVJbGl+IHvLDBtTdLguK2MNBIuhwgXqe3f3QKmzYhoRtaUJEsmc+v621YWQOHpLOtI
USACllTlbj5ngpB/PIHJ5LR2hhd2KHXb7654mtiY03pxF0wFKGEd4DQWF0ypYozhBY7CbGqLaktt
Fjqji1Oimiz6xCcu4afMmlrAMCKW1iMkNzR7tLDIKGFDTQmnFGQFBgLP1EViv/QAbdlAWw6TY3VE
ubbYDb9SLK+kTTp32EYjIDQqWOuXn8mTFkLjh6SUD7/N2Wo/5D8+l9WZbJyHLipk0l9KNJPl1ZEc
rhGzFsPABBiiciaOquQ2+qhcyrMaou5wI5Ah+O+LhtXn46om6ZW7kUkseimTzHwMs6mWJGnrMT2R
JGeB83ImZfVjRbzzYBNO/xw3irC0/19ZkIVyRu+5hAIKY1uiiKkZ7bZy1DUMqsMeASIUX/GkH/LX
fhd+MYevfiVkO8KOfSd2rk/NyQsbjZzhX/fG/F3IJmV4K9TF6MsM5CiC1p5G6PFNR77D9lMmWUYR
52v4UXFA3uxPzW3+m999DCAILp+UpyJfZjQDSOQ6i4/gVj5lCrDiSoPJJE/SDN7wszo087ydkTZz
nYZ1IfABeaNG0K0wChjUFMrfQx2hqZm3WbpNogScq+5nxo3qnWsb6u3zIRun31lDgJt05/DpH8qF
Mz6NvIh4cC/0hFpSfWRNWLVRPWgJ6a6MMTk0iCBxAllSg5KScVWMZpwyUBg+FQbVsUFfAKtkxTY+
ChGdoZ/Edkc7B1Xv6C3ueDhTbxH4k1zUsYLn74h7Uze1WpjGEQUPs/F/8zUmDRVyed6jto5d18vc
GXTjmz5li2IyYZD5kicHBJJ02VqRwpOSPgMJFsgPGwrZOCJ4ocyHEmoWCqeDoxMPcoBJZ0f0tC/B
SGorU6/VbuQvHOfGo/amqHvSmdF77QPe/oxmJgrjWZaqcAhW5g/vJUqzyNiYAQW7aBUdUejQ0nuQ
OdDaMAc0mk8Z3rZ/yj2BaP/5tQDDo3DTSbK8kCVOYD3Iu87uSEpOghhDGKuIpRhQHuDWMKabAJEe
VRJJHAdJ1dl2UjK+r6rGF/9hLphClu6cOWfCpsii/SDgczYW1apSa0Eqz/rCDh7AIA8yWxKobqkR
BcBFSb6TAWuzO5WTFmE0xX/u+vshFx1xwRnlDa+rl8+yx1Csh1n+hl4f1gd/p9cK5U0XojLGt1Zb
+hJnpjzFMhEwQUoO0EOwFrDXXPMBWpZxrGul7TvaVJnVUIlN/+DaIiBlug44Xyj0keh6SKN+daF+
rAB19sq1p2zuQNAXr+1eX0w0I59CNuZn9UyTmRsPo/fS+quUmhoyqolNqhaugNC1ZLSp2BOEcYAj
kGSAuNGHaTn0ze/vx4A78dA2In7HO7H+STQqctcZMertBM+GOq7ql/lCH3lQXjeWIjgmIWMLRYIA
+RwWAGEDKk069cLS5P0x2fsevp467wg/KB+J7BfnS/s0tw/N7FYntNP3a98sY8ogyl6sevTQU/2Y
QTjYQ+5z9Fv6w6lEgevbE8zImaHTZSx4UI9/cddWQZyvrABIZHwP8DvGvqCsIYKwPnpsO22eImGO
2x5WuxESUfNLIS11vTDUBMr+XTP90jw9Ffs3Zzpl6kgQO0tX6/svOmm7dJwEpveAeDrQSzzNqpLo
3XCg03t5pI88tBLUERwK7Ag+1DezO3r9bsVgsZyCQGsk0zw9xBnvEy36En5jIAAbR+mKuYWqvOjO
AEo+y6JsKWswdH1uMSn5xPcC0jRksa4UG0EpGO8BhnPdxh5HB+EPePLIBxMkB9IAork7szG3WTrN
a1ZpGQM3Bu/0bMBR10QZyaUtTq6dHnbZWCfqbelvy2X5E7PNxKCpdKpziVABruEafq6nUayoWAGT
X4UCPqGFrDF6vEIeWDbhzomg2Es5WlqLNQ+uSDnrxaw8NoG+jHbbeEIQpC1MyevVNoPjdjusqxc/
uxjg3YasqkHiayGf3Je9NmXHJpPbi9y+JoDLXiSgxTONqwyP6rJ64oXhwOvXCAsXD1Gne9hS1toh
tl66eZ/ub3wJ9ynTiGqgPJkewSLU0C4tMQrX0vUajtY0tDCMnQyzP6TmF2kd/1InvD0trSCT1bOu
tufM/gj6fmUP5xwkkA1uUn398Gs3N6IdCDGYtgc1rJRAn7/h3BOgMBUCesa8zWUHA7JgCjsHuYTE
fXL8nJyp1fSItxQ2x/CD7X1peGzbZXPmtrIBzwBz4sezqGOHcyNxunEbOZnTqwIieE3ub/zcsXoB
rgBxvkPF9X2P+hAeq3S719Dzfcs3sf08NX0MKMCq7ZAv1XojW5l+2M8DTp4cgP3EP9IGDUZeVeCa
kXMlUtESIZKrsD3fZG4WNKnSQOqobgyQXpMcUGfjRA5jlTiVCTywoDbSB8JU9OXXwnn1YBQQD0Es
ftQqzcOWHXFuilWa8CmddXOi5KwwsWu1kpbeZi8Ad2wqZ9NcDK9LFK9fq/bDW29YmVPbf8AJHdTG
7z1v5/5m+RiHXKiYQnsD3L3K7ASLqG10TFqwXAHZU0hymn1VYYM+JW73wxd4ln+8LqnyB16yupGw
d9LA+PXKplQizucXQYoYpZBNuys5TraQixbQjPTmJuZ0rOytj9PBxEZdO4jFAf2dy2FGOdvXk4e0
HyUPI9gGVWqvfc9E/G1zzOAk0H35ObuIzJVgRBfKzQyhtBlw5eSFUTutCwR8zvQwlAODBaeJZj5D
3f39TeiKm2FRocz1lVp9NtErynawyEVgrJcx5SFBVL7hwebQmpQjurLtVufk5azMxfqH8GBQ4/8i
M1SinUoFl42y7+DhCHRmfbT8Z4VUGVl9faXxdw8oe/V7j6Ahyg2foC77JNPx3gMTgGt6alfog9Zm
kd8TMRLnO53jQnwWVVtyRVABRhkVy4yUQ6f2FFl3eAI7woVdVicGsrLsjayOhxD1e3AM/LTK7J8+
Ik5hlb9QCz4GGQgH21u6/idbatblmPp2Cv4QGneSMBVn7+zWyTQMFkGdJS7aFMRBRGB0/iLSQgVF
J+GqempkoCTnP5RCnIbFV1rdCrumfm2xX20T4LI43/6OupBnT+X5WiOV+w3x9+zSt7fldeftK9m5
zP7hd1MT5t3Mk/46DRuLLZfTtYjG+6S9BL+73nAH38enrrNSbZgpjyQfwWP7Bf3vILcMi1C9Ojmv
rGP5b4yDpjVkeUtcnUTSjgWCB7A6sJQBqHvnnQ9id7Lg/14RAwFZl/Gfdr4vqvED7SKrJnHngDUX
gvpy2ok2V5AXdzi5Hy+ou/Bjsy89fVZhzBL+PyHRqIZDSrk08OF+QkbpUWuCUkvft3TOJ/a1Pypk
DE2Vl6WDQogLiOSTtHsYgsQhDIA+tGiXs/09xylqqphTVRNkOcMMsWmmpNNThjN5+YLHV9kD2kqk
uK5bYtm8JEZ+f8UithMCq32BZAWYxQCWWMyds5Drtpuo7LLSlfz92pwDT+Pwyq2sNibJ6Cbd8bY4
MWHJYeAt95Wa7EhXTWYkA1cFlRU2nvLYrfIht33jQTbUjLnOzRfd6mhWwlGUmkQBeVO3GncgZrhL
aB8eSxXwwN/urtyPImXh/Y3xzj6JGBuabIskItNXsI94oilRuSB6GJtoruNGasbkilpD7ZQ4Ntvb
V9PYRB5cuhKqBOMUBqkyMzn+GP1/S+p1Fhq7/phfuXdNAy0QVE/FQ/MOPOd834h0rPmAYQJQK/QD
Q1Jju5GouPJx/m29XGBHp/Is6hlZ5FSfjLHy8uU7l2mYgzxUVQXsqzkgJ0itNmE7w8HbwwyTYAGx
Lvyz9kDTo29XsbHvcY/yAZXyQVSqeT2rD9rDEjdcFkjLDYssxlW2IJ6QGVwGi32U66Ga7p1VI4rt
no6HeRXo72wK7g11UtB9DyzecPPxUYzmoSOXWLPBJGw2W5ut1laHQos5zv8xHCsHjDzhIycjr+tn
gZ7eezqXXCLTODrIuWlUFrQCCNfKIJwgbDjQ0t0rWKsd3m7lKxOa2GWHanBL0Igx2WQQuMBQNgRN
r4zxnwpE3kQnL4aduL0EQTEgkLx1A9vKXXbq80WnPF8Izjjq6FTCUscOTB0kCkIm0J3n7r8Vtk8l
l5OlxhrMwczjqWdNr7eNxyImx0l6lQLhEdN8Vv7RTQNvXwzGnfrLMjeBmmZkIgOJKXlliYvcdT2n
ZK3NDcQ2n+Sy/YucO45S/UnZMedOHCA7bOpyLYjDNL/GDNnVr/FCVxixqXvIklHk6mK4MLG72Vzb
lDahg0d86ZPTvoyo086WPCS2Yc/JbfwksrzUrcBLdiU3oEEO1wttmst7I4pT9LiRXmD/KfchUFNP
myeE+jIZ6HXMoqVM8/PzlbINeWwCOjfRI1ekjmlZECxxZl/1bFJMLia+DBb4oOMbUM2CDT9/YYJM
BJYuzHgKCqf9L4p8u1Ssyk7Tmby+A9NtHQGRi1LGi+jujUr6kmu+U2gEg+puOFJFXG09j+RI6tWj
M2loWuLYiFOHYG5ZKb/TG/qLu34TDv47vEmTrjigPi/kggpSEPFs9MS3Zgsxz4NbNXiiMfkrjkJG
ESTraJYd5AyZ8IabNZxT8JzrnvcB4M08PVLXiBEgX+TA62Ub9YPhZAJPqiJQW7yNuLJrhOOdXOPM
gUXeF1sV43tuG18EMYDaHWeYOgJ3Pg1mwCHi/fddQ2pwvj4jjfICwdNdLnmNkbewqplWf8MZ0Vvp
pqxyis5Pufv9kjAJcUrpK+LSvfSXJ7vRg1/heIvf2N18d4SljxxJh5jGkZgTrKc9/C3TXwptPrFw
M9+jXwm7Lg5UFl9ZoNbPxx/d2bRRUhHohvJ1CcP+YNyIDYGNVY+Fkl+XKvIj5yiVVJMErdKfbdbU
CRxLmaiXa479OtkimpwTs8kKfIvshSY0qb11LFpbBoPdjm83BbZF1M/0QVLfKgvwYi9xdj0GTWdU
QNLhRohMYdbMvgbeuWWHQYX1LcmqPhN6+QbuUKEWTnQ36E4T96k9m7JZLax+/1Ar0cmNFTuF/N2K
Wg+gXjmwOG6fuhu1CD2GllDGEasroNDNYFQmtyF6BXu/c7OxhqfUM2/lM74HoD34zrfcUyV2Xk+T
Ezh771HxsTM1fvgQqDjiVdJL84ps7a+iuJ+YjKnChdg5e6TXPecmQx/SYUBnud8Lo92uSOunkYEF
p2w6DXKqCghnH3/PpdcOskcbiI6bwKDViIXRpTO1ZIxsP1+A3x9FZv7H4E3QySGtmYEQUOHYcgwJ
ZFIkd8V+vZN8v2SDhg7mdyf9dzfdbD/I89MLngHQIxCfQ7Fnz7bwwu4/noz2+efazVq4jah3pfK0
YKAGq1ZdGzLqAMQqWsxCckzDQpJQRjR0MFos6LGxHcAIGsZTiNVNoPUAIGWoBFe5+6b3Hl54n0r0
zYxXR9EneXEDkS3cmhS2OtjbIUdaLBT/KQOU37iuZsO92jCDuwmUtEsBctO6p85Gd806TsY3Q99P
jYGujPtEBfnDQcvnGRkgGDmlgJmdw2/+/4KIxS8ekRFGdRzz66DnrAES53hg5LuRIDOjukWShVon
rsFUBpT33V+poMlq+e0FIXtaMU4kEix2QAub0l0RNq2NRkq8vOg6+n6bjobx730wfVPFjzpdaWU+
HrgfEu1jlEmAolaTQYqxjPRUXYKLBJGOmKriezFp+Lyxm/tH4LmTyIld/dJdzCg3Mfu101LFu/zp
7tgqkoQozbS0+ykUhz0Ucv+CdEJHgFLjUAwY3rZH25pUanXmJVf0JHvmaP5/gk3/jOit49gE5umG
B1wLxIBFqCaA8shUy3wSP5OZ/Cblt9TiJOf1MAXFVfHrT3ywkolHep2J9OOfrtatVa34l1oHrd7c
NuxygFtjDEQ8FogiyS5VYfiuZqeYsZ4Ux44IwHYI9sYEYIw8HFTRtKsIhk33/7tXpECxrlJHJGik
pk6N7/SRadFYcuQx0HdTLN/MySCbhWSZYQQXbdk5J3cqq5frHABJxaYqoIkRKbYIWtuMvtijlsKo
WbE5i0YGFCYxXix4w87t0tTKepZoKx4gnSjiUSQdBhsy7t69Lp2/tkcBFFmTWXwe1U0uZHVHLWFe
G1DCkX1w7BArud2K21mlStw7M1545pHED7OZ9GP0JzZOSwzRO387jnlrOK1fmNm0vV6/iC1Wxefe
NAuw6J0Fjkabg4cmbNofQGG6WBebVPg7vDENDc0OHMo1mOYPM54wOFAOZhUuJsXeDbHz0+1I/qOw
U1kji0GYn7j4jej3MhWnuzxNGwFbIFEAz/AlPYmkFd5Yw1vldL/7o83NuI5Hbj0DqAk+SCEIXtnl
DkAEi1ZNUK3TnQfwdIkt8mRLwGIk9FBpZEkCSuqhcmtoz/2eYiiuqqjJK6qt7CKVxJmmAXzvqpsG
KeoTQSAV9v0dwRSmjvd0kfqSfmMtr/JB9dSK+/6rm++sO8A28L9oNmZASveya9Vhs8/YB66imMvF
wNOsJJLs/5Zeg5PKRbZ9z22xbdPf6ygq/w7qnELt9Ooe3RoNPkQI/xJy6QN67IPk57RaIsnmso5x
e6RG+yg4KMpT8z4YSc56rFfKAgoEdZYAxPprpEqG2CuE9UyIU9aFwIjNCtUTh0WBMPl5DkRiG6g2
VTPKJP9fir1vAxTTM7wAmJTXIbauTczWlCPQxomsKGcXi2iqjsp0gFm9fxF+DfvZUvSdXPTyECm+
xBPPOANqLQA49OtMmz2ygb65bI7OH6Xxa4xphWSAgxRuR26PjLPYM1DFt9GitDlLV2/1z3OBQNFY
meBMvY6HEX9A8NRXbZR5ye4DdngHZVJSPX5CuCTOlUjz7YS/3jXTxXO1qopXZc8tPtZE8UAFfryi
+OHYQT6SpNhZs50WHEAes/yYgZ55ydBHcUosCqTQZnj23fHIlgE9wErQKTrchQUKeg4Pni5O9tCg
f/OvIxeYp431D90sha8cZph8H2p0TPwaHE5O1/CJvi4k/g2Dy85czeT75LV9EMVs1bME+HHaB/Rj
UoLnqEykdL+IZdUlK3xynhpefOfxXRClZacnLjU9LmsXRFTwPOzYpM0OFBOsRrEG53JuRaB/nr7u
/X/2D/3MzmHtiXAZkdF3pICC7sgL1i9TIgkODGpX4nuRQ9AYmRElfFe9T7TnfbNaGKaK3HQl/NND
4Yax9x2RSGbpXO6nWdYwaWhoy6t8rDmtU0UnLfvDaiSxAwJKXosOYxkHXNI4CUz4km/7egeulc07
sG7fBnmzVktiQ/axQQeaH82MoEjLvi6GEvQntVPrEKvdqMMvNIo0DlGvGG3AzT/BS1O5RyK9nQnm
zSbwQw1NaROlzu7oD/84zTEq4QSRM1tTpxQ8eVi0TfpF1v1cvbre3gbXzyGuYVqvxcfFR4tkPLSW
3wO4Jm8thB2EYz1zUyFbHNDHpi5uWZ5aGvaUPRCr53+Q4SQdRBLFFsE/bY/9H6J6BLgEVuafX0EG
OEAiakopf6MlahWmZCDIIZV6ms2JFNRfRJULUojOxte/tE0cPfNsr39ICZczNDhwnvdspGQqB/tc
hRgdWizkm8fct3Sb1mXHLpEVe9wpRgqLDb/4wFWm5nrgWJDw0Sz5KYvsX/dv+Yv8KCayKdqGYpMH
dNm9glCG7rooBEiJ23YPMZFPcuks1YHrQTcO7vXVjVi1fkAArqW5QZam84Zl5trVojoA45FUZ1GP
oNiW4I3zBiVy9RLUw4VBL5mMHN/+wrOxDa3laPo0WN7E2O8SeFNGN8y3AWPacK/H1c+3HvnS7Si7
T/EwiWUhqhosWEDZItEO4v66Dd55+QC5HpywRn0PBNfoNQSRpgFgt5erxVJDB9X5RyrTRAagM995
YUc9Vx6vnZluG3t/M+Mu00uY2H35U+r5y2AliQLipwVyMKlZfRq8Pou/RGxbCz66d2geolLGWe05
2yw+AQ8hNMwoyMtQasniRu012LfxkNfwHZAtPmQ4YH+q/0ylZaTS2Rxueyk+4zVRAhJr9dtTFcL2
TXEVjrBSw6KcslYJeX/Tln5OKixNfnLln/gL4TH1Yf37AMugK9IO2DiXslAt/eytGXmYYfN1N138
AWS7LLScMkKLuDEij/umTI/2KcD3nu94NYZH93s8MKPExqIknPySGfVAhOqUKnY181kA2YiR9iJ3
g6CKP4tqjfiIm342+8OfmIo7t2iwn0SbZnHuFK0YIV6Gsq1SmWORkhyDXdl5j/s1zYFn6iflkc6z
FTr6w9laHWG3NUxYsZFJXmpxSksq7X3Jxd8V1TUl/fjQNDQFb5d5h2fk6deprDT9upUHloUDcLIS
78wzotyOjrZXk9Heh0frQjpUBgSrx+tNjz0smRD/xPRIfuVrsGKg5RI7fL49ZSJc2R28umorCdWC
4wFeSCzeheP7dW9Ml96mExccc0W2Dz5WJtlwSkAsIUJdJPiRhJ4A5q8dxDIlQcoNxJQjPCCRup4M
W7dPQcWouOjsZ4S3tPbxNwlJwLC/D9kXjW7JSXr7znNQzqV8bmBybRaNVj9eABkVPpusb+c9QTJy
yhEcPYWDSr7mxUJ/WsWu4LTCsdiyvOS8GWg1kYa9YgSuVMJ8+eTfJvlaODwT+5nzCaDdARG6Z8GI
pbXTn0NnOUzYxhIdNBvQDwERy74l628Hxjl20TVJXJhN8OP0tNGp1eZIaRhL5nTmGderMDjjoN3d
NhWNi0ysXO56KFb4SpeXb98slqmrnbu6q6XAl+1BmLnjhwZ5YBZ5b/7olvNEVPOQq9Av9xnFLQON
aQtNo1RXXYC/DU6U1LDIr/IJRK6y/4fYB2njN0b4tZXWDep9ktaIzglhcJi1b+qlYm5tT7fnv+4I
/Xbf/oc4KoQJrAzW86GS8W2Ymaa0txuhfYaNpW4+fLiZX6V/+ESJ/INQq/s6/zyzYKnIFrJSL6kT
fRSMJBYy3uVFSWRQi6UDNED0xfY5te3FQXAXjTsbHb6xCCqhNDN9v8bhJoC/bLI0LmzbXLce9K84
t5LqL+8cPL2pTrZlzF2mVgTeAQLjCeiTMmHiLjVlfCGpNHOa65//wwlHM8Hr7c/gn7fFcjEXCubl
rP7ytJD5TdjVzZYwmZJz0j3HFCHhIhL48txPDGOOLtDBZtL7x/f4x+ADMpQYLrgXqtwRttuCCweI
gVrLlFYlNTRXBdSLGpS91wW7ma6GP3EelNDOXAmr2dwd2Y3eCpMAimn0j9VC7rChNug5DAMtQA1F
unl4Mz0rwy6bQrnUzjfh+xd7LHjvevNg8DeVh3xjS5hYk3H0S+eCmyPrOpQ8tJsBDYuJc2cnkVKI
JwUPy4zGZvcQwVwDhedlJQat3YVROu+OiOsvYSV1fQmSQM7yp54uAk6YqRHIPHmiFikk/l6CfhaZ
attEKatP5rIG+zwSkch99rHN9WqgWKUcRkWNdbMM6RF7KOaKCfAWScQMsBkU1ZrNddQnJgH8YEo8
cK7AYmR6/tGUD28Ec3QAwN2vSrnqspuTxJ6kkoQyF6aNeeuR0LNi9SdziOI6FOQ5UW1kk/1hcBcH
ffhU59Fqd43aM5orj1WYK+i335ZezKQy2vAAmPgb07meIuRhHI7/Bt9U8pSeV4Hpx9VELN12Lxhi
5CSVRUGy8P+HcEfOjZ/BJfnZ+161Y7g0MoKyGIX2/0xFSCfk0+5O0XZ3hyNxhQzM0RmiNHxRtI2x
UKkd5RYPkpTw0toKuwGK+u3gFJbECs1LFhF0GChSYuQTzIv5igFxdaEEi9vLcfzWkYotz+Koeamv
XX0G0n2GZsfFcKTsMEakDzHQ5GedPFFSyx3IX+XqRHMU8OQq08B1n/uiBXUnVjLLfhI5Sbqp4Dlm
TjYwwP1G2KW/FdRpTk3NMV0Eg6dv65tFoB22cvd0/Ex0t2g2Jv/xySo44JKrUyz6xSpFAm6+iT+u
zVp+Wil0okwix3i6vnyFxTh4NtRaSBLW2fPURfGN5wbIRCdr7tNvjZG2unT0daZwU1/obX6uqhfG
J2BunLRjgBdIVF0s820PISMpTs5tNGRABLU+XZVOAjkKArQRuSEAEw40XlZvvKhWErtqOz0qjPtQ
OiafwW2lQAAGj9dMC6lIJqopGwtWnLR5Pt2Fjh6qwCrDpfAwDLGwFqKQMH8rsscH9GwKItVc3XNP
Jz55GxX14FEhiTmeJi33btOvr0CR9Eb+2t4GOpUjpGdPnAdUdNElbAnHPHdYABQglvzWhXZzXrO4
O3Poko1GTCo3IbCxy08G5aVQFL2JqUplIsXHt53yusviWvPiHRUJo+bEZ+YUkEgdg6Q4033YTpIa
ywpDPn+6reqKsO2tZEILJbS4ubmmoIPGqUSOgmZDHhVoDkR13cf9i9+4Yor8TQDO050l5SWEIIHg
HK54QKMeKhLZpaI/w+0XtY2AZUPU0e/XHFNwbBNKSVbP5/aXJ5C3P5Z+HMtPw7fn8+/Fi53AOB60
25nIoHhMVRqr6G6BKg+L7bh2dIs92/xwSQVqvRsavcnB2AdDAYSm1AB2PymBe5SQKx16ACGQHKVr
vhGdQx1B+f89v1uILEtzzWS+gbE8cV18UDcj6xWcqi5LfqIooL6xzmjivTW6oFFwCfe5WO4D6Rtk
5AM2X39SLbGPmRXZ1ZjDpT0Mp5yZLROe3d+j6Ozo/m9m+tR19ueZeBjXRmbljFIKmqOhbq9cDPhO
Zseq8s0jWm1JhNeZrmHq2QGXg0lAetFWSASbT9+6I7FEd/0gSiEGEH5xrcEJNu9rtFtXVARRbog8
ZgqWCYUigsXc28Z2rRrojuXmGq+Cp82Hs/ie9M8qAlwQdlGDQGcBfevtuL0xdlEzTaP1c8hCAEIs
ec01gYwMjwx++VxDQIOGEOlu7PjT+mxX1M6tQ/SR/MC3OyzqRH5OKGES1TKI8ssnDmhfO3JwUugA
JSJ7gFg1nq8zyRzOwY3pADTWQVtYBSn8vW8BTxC0K5kq/+Pk+7NLYzN4Zc3y5GwKzMLQ2w7Um2/k
VJQgwQn7hYmtqW79qsBB2P8Q4cgeWMfwMmAeI8ko2EEtixotIup8oYQUhyOfxTcmUb8EtdVNSQkf
u7LZtqVEibC+pL6OGyUHsJXJg5NOgtFUECeJq7is2/vWBaHiNGrWHnmzYxu0kJPVw0byv3je3A4B
niaTXeY2AKO1/aOLzKyFg821rv4GlgEdvMcyGW4qHH9xrXDyfBCDAL8tCCJaQ5w9NiuGIBPBMUQI
uOiX40oVp/HBCZKRmJ43fMxfcVVB4M5wDdtSjTRCRTpj37+3eC/xvMT+8BxvtUgZT2HDt88ixRQJ
hF1YqcswO7LGjos/xP2DdO+0teLtuxbEO1UY8P/+cHmBOroWuS5vkFrteQU1SNl+g+0wPlMvE8eT
qUcvjITP9oArdRzsE6RkDHZw8g0Sm/qYvoqu8atCfZCUJ8F8/MUCVMxDrmjc1X/pRWR12lBHzS04
7rCn4WTzvly3ETvyuWR7vjuncaWtR0H7d6p7gFCDaDoo/b1GHZuX9ROfvEhAlZJspGLUP0xbqUhS
w4v2Ychr69CwuyXVjFfvqu8z//0SC0V7gbfPWxfl+dvHHg/3IJOIA5uizQXSswuAcGnu5L4TcRU9
SJOXz7IG5Gb5nf4K9ouGJntrg+whifdWbfepXO4tbL2jVZzpEYtRXiyGpFgcvVX1t1mJe+DTJtUh
h+kYaNGpqbXptrLbbDkylVNaci0+CqwAoLmsHspHbg4G/kK55gqF8lBwNWRj46trwdkip1gBZeej
RRGs1EQtmYiFpEBKw7JgzoMOvDUkiRVy7srNsaCq9e86pQdR8zeP8VWVxZ4b4yjJWUb79mmaGoPB
MiH2VI1ubYFnE6kexWytsupsKBq7d6cqyvAx0ZhtzQAzO2ko1hLHbYbNxO0P2u8AkngJZXaIEo9A
pe6kTZKz2VH88dW3Z3fVXL9RyPjM/h41zk8Z+hsO79VJxaPSqaemskuldIMR4h9YX+MHVpxtGny6
QcZsg/BeY3M46WCDy0GAHKKfSGMTuRheayzyYc+n1fLeKwP30Y4f1OO2UnaR9Rv8+dcBI66PzfXK
dD1+9xA2s71QU+nzN/MF+nTs9U7diCyUFjPNdhNu4qztWQM5sTQhXTV2Q++upn90kO9h2j72qE5S
kT6hZyzyEOYqPQoTool1cbbwrfEmTEI76a4LL0II3rrNVLSDTWj3VFu1UNJDEr8D9leGKspzTyYC
h2+xnDCwbZxJJC1ZBxEjh9Uis15nerYirbxK1uv4WymhhDohoxfA57SM6WdsF6KZyDbquxAO0R1E
O2MBBt+EKNTqw2mthuxTI1oTQo8/b4wUNJzneIjuFCBtcS8UBZbZAD5j7mvj2gPi4i51OUMhbHzX
2t4AFqZk8teYQjSTiQS/hGX3BmMNr1gkkhKgD081LIXnJh9G+3QcITkdlPD896Vi8b8Ij3slHehC
OSbuvM8zfrDO3jGOQTWQARqUUu6UpBuwJQkRI1AJYkUN08I6TIc03X4FtMtnfI0s0LDhSQEhpcNo
fSjgvQZY0kc6G88y5+GspOhvT0y+YuJTvCx0t7YESJrNka1rgdf9geu8IdqP38s4GvctNzH1ckB8
J6MkBvGX3Jp0RVQofgA4PeB8PqwQgtKN3SCK/jzMtsXHknMtxA2k5QKEo/iwLTm3mxXDTVRxQEB7
c7OoWcO6HJh1gGLZOZgbJKWJAYjxq50piuUWQoDsj9bOZALxY3MEFQltfWkOIWvZGmrretrOFc9y
HyDoFy0NaTN1BnIxhjSfAy0pIlbeoLoSRzQ6OxmULlBT0VhlYqBR7oJaHl3vr5dzUk3s3oAgI9vJ
F4wAgugAifGvq6pKiOyBhy99/qkVpFD5fG/vdMy1tKmfHFC2rf7Qkqi/9Bkz7xAula2Wi5tbSvMb
ptI0yG23d6cV4tPfnoTRidzcSLok2AtVtO8DW3v1bgw5O4epk/B+oOXLCUH8x4/5Wtx6r+H+upJV
o5kCKX19WXUv5TpsUA0LZ9ovqRYwOLpPeaIX6cpGaPpFPcMidw0pm9p4QuBN3KR6B+0VmGMgXTLx
9qsYRYfhFCN/W0/iOowuY9X49ji2Kgo+wnfcX+Os+MEr6L3M3FyqwMfTyUqfdmy3kZTnx+LDKUfD
bHxdlMDSP+wRcMI+u9G5fWABmFe9BCiPgD8vGvAyajbEtRa94A9k8+DUlRIaV7e9Rkb7nwkT3Sfh
Zn4X/85pgS0zXpLHvStrn1XdsEvNvu34ADepEh71gX8FvlWf5XK+cQYzMouUMxZC6huOe4qL3J8/
uKhwtYjMKL1NCA8BUjHWhu8VDGADvbM0KUnfsYRBkBS9EpxC66u+HKgKDakPDUbGvvfyvKrbBx3x
Mwmm8SdljPs2O/w28P7P0SqlfbJpCnoTLcXjZOvbMEZJs5mvB9jf3yYISbXd7vwsXMJoYZHecfYd
b9EXWgCVVV22Aqu+y5PQejykxXqsfHC0qx525qo6svYqzk3YuMDcdciypXUIyLvpUNMAOGpQjYOe
59k6TXUg/S5bpGgGewJxRN4AFPMtdkDDQBoBluEVSY8MmemcoorrMVKbkWq/07gR8t43WkMPrkbN
ti4hj9Ve6+hQLRZLbKYsYS4t3uhqXQtDL7ArV5Kh+r0/ySyy40wiPiQwWmUZTZzMqepju3TjcNWR
+V99titCFde5XC4+5K60OeVJpWsBTS/hDA1SzzFQxNR8x1CdUo1AjNxqi2ft/ZMrOwouLAxIDDyE
qhnnMkAuPvrI0ga1ahSrChYCzSDg11rl6QEPWI6v6/jE8SaiV6d/zGlkf/BEEO+Xv2cUKW39/Go6
IwKtOl+j2P4kahzlLyrZd2zvEPfBEJwANHydg4UKhGKmpOMk5zT4zHpTuunc6AkkYAxVeP6Ovrc+
l5adgwlS/tt7v8/VG5c9iWbjXBt1TQoE8tWraHFCWPTIrCfYDLIFtcuGBECNZBCEj1Q7gIX6z3on
VMoDSqmobJHd+V08jm1Ty1YGYCbCmsOBhjGitTRXLcG5HCDWLet5z9iqV1S7v4sJ3Ps+x47rcoOf
SB5dzaxhCtDSCdlMZUEeYeznvNpKi/6WGisrcYLuj94XroZ3HNxUt4IxFMAQxBsZ23SI3HsjUf4N
NMXc+qEvu6WWnFdr+eRmx1Ry6/orUOEa+YElgkWkilY3ie/DeDlt2r+jjKZWcavJ837LtwOePA+U
PlbFJ0eMMkZlAnx6BP27hmxcLeli//yTL2A4EWvu8FrYSmnvYymJrFnz7WPNbheeRofegeHXzTqa
EjTPIRCjhn9hc7uZ7j1Cy+b1zcqnCrnSHaYnpyI0z6zFnvGUSHcqmpm1cfIeRjV4ZvhNkTqkVrR4
sfTB1Ro/hqhGHlO0A7dMMdrRV7qpdrVOJ56gTzyGLDrNdqSV408/rNWWPnSlQf7DgYD51lHVcnXH
/3ill8GKFRZtWlaElGmnT59Iu7TUjWB0zcgLB4MuxpHzt2LzP5o4ORA8EtC+duqclVwNt9xWQV5Z
6FRi7U909nWN1/nI9WBENdrPQdqja3g0U3ubrrnJpo7L5Iu8YowmEwiVh1ZMNR9mjBoKsou+vhsW
tu9MOa1PrjO2jNyzBfzLg2cfJoqvMBb3VNMahae7J94njkDzucQOD/NrvM1pWLmsFp5/La0ca3vW
QIwPD5zjEA+Zk0t7a9ssu20293QhtQnjzdb2GoUEhqgK2lXSEBqKVvcF+NiPKmeyF0szKsWUCc6u
3S56tm0F186HBdFzMeiOvMxBICp+NaqNVmacs3rbuEzAz1CYcno2GrGc+ht0loCY9OQlEratP1lq
7UIM+H1jURXsVhA3tnBNnA2VLhTYeCyEQJrT1qVCSQbcLBedExe3OJunIMDPDpnNALRfqY+dBEkN
T0cm63R/nwjRjoPZUF8xgeIXOKSq7QNeE0BpLIowHYEH2QUrVMgbAarR+S3NYUSLwbXiQKqvfn4D
a1HdygWZ7Vd/BjljMceSAxx8wDWHC3kbGzM0/u6dvZxUCmaH6ltDnhEmiRS4PDXLtF9eyDtEmP5B
F8VTdO/Zhp+vv8jnBNf7Kiol/51Vefu05BQnbjbj7gZHVzGAHuFotrwPu3qwWTUyZ61rOthK1MzM
Ufqsh3vpcxhblh85RbCk4rm9ldFPP9Fb0sqCI5k0uhU89G4ILCzBNCyPx3mE8GWzWcVzpIaO2daq
TG88xQtFmdjBORFFpWFTvbzdhURGX+C3Q5MghgGO8Frx8XlMFErwVWu5gbi1IjIy7u6J+h8KC/7h
E12OQdlwpkyx+icpD1P99xYLQJscw+Ofh2+LTagMwhshCSAPRdEyvBjRoJBQLOI/yYaqb6VucmBl
oG4kbo17EqLc1TlTYD9uby61j6xJWMwiA6qjzIrhkmKshhi3UwqWMX4+B9Ji/BpvAIv1lNb8kFnh
PA4Nqf4qfi9H/ovcopLd3iPCD54SHIh+hnQnt3bBG62ryg1p1j4mzxlq49GyAbfkxvYsrWB4jomT
N4rPHXEBoGcDTE72htMCx2Ug2cQCWdlByUVZmaK+aoG/Vcnj9MfhJaE0dOUoAkTZc0nGzibduzuv
vRkhpkEJsojErGJzd4hNEr+97CHNk74M/rYXb9ORxislz7u4avcGK//tPnImZS/PGWZWZJT+37JZ
fDDJIYoVIwjJkfoziBUX0KR9crUi23hSVb1qNcM+4ckBn3XfLcjC0zfFNJ5TTeiERAjhbHcU2B9i
HbWrdynjpQetiFYiM1KfYrpRkHGDLu98V9MY9IOBqja5OE72Ap36HfOOQQ32NyamcUxV5f8iMkTU
UaONZ4GhsO7494hPYlfgXVRsmHtaNPLOg3MWl3oTSdyD9/Qn++8AJeWp3SSliowxAu/TtgHamctA
q6r7PkW61n3SbOV+6+TZPppD9HlxO+Jwc2P7AFvUpRX5NubXEJjBYZOS22Sw0xWs4A+KB8WQQMn0
ZQ3uDXqQKlP4ufDAzG1hxu3RNv0AgtoIZeqOricpZyVsrn64+c2yd9sl1GuboxQOJH00RByL9gSc
u5EjIMcLQ9xuLWb5baXPVakW3pDH0kivx7Zw0T1T1jrw7mV8JYECIYM78kFyCxH8noNZuTNXvaYa
DHKxurAVsjCr7twyNdNet+cxcDEEByJU9nkmkcSawQVpjnY6GYRX9kCE9XMHpzdf8Nm4xx9BFrmj
HBGiV8IwvW4DD4o+7Xk9rdPg3t/fCYuNU/lkXLRrMWZd3bDGNc5rAXlQfz4MBkoIt7aAr3KFmQKf
zyy74FvciQ7ZgDvspi+4XCOufoaETbnhQsDBxQWD6+EeJsQroVVRE8Ipnc1ypTJ+86Ux/5DjavWl
BamrdkWSHhOrsLPTaaUk51eaq0uksEk8FN+46lvrNba88XCQ5AXgvkF3rEsZbOFmURPAMzEhJKC7
Mo0P4yEOW+BHskZ379YDx4A4ObKv8D/yOOrHu14u5wUB04t8tMbvOKcBezHwMK6f5/6R+9k9K+3f
aGUi86kuiEqAM1sJMZXzl3tk14XX2r6+Ah2bCRgiRzkli/p7Yb5ofStCJ9jK4xYELIiQg5D2qpKe
ZY8IGipH5c7za8TwZZHUycY/7w4q7oubnyOp4y+BsNVzM1rHC1DD/pK+eYTZZWVb4PJymIhwpg6D
8P6EZk0v851Oex4gQzEIAZZGQ60qxLQWXCnRyQk8CvRaSLub3gPZ5a1uAAd6+1XwpmfAyyR83zdC
ZxGXSOXLfpd1KoY9fiCsXWq4VufUWzVFZzgl1QPdy4+Ie7nKihIwxpdh3NVT+5icHQxs6JBldUVn
wmFgxBkipVmnmy5hm5A6b32OkycA+/VWAi6a0APmPwOeI+ehfj8g97qSYu/W8pchNPF6Qt3wIjrJ
QIjuKx0IsU88e1gxfTX4G0Bi9Z/3Xv/pp8+aQjSqLLakIzeI4eJgf8A86fJy3kWP86Wvc/LucDCj
yusJNNkjNnk5igwI49l9okLssC3rzmp9evZGOoCdLXH5/OpJZEqnbm+hnL2cF9w5Z/jIUexGr8Na
YZiMldjwxdjrpsYpNwGTpwpGiA4KOwvSzD2Aw2ZjvDbOzHGQ5DxGdBuuV7X0UDglDJ89aBYKwIMg
8XWHMGWp+HqxsI844XEHZSxx3ngd6HTDjdjQ2+mIUCehDRzSZ97qdk9k7Wf6VkV2z25iok/vibQd
Faujks4jX8M1JhhDahNKym2F/AHLdsVLcMp1L65jklNx3TvqPq2cr530oUQt+joEVvi57ZsMU5LY
WvtU0w/V9Zhy/pJST01VvURanECqc9mn4v72294OoQ1zbGtR59bwx51oKDJNYtMoHISJ2Kj4Fl+z
S1b3WG5Vd79jyfWlriGxlsUkZzDQeVOE0R0EalBtxDxB12+DhZe4PlBzeZrsRu7XKiSgQmb+Zv3x
WK2aZ/SG2vCWrcAkezdtgs08KomOHnKOMRK4BEdRzWDAlGcqFsQgYGU27pilyTDV/U3GGx1Sml7F
pxOs5dK8Osk8JZjk4juNWjSRfzOgRHSRy6Jkjo235wI6PnDIfbsLJOw0Dj4w+zGAhj0JeTV/uHkA
tbNGCSFa7WJVB79nJ7EilMXM/XYTlZE00NL3rH5DG9oCBuj40G9Pgjo7P0j1Dss9bJugO4nHaM2U
vuVXSiPK4qbZ5mcoT6CbPb2K6POrw2l0QPfYlo33SSsErFGekoDFryurYC9ziJSIhXZdRm+C1aNP
Lss5J1IIPD5S7+H7tSXOcpzuMkF6uPTrTuBNZHaRNUq/V5M/YlY5zg96DZeBXLyMcETkoBeLOPlN
1rPp+wrGZ4CQwcEYV6gub7H89KsxJ7J0MOGKz3cK9uWdoH84Zt/s6JxlgY50NS5uWS7or548/iok
WxZ/lTy2+Cjpuqe2pNWmO9F3UX/dV4YtUeJIKl6csnb9VoJZmMkzvVYYNYNBbZOS3eqJl2PfaqTy
e8xvS/f+wrMHzVZ21nSNbPvTNNF2gSYDule6lXkodVaKcTKU8fg2pgu8zhw+pKjtHWkRjKXkZbl1
lYlqCbpMva2NkcdtDDSeybQ2EwuUPOg/wf1q18CPMRDyxvNB6urn85zfjkorxjMzmvpQYPVLeKP6
PgZLeRyGwqorSZEglxwXkziiQgZOvIOh5RHyEeyiNMNrdEpDU/YBNEbe1ovJjPloJUBihPcJvmgR
wDwsOLJegxaEW2q9YIVAh6tPd9V4Ww+Usy17/cHTZ6XslNUg0+CmnvBzE3OjQRCI8hf8rmhUngUy
J2fNLNtE7RyVs7ev+QcQkMM7ecxdamZB0tNRK0qWPeFLCsz+234yvqTVqLia/xGv6cBjDImeS6lO
Upudp41wB7UX3zeZKYe9N6KdEq8EmcEDdLag22pL82EkBCFwi2pXvPBPPmHK2x9Y27+KhY+OtJMT
KycEAQvqmFyAnpA7UOKdsWDXCjg6Oujmg0unIYy5rWyWmAGMGrjDx+6E+b6Do/aC8zquWsL4Q0W2
I38QlXOXP2xlV61jm2zT+7Seh3T8hyvBH8Ea14tLzDoRYrKd1Ea0dgYZzlh1AaoXeJ4ojqX/5Xn8
0stys4IFDsjXPSlcxcQSSbI1jDW6mmmG0fc2W7vnyAoRZNsTJC2FKr50U6d6GNF1bS0vSbfW+F+U
p2z0Gp34/Db4nfv3JIgAnl867it7CBKXjbzXLM2sD9tjCQupQ2Lo5WzqkOqtRrkk0/XkJzKEupAU
8B7rude6mZkB2jAUZSrmVMHA9cS6C2Vixrn29H32l4e60vkfbhfUynIGyV9KqUKw/TRJMGmrTAvL
FpI8c/ThcYily6L72RSJTrofL/6TcpDfC0jzx6m03APpxFjyAxAhqxp/Rpd951l0DXreG4lrgYVa
cv86YiZD7nA7ZQ+1mSfgutlrhrMwZ7uKLlzzIAqhE1LZ+XhhqCGlZL75vRTz3aga5SuHsGWuurFx
Kp0aP+3Sc0q56Xzlvjevey9LlZJ7LFPyMlBA/QvJ3z0j+dMMhz2QSakOV9y2lBsrztRIo/XWIGN6
vwxitrI9Lb611EdFNwsqNTF+3zJDWaIUsVa/pm/+vO/ig4DdcQmD2OSdwNH5RledSqfsayTM/U64
r3ib+p1vYLMM1rPmMRVaPDIYuVMchXc3IHHbigFrzG33YqVBL5KJJOmSExqxD6teEqmVJSvs+iHo
FKBr9DDSjVTemSulDtjRhhELUSrBIpLcTQlwjkvxXOVpviajh9cv2CMVwBL0j7WzLEIQt3VB5hxN
lwdWB8BrvwAGn+OQYzwzKiFSLaxGTLF6CrY3TOrlcy69DR4P1t5whlWYhc0l2JXUhb1B5v3AChUb
pYeia96fQ/iEAhkeduyPySYU10manlrFjDN68M7CI65Wr7OiA/tpun+//gM1EBlBSYp3EAyg34gC
LHAzhU1jXxb0P6jRm6g4iv6d4bhzx54CMT44ZjytJW76KahcwgXVctbuELj79urUA5PRq5JJzHg7
H11RWAe0cIXs6mUrthm+8BlJdbw2t75Pa/HLzKld347dEumRLoInv1xnflMwozlP5KGha87qvseW
mGcEYog2tlP1aHDj9pu6hsIMZWm8tZm4Tn6bGDATWxqhPwS7vn4iMstl2/sycj8Q2IH8dXNFcoW5
/ZgENvQ3XUTe8q7ZA8KSRfkKv9bAOLzOI5mxA6cfBQuCJsRUf5hCrckTXt7q4MQmh6VVUzpOTmCK
rieHYZUYWzXxNA+BcB/8bCHqkpDkJw5gTCR50GHXbIpj3o1vPIQkimOsKCJPlA4BMc4i//aCSoDD
RrKTWsaWO5S2rUZOxwlejVMgLt4izAjll62hYc41APW7cxVXSZlF8Fcy/D7itue0n5SzugGW9nuH
GocV0PG52STVHorBkTUP9Km65GSTFgNcFQqDhUsNCJ8ieBf3OhBSOpNTbUzPOuUg7kWsV7l0Hvr6
r7T89gE+3ubrOKCaqLPZXoADVPpWMm2Yo8Hcb8Y0kaEHn/D3aRVvQdDiO1sHWcr0E6x/Ya5+xsON
nFLoxGiTWEIPC12bXOVWgNOSOx3hdCbTYSMs6Nt2Mllg2kSu10OY2IKKufEbOSC3x90w9zxZq/MG
Wlvtsj2K92FCinTcNsyAjpNpNSV4SAbKxhYnD+s4WGcpGsZM8DfeAj1sZneXdKbZVVkZCZzHiBBV
7mr1kOzeXKn5xq/CEnnbxGzJGydRTCKPKucahRYrFTnfPlN9T0Ipn220YysR3GzOj7/CaaFrmJRG
+f7t5Vbw+L46zVaxIakDW87/5c6Ou93WqIQFJjQpVdMgC2WtQL22FIgqjGyX6T9jpJTkVpRre7wc
wJTYR238TwMfZdD230NrLBYs5uajnZeC3IdnmnBZiOV0b25CtHMvLFl35/5SC1Vdw5cNoCItmnlN
JoZweLYRDtq1oDGg6H/v8A6Apuu1lVllpZzJwLy9avMdHiaFHFmZnEQ/Z9LzxNrqs4lB5HjB+e45
WP4+2ae6O3SJ9tI8Y3IKL11ci48cSj8/cqpDR40cZ4ciZacyUNxXIiY/aDDs79rKXSSqwlYd7IGB
7RVnfEYp5z8nD8W5eQUc4wymDiA1/DWZUEnItsXIccJjcFk6MvsBQ5tR5Edx5VSTjwBaBRNGY1wv
n5p7WxrDHYj1K0KDqQ8kOFSZ2Xdvv3ZFwIOAcIxBZvPO7JU/9Jnj3CKiQfEJtemgACL0brPoWQWn
VLoLgUuWMrB4Ob618M+9+XYWnzl7cS92d9BilJtmLWdUzbrwUf4gr4UfjLnpqOLL8J1hY4V5yog5
g9xg1eIckxYIbgLmZ7cHoipHPer1Lm6mPJMstzViAAZlfYvg/wwkQ1UjmhJd+EsqWfjLoFynbXq6
cYcgzdsmoanBiO1i0YrnzZkCZ0Nex2dyi8sC7KkWda1W/W1V9NjRnzVulUerzD2ayPCwRUihUJVy
90JF28Q2xKNEL7BNYeF0u8ueg9LzH9ef0Or/xR3+9cflf/TmXSk6EJvuzLJIHoub7/XA7CBJKVSj
YiCFTeq78rQElaMTh/4gHPHQEiXMMjJFPscFHvD8ARaWj5XOTX+gfpj7mA98kFMX1D09ECcvCULl
v4bFA93hWHVxupOTjoqBGSGHYwPrrVB0yUvthZwwEVVpbneCvqjVFeI4HBd6uDx1oVCI4V3+ojB+
2Tbq3LWXFZ9lTZRph4oJYPkjEJafFstGfDluIb9MkAL3WhSR9c7EI6QE+RWTsMiBPL57jU+k3k3v
bOPhDeVFsBGSDyDAHaNCv3NCoqdh2SFLHf+0weKvsc6pm/LcdoIu7p9coI7lZ8P3xrjtOydLhx5E
snN9jW7+ByVHG2oZxaaiQe2zv1poq34Xc4eNemGJqqV+SHGKEC0ZnWSea0EwjJKiXYVR/YbUfr73
vf6kA8MzvFbE5+2C58TmdPUCnXa+wCjzektorG/UO/Z42NZ6gONYhui+eHka/fQ9RonNugLoXqgU
hgVIfb9X2SzL72pR1gkpxTMwDoj96n5j4jEgT2mKrQDebmssknjBkXTVTRnqMCqf2bsjUZ9ASeaE
jOXby61zEEg6NXZFGMW+7Ho4x0RLYe+4PgtvY1ax8yh2xm6kIlOI5eLPnS17r0+t4QlkaltqH9ng
7kIGJofdmuOmfGawcze/LOqgMb6yaQPCkqVsPH5w/H0jP8VPlRGkPryV2eiOpAUDPXrqoYV92sxT
8woAkOuOimi27gKE7mmUq9yEfWxnHKbrI5WDFG4OHqegtRfb8MnD8lGR84tRybUTVlzlxWeJl5m7
XLjBbKdS/ExTlSVxR0y+Nxc/OuEFBxf2rXor2I0ZE+IT/OIRH5PZn1+bUCc1LfHeMvtMno6czXBd
07BL13AB54Zp7xxnLB/O75s1PMCfYsYMt9m0rto49Cy9LMllMcgqTrG+ymt4giR6bXkRFgDyOxoT
vEAdJxi3r8onu+4rsx05d7/w0YXPgWRmtvx7YOFOdCmLqw2UrY1fLIDIPf0pckL+mWNI7RBg39t8
gCRw3RkF8swvbQGQ2TUFVLmfis5S1MjWVROV1J3/HLAYf3IrPgiexLymtmmHD8qVkl19q3Les0xP
HbnANFX6UhMh3+GuKR3PB1czLJ2clY+Z+CMnMQGHJ30MUKK0vvPBF+yoCeYuQa89rRT4tIcpTNpJ
cFtb2LUgf2cAfSulogJimneSWFCW6pRWJIbx9DaNnodbAreB1PXgVuH9uYNB4dAAsOnWJ0t2X/JO
KQseaH70t2bUqy319t5yHYNAemjZUGLO3HBaOKh9s6+MrSUmfHE5EoZAhGxr3NNDrFdK+Mbhvhpd
DLuNWKKGfn3omWcEllMdFzIZzatymsa3I4HCcVDkUdQ1C/2+2dScufVFkEJRM2+M4AV9ywqhTmNw
e1w78lzM8qi7vLLIsGV64m6kIRkg6agJMYC2uWNFWoKSVDo1RxY1ZqVraCJV0tjN71paGwyf9fST
wzxDvrl9TToQ+Qnivvhu3hs+zkJcO+oc1kCyObFGWNWOMOjSGHSNSy4CiutgKzOUJZXh9gqOqUoN
N7vuk0IKSTQMRwXnsJb4eTQcu5RSbsU2cQPiYnLE5wBjkUHU2rd9MIdjw9REMPXE3vtM8iZsLYBS
gVQ93CpXCDnbK+JnhlmtoGSSVkI3lGjJcNOVRnziHzhzwOBKx0fb3bm/skbUje/LJ63lVjeEH9FF
Sz5aPEUPu8JDfEN7C6r43Lj5bTrvf+OENhIEbpu2VSPxxBbN9/PVcEYLivyz3hgJVnED/XnJgzbF
2OzVHGmIeXAHrqF6t1loQl7vHdRfJ/jJXNbYXgDqWVjaAHeAJ4qP5RM6T0qjaGMXOkUlXfDc1zXX
w3ZB9km584BRSUvPHUTWC/B52Q29LAmUblxAXQv7/tW4bsTgBN4/u3HOQKn2LHUOF9qVGnE+R4Fm
2HV/OupTBydTD3GO9ULmtxz0wdX5/960EBudLQ5gyPgk3QklwReG3vzRajbnz0b3fiH1oTiqihr2
5w8u8/oMTImH7tNB/tN6CBq/5rcnMLiEFYZAUutUSA9m7QfHaMFfy0YlOfmq2LHAUrqKBoY3LlxD
mWDai49w/6YPmm3rUwaskbcRdPh3XLbIwYXgTMkbDpFT8BJlo4eTItCwEMTKoECooehY1+sK189o
88zsTnSCqkLVkXcO95+o8TgKpIBJ6EdIQJRJSGebqu3lln/pNw7AZT0vZ29HNfAhk0o/EiNWICfR
bRWcdVcSYab/C/AiVrmDmmkg5QI24d9xlfEJdVx5JE5gSLRi4Ru6w2A+jIxoYX4jYLDVNgZ0fSPq
wmF/h7aOR710MRTsicxo3mWrc93Hc8ZNkYgqxlJZhEkuJTQcGSi6I8KAcfeNDqq3ZFiC70edwYRz
3cR1FEvZhwjtfUtDP/XE6OmhlOFTh+uvydiM1B/AFyNsHEOT3qo4hIVx/BUxDXsYOQqU6BjL1jwH
L5eUHnfGe/a01WiKWTCtTWXHsVnNi1YXxtkM4knBktQoUM9XrxSaLMfR8SvRPtZhblTjMG9+6pdJ
Jv3IWaMVWzaEiDmcWOq9F+PLT0JPPz3E2GGF6MZ734SUgoxuNpHkJKMeSM9wCYEu1ilbXOyaImnD
j/sgAklsXiVw8XTRBngKmAJw8EvD3pgecultuXS80eL4Whg2HOk0Oml+bUrbcX+krDXy2dJnkyca
zJwdQiSSeDTwDffaHz5SRz8fSKJaBjbCcdDrpdKUV/2TYtSzmw0nXGWPsrBcdbnR2rwqc0ujgf9v
0jRHz1V4jiee14UG4LHV9lJBDlHHcpvAkMhLxr2gde8CqrCb0YF2/2k6RnzoMK9Q5wYVJdPmwksQ
FV9SRZ+OeBQZ+zQV4IMdJ7KndjDcwGroHLtTfBvpM1OuCG2os6nSeVsCDti7URu7ela9lpe72CL5
NwT/YeFUiFM47P5hFMmagD/gAmUlVL8jNoVGcb+tag9LsKBNLYD/xg9yX4ZlzNloOgSHoleYGQLH
t3vhWUxFrVFJDGq3o/y3cX0vbRSZqGeMJ6wqn3v3C9EqKON3bMVZeJDur2ypRFZMf1qEvSVwTrIB
xDc6xygYBA4yGtwHsIaGtLzIMDax5Y6YJbfG27UimShqAI9yTBYm49MqlLdP95Y67s8AzSmUi+19
O4mZvEMQTVAGZhE30rVcP0F7ewpYBlXsetGOPCfckHfVibCxPr97Og/oURawzcAJ2ROyCdLysmJV
kiaHSLZnsLIaYRHBivAH0+AbSYY45kT+YKkG9KUpzpfZXvP68X709d7AAy3cTiT+vNfseKZ901hT
TPHiWpu5W49ax61nSMvANaGwUJnuvFfRLPGNe7GfnE/xpJ+PwLDI2SdFFGlcdvOnTbazuCy7hba9
0zKokE5M/9kO9rWkqIH3hAbsJ+zo7K/zllEBCUY0+sTps6wlcPCJuVJOaO5svIL4Y8dOlhWmg0Fb
O7j3ivvPB/ji9tr5W/ORTYJypXhF12cGaXM2VdFj5Dda4rkPMCYcsfJQ6EnCrrPRL9yBfH3BTLZW
5iga74KndF6x1HRlTLZr8lP4HTcugN78BU9hbLoEPLSnWtgRn9yuzXaX3Abax2Z+cy8MnAwD2BnY
THo2TJT4/qzRCo9fp56GdXzR0JRTVGnqcqF8ggSrUgblX0WewrC3PrJ+9yAzfRpNBMaTMbTbBPKc
TGHFZZ5pixFNGEdST2JjcRdxq93ZPdDsO6+0VLs9xHvvhXH3JpHMRYHf9uO/IrzDspTu+lL545az
rmZdrw25iY4ejsI06tffM4iTViv3pZAJ5Dlbc+ZgW/r2mRotNLK0wogbgS855XomELdTUQRZWibF
pPI0zuFqtgAPmtDM1lNuzlxtQQdk8bxiMNW7j5fVdgSztvb5sui3ZqWzdr8lmD+WeqW/exOtM/+8
kEPa5GlzDhLYRPghQjUgwowk1cs1+0+lScDgQY1gTnBUU//Q/HNRpGOzhuGo7ZsmlpBIB7FicGmy
4p68Lc1+fl8pZY0WwfDQpNGgz9V7i/vgKQH0f22KFVfwdm3nPrlX+2s24HNRFOrldmfgvdKAPHyP
nujegjivfa0IfebEyDDD4FEIyWxtGM+FTa1P3Qq07Wx9Ght1mpS/oYjlnyOTG5kBPrkryKq3JZXk
AFr4T49SgbLLf+dqyqygFlCHKtHaHt43v30IxbBm0SMei7yeheXAMZoG6/gukVZEoAnRGq8Ta+Nz
9OS6y+axiwN+yrI1si6C2SZWwEIdZlGhsURkpktAvuMMQBA5R2a/ACkzzL5F4UlCvLCV+A8PVEsi
Rj28jVXMmKDUkTXOON2oOT03eQ20/8z8AKzL1/qlUO9PddMh6D2bsCqOk+y97ax3XuAs8gqm7AUd
fW4GbCm+sKD6KekpYhc2z7Gh2rAbdGPxRCFXWSXLhXI3qgyMC9PgYDBErhcTm4eIz5dUwPoySgNq
9ZQ/AZQb8MK5W2qtONGzJ/pDoQ7bHG/+jQ/CqWlPgnqw7CY76bMIg9RChpvBUtRaLlLhAJ/wnDCl
wC5JpYoSm1kDIddfhycND4Lm1u0xIIXn9k9ECtcp0Gg0T0pAbTLkY7U00JpBz2pKjS35DU+YzFbG
pjC3cSn612dk171UwtQbg8GO/9RFunJLRvN5ge/kQm+6R1lr4L9NBY1OW5uF4UHkbniwAXSTYexM
Nqy2kJL/i//7CYeRBiIQkovfD4t97NhFNcLMSrqYzdOEx3l6o5soRr2trDGypXRupSGYrLeW0T4H
Kq8wvxqNjo1HXtFq6WYIX+5AMUDlDyLB0wpg3K6n7lhCuCk1vhEHqf5QshCs69r2KH8Rt62LoKp8
YaXZOZUif9t4k8NguaujZJpKP7g7+qkQs+m04Wc53AtJYep/K/+X2cvQKBqszrUydAzDuQlzGcbi
JlMqSKzOkNzWGeU4PP4VWNA/5hHwTDME9RLLLWizX6xVeF9vm1LA03mIKi9Staloj2BZsHZjP1dj
zY/goLVLD8vLp5LO12J/IO2KVlfXT8R3SQbcBHlnTm6wLysUmNvUfrtpVmch0Une/VySfFv6PMnx
YFdfhtPDxWl7bmZxdS+sh4iIyWIo/PfGEv5Vf3Da+q5QSGyOgAgZ7Pfl2sN8vbtuilOjOruq1kLJ
JhuMJdmLz1X4PHD55nfmSvE41rB/wCc9O2eoJXr5LfGqqSb/UotJwaURV6FNYUO4ULKM5ywstRCP
r8nUvZEfAoAuSt+LstvlH6iuRXg7El0gJs5KNaHIbLc3eCO8XbWyt+tI1zY79aRlZW/zDMJLYMX7
vx7F9n0o8LE92FQTe3iuRMywKTMvcTQtHmHh8hmXARW948qVGvBqEdeSuukyXwuaXkmutmlkJ7EE
ZRHLY7UyCMWf+sptqs6GxdD9WCtg6bIg0kIeMZBf8J3QB087tJB3Dhw+0sCIBs9b5bZOGnLCITr8
60XipUQ6mOd032eGHN3y0ws0YbXZK/xDRTF+SYMa81KWSH678h3ciKkpdMj3/yyFmhxO7JCaVb1G
jj8bnbeK+TZ6Z/3tqgQ1OMPPSSD4Nf+IzKVkPVI5JvvYIvnYy7BNn9CG1rSWUdufeVzBG6CFnsKX
AsKBQ3hgUD8D14H31GgZVnaDbWCLkf72m5haBxDWzimvHaSS/88dPk6kZc5MXmogCwTo+eqi5XQU
xOkR6kaLUrP9oxBq+1zOMRyUachwzsyg/qWXE7MRjSoKZJRCIDtLb9QdCTAgJRHcn4lh/rtCBYR/
nW5zTfKji+uUfDXPqjp3sC57+LCyXT0xt0Soae97BCqm8Nz9oiqS6ISMh7j4oT2Qk1bjxCKGzwIL
wbpew/DZo/pZPRadSXuxk7tJHeajUShAOlTQWUSGjG4unbKGsesOc01cOWzHQSzFLLLAAdSHPuwa
8HAKHwzHpe0AlAbnHXXSQjyxTYRMfl7o6FagCtPtqIgiqv2EqGlhk4uwbgLJ5tAO13sJJmh2EY8F
r5iyuz6vsl/LpDURAY32TeHueky31vXWH1TngFE89EsIKKYwUYQeV1xjwGKGHlTigRdc7qJ2yllw
dL8Y0J2EnWJWM5+s+M3BC6djVWNghxNiQRm7yV3HrLEiqtQGafmBkYspX4QO307a2KIkXtI9AQbG
I6VCCJvXJM133r2YbP1XkjBRCHaNV9W6v2QCgftSgA1Ca4iEBlHfTY5yomY8EroN7R7xQ6Nk6XMP
51EeJCmP/k/89siLNpGHDrWZOkXlL82yXAYmjufz++PucUZCqOCsCAOhLD8f+muilGkOzxrtM7nI
da/bY93eTxUrHJMyWMcsM+JFPQjgX5oZj0Yv7aEcxfkPAdbp0U+5nFSeq84eFQBg3keU2Uo4rWS6
cFv38/2j464p5943eqyjJEKIUTjlfRRSj+g8mDR/E7ZLTITOL3arQeV2l3weXjsIsYUnlhyfrHPM
bIIGL+1mtdOSR/cGksbGvRfX5sjsfCRiv81KEHZ5vhXiznKtOT0BwUnAE9cI2Ciu+RYC8jxUcFDA
xUmlfo0hlATof7+lGS2YYhfnUbEaIKaX0DNhDL3arGvDbUfqsVX43POqCSAPBm1gHkzR3NzvZ6KV
jLzenU2duFGFpxwvDcvcwKLd2qlea98Tl/cxkMoA2RwzSFyZOAjGhVBLi0jp2NyrQIfFBBcVVBud
uI97+mSS+GGYsrfOWEp6HWvaYlQ52OeSglgL4A7jE68hOr3lRsXFseowrPaYokMkac1G82doyFme
jnMJAdZl03lvigqPb7H8GNRwrreOhTdfimVI2uHaRw09FpbLsJ1/zHGOmZFuecqyUX/isHxv2r6q
MR29dr3mLB5rCX3xnwZa6Wi1Bi2Cs5tSkvITeCwIwx6uWqdKoiilyedUgSgKpPsM/YHEu4yGEItB
VUEh/L93YaKl9Zw2J90I/rmw/Qr/aAiMod0T4tjTWEx8lXeBBntFoioflku8mNPFxatY3o98pkzJ
ZSh0K3PE77RzwoRgXeMFX8gJ+xw++mqo4+KNhc3/cPhreTr0MuWwnFY5GqEvjt/vYGZutsBt/cr7
TVK3ivt21fvQ+5GZshCefmnlK2SbU2b+jq2Bn/uIpdaWNzZvR0SQO1pF3KLtk44i2ka1qzwLAsCy
2oBpnsOAaI7rn/TMQOciYj/mckJ6RnOqn2BCCDF8OgekJ7uePq2D/PSqLcR5tOXT5ybbzefokUSd
F2JiYL4nSBgFCTI198jgdm7CUCXVnqZxoCqKBxaL9EFKkWPhg+Q/6aI9lC7iqaeaQ5I2g/QYJckS
R20ymQOqw0CXJTSeV2jKZ9WZo13xFRJ9wCuLV4tQp60OGvIopXntHtT94rniXw/k8Yh1cVmTpLpV
BJ3d5srOOt7ODc0v65mq6LEVyACmeQjG7NuJZwgG3joNeI61iq51iRGF+NHUBFk7AVJrJJDff2zc
uMeZ1K03L77GDX1hz0Pbzb4TwTfcWKNMVbOVJiYRvjKL24ZJniNxztLItTj0yeaaG8C3bMhoP/EK
+buqJn2q7DX7vcO9AHoBLKQlEEDkd5l5yTYMQp/VYc8FPBjBo+O/edn3UlYpTLnGfvIVhdeUSFqP
kQ64OS65oHL0498rVFFgvdlCdQ/ilFnWNa+wER6eEdJ5cV6rp7PrU0K/yE2JFcD5IBH91d2m9E4+
QRkZQXbuQFT26VTD2evYf0/e7SRAsfkQu0VZXsX3GuttxIFkoGQ68JAZ3CdAhrtTpq2vF3mZZvLq
y/dOaFEEJvuqy/DrGMCd/8wM6+38UnmInjSHCbLhFRrLiOYdJbA6xr3j5xMsyHLNHzoNq6hle1CZ
4sOmK0LwkYK+p7TdT1bkPYAdOyKSatJuQ8/b+99AipM3OJCy0bCpS4qwVORPKs5hj5zDmB4tEQa/
PkxuE9K7/gg/IooLSwQdGpTs40+i6g+Fxh1pup0NycemA0LDwpB+xp/QkUsiHHTeLN1dc3ZO5RBz
lnI4mTLdhcHwhEaa8v6CMxJVY+OEYdlhgboHljCJOaKVqbTeiPxwfymh4ZueOtVT4RBsBRqeSz7H
ZxTGXyPmpU6dh3UmKGUCiFOe1PAw+Pw6ehhBf+z+cajR3lXECYqdfb7cNaPK04eBTn6CguB6LCp2
LntJeLwVPWwlUDzL/zBbqcgnV+/BIgqUteizlKoWmW7KJWGFUn5ozgxcLWm3oe6Je+oJ3Ir2CErd
492Ku7a9s92VGxy9Y556IdmQY650F8wR3iMwYhnsf+nT6MlfNB2YGUBcEU9nXAYNzlDv/Z1+fE+8
g6WZVLPuFPoJyjYphCZyvYJDLwBgUlGQ1WQlqGiv4uuAVLnLaKStAopEC3YJvIC48osSjklqwaNr
bY7pC+HfXLmC4DmbN6kuVI9ZM+vQUu7+Dtx7Dqmt3hvfD70Se4vVVivWcY4Ye/qxCI70Vfnh6lpW
0rhs0Z8osgEL6scEASoBMWicZyD+5qRVj8mlO0HFSpVj6BwW66ZdSih0aFXvf1GH/AnJYzMktJ2h
t89iaHLwMYlQxPaYaql2+dCTwtogxqJBZ/blVoHWu+HM8wN99gn2r8GoSYOs09+tQLlNpevi924s
sGp6lhmL3OITK99L0uNSJ8C/uwTPYGa8SnfPfTjMEAyFqeV4SC9yFM+J6SaXt4M5trqEQs+L1xTd
uTZ3EPUdsJ4tLxJuy1t8qELryagh+aaQK/d5MO09HvTN7ZPds+o1y+6X35FoMAYEOF9jO5cEwI1E
6SJLrU8hIc5tGuUf7zhiJg4TbZ9VWaIJS1RmP9vxKhEbHjTanSQRgrBSXimMs0INCaFo8gjJyE6l
tSJty+430ylIK2xfXJ52Qf5UIp7CNST46qpJsUk7ILtYEEviI7LVhULeLeO/7CvA+3evbt0KbIDh
0cpgvwjqACK7GO0f1QHjc5mXooLAKe91zL4kBYAvM0Z63zitxBXRJrWjjsHK4M27meVoEMZTLbBP
YfprMlvLxuK/8PUpP1fs4Kealqn/QNPnN7rwO8E2XxHEAl4VKFlpZNRAH/bnEKyEBBGcuIIp7Gvv
P5HjwHaQizmt8gpGRAN4Zjdrm+wUcRTOPOZj2+9f+ZuCuDqbciPkKVGdXcBtUYH0GlRD7YWKKiLD
rEQqL7CByMtRMU/OYumWlS/0bCIID9qvb8V5n1mQnUg7bstblFBWEL3blZC3uY2WZWH7J7TBh3XQ
eYE3CwzOs/EXBnoaWAbKN3IsnPjQm3NzusH5rIAVrR2UA4ly/zkqJv5mPxCWxBv7Lav+0tt+kEub
Cz/GVKbTO/6+doB6xTJiCvtN5ynuimDOqIoiNnrKT2s5M9wIyHKaI/qH5dnn8iHjusv0WaShboyR
b9vYw5poPN4Z1J8IWJgAp7LetJ94BV80ZNsO7s0oe+4fFLPSsqFuzxKmDBfdEUJO9TGRywTGnvpz
1Ru2SXsGSOMbyQ2MQ4RtXWGAl2GR2uCe3vA5fARMI/5TMUcPBj8ClMoN27c38onJjmJ6m7bLgIWt
vNtkc58PQKgpK9LWH+t9pBHcKU+rrHYAIr1cD88WTc6sHB8uatNw31z6u3D9tfepb0PAsPWngnjt
zrnCBmq1DLCx8QRddXZQ4MRhP05eK5G1sqntMYVfyRyHoEQJokyc5d75+5yK0rKYohNP2skCUBn4
xkVajw3qeyY7qKd+jk1WvKl94joKZZ+B4k93Ae8FK1cvtaM8gVT8KHmxhPEfiuUnaqLXiCZykPG/
1adMrRCaB4kJJv5v26tPrq/r7XkvoEuuOItt5xboza/5/s4SM33S1f2fVoPJOVUweFcpfrLXVDQc
ZMmZ1d2bMzthneCaK8/iPKFpLCuEzRfykE/9X3NDpVwYPEs3bzhO5akZg65+rvJSmCQOeEMeds2t
y40BC/mtL4nX4TEeotzoOP9V9WlGtXhKGX1HTuCDWyw8oJdAiWsi7pmrMLth2ZNTiYJQ04tt3E0k
ucbaXnm2EQQxalvPcF/RR7A8H9kM+vc6XgzQNf5XA09c7XQNIlG5B5yXwbsj41ZuD1wJ5Ida6Vp9
YfPOWjZchgvfWMx8/KHzfFUykAjiCi0Fdv5ArCGmT9nasHB2bnA2Zi/p+7HI/gbLq3et8EdMVQAi
27YzA5/UWgsbJ8nbGDHJGSq9DFjGPomFXe4+ymRu0/OYYK7fc66w5Aah6xLpYyIZ14xcAo8i3aJp
Sbder2nBAQnrqCbF9WErFswzhbupKh7eN3UsIRHZ6NVeI/TSr17xqM6lij5bogfx+DT+dnxg1N12
7G7kIzz4VLqxCmGUlyq1BCw4BWwqZ4rcOFf9pRQIMTiel6a05661wYYz1qdDo4JeF1M7KVMps2cl
CL6tIqCMBbf2ljzfwswfPVjnk0hwGW3accISvY0Ok7tPKE/q/ne0okn7R7Y9L8M1XgbwCyRBi4Vx
AHYsLvSK9q6aenUmDw8vXPRtUAXfYooIPZ805p/vrYvZaZ0dFI5CG8SzzfeRb9pmb+ztPDgzuqTh
lbxWC6eLlpXr1DA2kIhdtRUJrg+31SWjsBf+whbVtkdUrh7rcRsHTnjlNPgdnleJAKSaTQskdr1P
IceU3rbDiQlFFcROdGkWuYvH2zS5/kLYRjJs+ODAuysmD4pb2C2RR+sS9QOLj9o/oz+/b8GhCf/C
qNJ7ILoAEnQBTn/d1cbLCpvJMHLRhTzaYKWAqKK/n7CDxVpFeSp2tsY+QncSaAKX6lYB0oS4xP1n
MiZOjqx0KiRcMY5TbWDZXLZUkrbSGgLE8k4ZANKh7Al2yC9lfjfFMHLPCCPUzwAhuiKzArEe6gdQ
hXuWJvaZyY7crjekUsJ4SGz/k+dIgSeLxfpbjgFuTzWwTUPYnjVL6afcs09ylSCRGbTV4QRLKpvQ
i7qfcL+cJmMX6ya3WWOLElVHlaExLIAJ9tq3w6eE+INqdrSa5JFE94arHt+BwITR9JF+GfVGafv4
PepiLqxyk+lCYyoby3fi9lWM2B9eP8ecySeedEvJMTCLBMXVge7GMh569xdAd3/X5tax1jggMDHg
2NvThXWJeUYU2I7tGZYr1v48/LHe+VnhdZRhnAsk20QlZxfCc2IQ/eCZ5lvQFCvAqij6trMXUGt+
O7VfoubXuH0uGFg52PQk5/tl0gdVpzN7X9bRl9HHO46hF31LZREC2RFC9LQS6AkoyMiFlp17XjAa
Dw1hwic1/bDljBELxu4aONxfpqljq4pIoZVfL8rmjI1eqIq3v1+WUlxJ0zMgvnUTBoKl8POgznpD
Df3NRC/EOPOfhOUkj2ivvhMaL/vPW0HyLhGIWUmpqFhoOkzUgmhR2bpEur0rfgpAmyaTavCDw+ju
F4UWCP2rU/zYCn2L0jUt1ZGVeNfiUgMGa5TIQ6BPzIk0nUoYfv7PE+lqnETLMLrHNw13LfMC2IuA
lTnr1i2BP5la02zei9mDjmk87UCsP9MbbCT2rU3V0Q0pSz7WI0t7DANNOu4P3CPltwOuoSOuesXI
kxFlY54ORK/llMUXfA/pFjm7y05mxFaj9qdK9fJQWaKObOzxeydzmpz+kqYPGUBRnveFt3QRfJ6k
9ZiSaUOmTyjA1V66PgAbl+YYrP8LWxSonrlu6lr2PROw/UqkWPa5o0EyYYYUIsZU2Yxf/Vcw/RJn
jJfSqg3ggnDRT+8rSfl0lVS2Mh+EM0mXkb3zPR8whi9fqKQn0DeHHElpAMCAdztAc+BPBmnZ3rtL
IoJZXHX/TnwwF/OsUtApS7djtYsOcZTt0r8hcdJIILOy9D3yRTpc91uNqjsyGrYMyibCQNGri0mJ
uE5X4E+iOOQZJd+UPpHWN45O4VAebwfykolINfZxS9b1TQX9576IL7eBZdermXgSOzwGpEwP/kOW
Jk5LFC6xwOfH1kG2ydswyTK3zEDs1BssrFu48SPIUiOjXg2ZMho3c/Uc7fr8XyzKCFzvm2hmkhq4
V2YQlBqcOq3NyQHZ5wWJMZZiP0U4TWBZITOUbmrimCmQk0xxqcwMbnpQK9U9Un2f4w9zEnB3s/kA
yyAx9tGOrq+HNyqwH4cpfYbt9VlQJT0DY0FvQ0Lv0nVpm9rVtw+vNO0fJyr17X08mhwjynd6wYbB
A59cmU/aSTPWW4DUMLI3Zy5b8oeVClbkRrK7akOShLjB7eOsPRUcklzD1ExbL7otWVgD5wtgXq0v
CXyjPUw+rtTpZKx59PhyoXSrnVRJTWcwe8fX6p9FKQ5s3/Vvv8G0hE6VTCXABKkcjC+6hKhoZmnm
m4oiIv4EcNflG0FMMKADVvMQTRXEXSTR+ytdSNEVEh0NjDUI13W8K8QRRyqHpVGf+ZGz4D38g440
Gt12eYuuQXs0CW+3KmORjy5HCDLml6khVUXR1tTLjOnLwm2yH6n4RvL6UhsZajJfXH9HhK2gKSKY
ADlU0KSQ6a7yN5ldf4dpFjrAdNN4nhaxoK/crXw6AsuY+H3hzDkWzOFU1tbN812xW9yMyRy7E2rJ
fitWI6G58RyExsl6fOE3W99h0igebVnss16oo8U7v/Ru935rM38WCQK45AGOTz0Uvh4YOv4zT2tw
UouX2XhOCk35tjiNFH5CDJh7on2mGyi9CKgOWr+M7raUG335aBBK/pcXRDAqf7iC/1gziZKfQe47
gZdX1adp8Go6awvadO5gToBk1aTFo0v1I7kFcoByG1klTwqY0ih0YpztW3Af7ljgMF7T+NXSGWSk
81e9eafVMsT7bD/+9U7BqymHUk0NZElZDE5exFYYmdB4CXxNrNOVOCFaCAz7kzbzL5+kQxUm8o8E
w/H9PE3sCV+2s65ZvPJWl22i6SnU2p1tQ3JvFtPFfDHGCjEbgOa+hvX7GaQYjwAl0dFj+LltHbGC
WaA9fiz/QZp+chVV4YSt5LfjPjLuDKlTshg1TyCFu3/pvcHB0LC41wtUAcWjMv9b98Adk1X6CJlC
q+8uclgN/Uex3rDHFn+ySJpIhdt1c4+eunez4Nm6O+Fs3vNQDIb71gVXHluoJxOv+ji0XEArC77V
aBNS1cm68WMnqkZN+MfMK/09i9Y05GFu1Qklocg9Wk3tatqYu+7Xv71Cfn4NfGaqiEOzNauS3CRt
bl2AWVpVt35b5MCu68A+fbQ3C+BwwInaK9NQOw+cm5xib7wd07HstnKtkvaVscHm9lts7wlvSzqZ
MYL3OgYQdOV/DNssk0ARx0SMXkAhqx4OcH9DFbpIzvHwf4OgFzI23ZJOwncNz4UHAO8G25bODX3p
A5Fkugu9ogtkf6+jJkY0kkL0/2tvHwCB2Xw9o4EKb/0uo34PGe3gu4b/X3fqn1GmlTLv4bcMVY9x
3QIj2dzNG4C40F2tavG/x9eeET3JMGqe8BzlShqtgWu+uRQ2GMH4qHxCRZqvzp236t6dVdMopjnR
b4+w2BcT6Qq6adWIw9Bomx3skIzBDjgaoQ3lj0QuGmW4gMC0auvvOcu4Rum9sHQXtoaJ7+cmSV2A
XQlGcyKl5uCxPDw8yCVowWPCXUWqR6vPaybCI0rEyo80+qsnPA1lYjNv0Fc9MJVT7RlJ8xUcGs6W
TioZhdpe+1aaAE7+p9uXYf3m2Cu6kGW1mQCx6EuClpzf/oer//yS9g/L2XUHmAtu/CCYuVFhYmGg
9A30/vO+uDdTgCQIZgSDnNb4HSQ+86IZSSGxbheMihfJFhn/Qp/2DX6f+sTMQNhACe3m7awHGs+l
WDAHRIg04Ab6Ck6AU5/0q44FvE8zeSoTE+AUJm2v3dXfk6oJ6O3p7dN5Ovex8mEjaahBkzYbOjRO
pXZNs++1gjRBZg13gGKKI3LvoaYNZA2GqwFDgrPP81pC87ZB/BMeuUcZPGt0Rm6Wmv/LSnF6/rzs
+HPmGRZDvOpjndglfM4wSURS3JVynXIAnVpkyOaGDfqqK5kAojfbmccqaGb32G5NhFhwYjKtUJ0b
IXN+kOzl7NVMfz+0VDwWv4skJv+cVBwVH+bnf9o/usT0z9z3qIQuo6etILk0qhjMZmtQYfZjHJ8j
GtLffACEHyaCq+GZtJqZeDHEizQRwmUBYyR0KmG4sHNAbDeVg02AnCrGG4fh+bZPv31GtbSTvoXQ
EVt4/1WN0nbQXF1/RtH5qFNJgNU9n5cdv0LWhgOhQxcU/VhfJZcj/JaOJsP+18SjZ900nbOIuKrJ
iemvl802HPsgwhRBXHbnQMav4CxUHU1OcJC//fnYabIZGja1JW8CkY081c4TJRd2A/6a9ILBV9NK
eIv/n//FkPcoQMgZYaGetRFTTktBnaMceGl+mfO4gKiYtAiP0mh/8rq5zRb1nxYYi1dsvzh7qo7G
5AM12UCdMBPhPpe1XzZ8sUDL9VAsxKEKNX+gXQCNfrvMfaihwHGDQIby8H6yByBJFsYUgS8S7fPh
fRkt0GVhDsIBsXYAoEOrNK4/TEpTC9xnQ5/cykai7eB6gum+Xvv14uh7D0+BIui4migprasp8akQ
5LDBK1s829fU57e2eYIeIhh1fQjqPt4M45HVxkfk3Y2EwD9h5fARbwV0LvlwWXyEvpXOcrP+ELD6
2K/l1QzigrM6AARZf3yr1EJ6JYUPCOJYJ7DSNFh9D6iEAgXyARM0inY5wAYGhqdY8oLH6JIlQQ9X
Q3ic7VUms9Yb+FCheBazQZRCEfM4b5akKDFLvwjCfkVmpSWm/tT/xKSNqf6qqCmhYJV2418wKR0y
ZnI9dhAWtMJXrNc9A4SMwMUZSVY5kbAHLefKlE+ahIUoXRv+W8Jw6Ui0+8qKkEyCVw7chd1paftt
i9OorAWUxcilH8Anklx0cBGnkR8QKYQg9xCvJuKIFFYb1xJZPtKdLOoKBlufnBK9flYsV6zu+nf2
q1mcuV/1aoq58B7eqWZe7kR24M/4ZaKxNo8bckQA0RbuDRjFSwSVAwT9uZzEBy3uQXOvI6r1b0si
oyWI4yfBAqCiBefDyh1VqdXn64lPjdb4hiqKZIOQjmS4Fk26mn/DkiO6C2ZAlS+oIiTGwZ9Ks66V
CNsIbIYAdAIJ0LyOmv01P7f1wzOSo9GjltMLDNyGrhArwtSqsXW9FweZTkOUCKK6vkNhkOAztk6p
mDTblNugG4QS8qkUwn1WIoF7r13jU11iSh0/m94CV17gmec8xn9iDICd5/PqWM5XoAQ+DGsKJLk0
vRllmuKy9+VErzCDQd8n1YcQeacF5Tdn0kt2DNNQqDeweHI9/uuAYhPFn69xaRqmUybmVgzTCy0w
Vw8vU3D40hA71808HC2mznwDfPxGmtjA2Cs7ibuq5FGi4xkdfo62bOaMCu/YWpTuWBV1iiuebjVv
ZvDRp7m0H6vWolpdMbcrcBN66oKdpuD7/6ZTKPgJd+zeHXLUVoQ0H9MX/9F0FG30rAAjqhLFA5qI
mz59d1MIDeJBT33NK9oLME2mSRI7tgRtx+6yuHmQc4Yhy/rbmUz8d89nUTIrDiFpPrymBVMF6wcq
ptpKwOntkiSz4PI/Fo6xTfFYIoIM5L1TVi+DJbyCJMsT7jNZ7saKJuspAW4paXwYJbFSEMHrjAOC
Njj70c52uUP6qECgZEUqO7x6s2/q1lN9439bm8Q+fAbSsDz3+oXCuCHY8X/zUOqv1Z3HQg+fol4H
v1CBg2BUfwrfkYBzbKZXcrjjwIRhz66n2EB0dmqGcMEXvOENdVWDgEMYZ1tcU9IWCQVAQWYLUhSY
cacdYy9yMZjzhmBCH+e+CR04oJ1NhLguvdqAAcxestUWSnDwxYbfaTpP3unSUgBDaow2YXYmq21e
hbq0kj5g51cOec38NdhqCvbimNX6s1CLfTFDxj67R6xSULjxhlFVYULhBZMSt/Wh9QVCPH8C/V5Y
tyTxyF6tAFKkYxragZ/sVzEOPWnCpL6a1iAjmp6W9Y1mABbCVzBELBBLVLT82eTsdfO2Vk/FY36B
y+mtrEM2DQ/BRdYCoc8dgiFVuOWfHfN7gl6glyxV0F2lNh2VksGKsT8ePUd7JT/vD2bamQYaUk6t
WKBZGFwV4vBMuUl4/jKxiMf60ZomLHhZK8YLZdTfQCcCwEoM1vnm/j9YnxVFqAF9I5ch2LSdGfOd
Yn70Z0kS3622KJHJFRLypCjC1BQPO3y5oQqsyqvP7Vm3VrI1Q8p56gJtJXo8Nl5PkrNBy37Dof5e
8ZA0o3kV7X9l+I6uJiJoSAyGMBtmj8VqZRXyH9X0MYk1QQ/H30GWl9rzinYi+qmk1PkRdrK9hcmt
K/yeUTut6gfbInyyrDd38l2KvoBKJvecOFV73bPLH7WXGY3JAJZ52LVkPoDzS2no+GNTGI4qLYqC
AxbWz3/WVT+Mv4gLatnAcJVNeXTwjhASHUkVEzVuRjBvnbGYJhQJ/Hus0dSl2xxFq07DwtYOL3Hg
z4oH3nmw1TdRBm6IDQ00PQ1nVIRezEbejOQ1zw1zVEKhp6n3an36yw53t5x2kUhB/tuhyvnsjzQU
BW2zPrTf9GFs4/A0+5q36kbjiOJgJdw5AFM3rrDO8XuDnd5StZ0NrjUTsneR/CWQL+Vs8i/iqG8b
K25afLbCL3fSLSa6x5Ucmdo2mQ+Z7rqpUiuzoZicjJ7pQC6WoOpnJYtgbcUVIWxnI6xom/U5KDHl
kzk2vqliChYFVRqsfxzjW/9ev/3rfeFzNpAePxPukeXEJelQB1p0hr3pQtbIfw4ZA9K31E7G2alH
2/2EfQbDKYSCq3fLL6/4Zj4wQbY/f0oJGVsq9hFtQGdB4YpaV+0KVbMnixk8RJRk+UX9mW64XJtr
bh5DBd8Hv6SmqrIWTgsM0IW7NuUwo/ARV5NqPIMrWL/E3q9b574JsX39YZWFBgqYRJJQNESWGf7Y
NsrKTOHGJdsL3B1vpJqF/G+N23tr8uD8ygX7LSMQ5axYCbildwdS3j4JkSFobUdhcyE569wD5mb3
0uG0u8YcWguFdB3gt+5709/F9jrsSfpOtdzzlpHe/cGztn7YNaZerFG/GirlhiUt4xRtqE94U1Sl
36Nv19w5J/oYMfEvwwcfZ5NbntjqD10ci486QQy1UPc0/T8FGFyr1xuBWpSoPVcO3GtjXxjO9cek
AcZslgEa9+l5VVZfOFhXtkXXUsIoqDS0tVq92hGK5rOJNl7Aawc9tzO+UGXh7K2zwlcz2p+wzg3W
7hzf6/KZ8MMUO7Yc0EO0PJc3U5RnzwPCfMu7v7Ki30jGWcW4cc064OVK3gxSqeYoPpNJXPVg3PlP
+Ndplt/S/7Llaw1Z735ASsnMulLd7QtnFfSagXv95MU6vxD3D9NnROyxI7gayqMvAdWfFPfm7kAs
qQXXu7G6L7YV5lU7ANZxZ1cLmW6h9Oo9YNklxQ+Nc8q28mSt7eHr0VCM23SWNBTWh8KuhJ8Fljwy
dsigvx/zvuRz+nKzgfAfCdygpWMTpFUSw5OZtiUfrhmhTAo/DiJS31WzDQ8jek2lEpsbvJUJXt9V
lCnwcm5/andeiuI9H+8hgojsoNDQpN31SC5TnwAx/aukU5wKMTYOwA8Fr3KKZtUI8TF8D4U+1kRi
EwcZYa/7eo7xgHbqBOZi7sEX9+Sr++h/L8uS/wbTMUVvPgnXM4lXUP9luFgv42heStwXlVBhoU1B
H0SBfH6RuXcagWUfY3H/R0PSk+45NJ3+VBBHnmkak6Mb5qrBXRQk7+3xFis68k+SGGJ1G+UOZYbj
TQeS6rxG7CVXvM7wMN2hiMA+tw5fHOh7hWQno9O6IFq3TSpVnBP3Zg60UsZ0TK7Xr9s6IBTMACUF
UOn0CXg3g4CPd69JcfnWofJWFuJ3paEUtNm7H+Md/m2XcjHWaFTjyVfd65NeIBmdPXcwpOD/LJf6
HLqwOo0LAON+LlINZ9Bz+9ftnzq93HIGFIF4Jix0uo9sS7xKBFYOtUgwFm54vGonxNE6dt46bup8
S+vmnsqyPu2Zenr0Wn6RnTcCXpuuccijyBth1plBBd98MsGWu7W06H1TeD5BOevnhmDy3fFKHsUm
0bfJqfi0uMPRA9DNGvYTHJjD88iR0LnIGV/2u1a2pTSJlVCRIPqYep8N+Yf2C+U3j7K1+sUrXdEt
e7OvvU+v1vQLTJEwNfAY2v1Th/8NRgQeeXnMDryaqTlIXCz/A+ItAAb6QdGy5BEpKnb/H+rLt0sZ
GgK9rYgZGlAlBhQr7SAHIBHIStQVwRL79rsKiWC8emRP5iXwyOGtHCZq4c2m3E8OO2vOmqlvJp8a
n9VPbReYZ9mS0e9P/ppyD09hryiMOb6MQOJe5gG+H8H1qrp2aBD274j9rV6c/EW0EsUwjqO0molv
2czqJE9KJ4DlU4vVmAgTJDvpD2dOOhqH2zVr/V492SDuUmiV8ib7FgUS61DJlnv7rAU2jwO0ANeb
tIGE1cjL4IZW3sTH8WrHFagVglF+9Icq/6DGeb2wBgRKtxKdK9hcd1uwNsHVU9GDJ3i/FT5QZGQ1
N6RK/CtvAnDtYHdqrJTOEJdAoSEK7a44+rDU5GRXWd3rtCOpNoUx3HXb10ZfXUjzG0sZIZG+l5lb
jQHMehPNOFkyWc00sr7IRFcYP3h2N9SLBE9461iR752p2n7hsxk0TVkTy3QO+3nDVTXnVc9QwJeS
XSTujz37lVTJEgyP9SrkmFBSjKDxt88sKyXP61bmkCK8Ggs2nAOCIZt1VqgX9BaLTE4rOuK3N63m
+AT7D7eMGfI2xCn54obcuk99jgRI71HRgjRynSX9oc06gNu/YRaXz0XPfhgyVS479FuXouEUvCR5
QPhSlCc/YoJJ/aM/mGJN7EHYaianhga2C3K4TLOba9DJH+bJ6qw3g39K+kNuSz0NXITzX/sq1fim
0Tz4IFJz1Snb0cDEZBByiXlX4YAI6ZMks07k72z11hUz1TygZZS2AI+hCoRW1QNiY+5gtT+S7asC
KYPF9vXtmvE+qqDfumOAz0v1YMH7aKG9WMou4IZJ8kymoqRSR7c9A6uboX2hYxH2bEoWRLPZ+0Zb
H5gAGgaHFLkm8bo4D6mvJKfKViIPUdgslzOcBzJ0FbudNiamaP/JZ/Sb2krhep8spZJ7XWY/Z+gh
uRT0uICJep3vUdeZACS/FusaZ2K5BLm3ntJ7AULF3Y+Y9nKlpzW1lAedAz8cSWTOyCPO9vu31lAd
QC4DzGwqxg8vQcEVurgPcNqY+JqQFsl5GOcCTJJxF28Wfkxq9TNdNh6qKMTkPppEZhCShMgglCzl
zlILNeom4lRvbIRDQW2PaXLIWFXWqe1Dle6h70TFLLKim3GIb5SaHbVkaTbaH2VbCEgjfOpo2rjN
gjosyeB9pCTM6lW4+Ypk/sDAjDqnBPWm0VygVi3E+b2oG4boBBdSBxL2zsuAFiqn3fQCu+9o/hgV
No+7sEZ59a4DkQ+2fmAunvgYw1ehIhCBF4bho0AMNUgr+U4/0tE/x7OJR7U7O186NazPY/BjuDrK
Felq+rqFK+MV7IhfUiRkpL2EHWqMvb3FZWwMkdoxGEgHSR1l8DJWi2Amx9FLi8m2G20Ql0bjvr93
dV8Y7M/559TMjI7+tX3i/sbOLvd+bZDOklQIzkzUWyCn2WD2eJnnHBT2L1HNSn8vdwuJuP8BocoG
D0zspulQXTTNyc/1Mly2pzvRG6RZYOF2k1388vbrTLdJILeKD/lYu8m90338H9A9H5ZI1nycXl1X
1HBChvOqHEwvjQMJeq2TKLeSLmRUuA6Q2ckiU03cia1GLu/37RtnRsGhUXLSoRR2CyrIbUAyOtyf
qSIEgZnyK9S17H6XCBBcOGA4CSg+7xx2bY1ESBXMxiepHzwZlkQor7xCFuCrpqAaB5zNCObaJ1eg
gtzXP1YtxMvHnzTZoAcxfpuKqFyN8i1ooDYxlLEx9LA6HUJI6gl89Sc6BYtt7OeXc8HV52OAZk0C
YlcHZWQUpz4rjzQmMsBsxqoqM+ziX7B9jV3cul5NvucHAiCMQa/iyKkbXTpcurvKT9mF9WCcqJqw
WiYeqHuxzNKrCJO6Pam2PJnzgCDvzRz7S5mKFhrwRDgVgqW5SVcsa0pFMBv9rtgGmhteV/d3SSkw
n+dN9cxm2mcm3LQf5OeOnCUEvHc2M2afYPN/X5JkIeEO2G8DRO8OxHHZTn1aUkqBnErs1HhBhMgE
agEi8CCOIDosrgjncGk28V9cIrSfVkPoLpv2s4gD7w69OO9CEq1YOww+PevaykiNbEK5wRLAoBs5
7WSBRc3/izG9gKh5sxnXvL26IyidmOMEGp6WhS1VFIborfS8JmGY/Sw1rRY2g1vUa3/MGyGv485v
D6BHeGSvGigiuabMDy9i6B+AJ0m5WMbAKMuaeWezW0kktAXuydNUkPq97b+4rHzwKLgjrHdrMriK
GWnFYD9YifrOSYPx/SYFB4a2qj/5fQVmdApanFCRJL/VTuqYQPAV44ihsAcu0oirWIwm2u9rm9vX
1ONJe3y+idDJXeiINEPdXp9YW+NFc7NYM1CM3szErbxNfXjTCtHG0ScfMfYgH4FYcKlc+hjkCPwB
X43CGCdhlO64bLzv8lT4zhFqA6/vdhE6wAv47UIG90RqmqUaC+mX1PAtLIih/Elm1Ae+lgvEALcc
pDmdKoxU4w3N0K1lYYQY2RSHawK5HxVnuPBwrWlQgG6hRpslrzB794egx2CQ/eyjQJuHmBL3RijD
MSb2W2p83qD/0RByzzzub54gtjDUmxWvYeUyx4Tybs9o1pJ6BBysv3i9xNC7f7PXRbMyfj2YzLPN
ZSv4ujMPGOJxCpNpA/XcAbhfUQGpsHLq8fLmP1dYfZyT3Hdsp4LOjUq0GXF3xK1DICwJIbbFY2+H
PveS6splvNwI4AIt1hY4J1R1BEE7LgzbPyhiEP7gc/3sqzocG7yyNmG69Y/qYLDFNA5Kgu6VwV38
7RiGRRyw5F+8C1F5HSdk+et/5cX/JpmWYK3YcGxAWVju98punW+voRWXV9Eoz3cGkOY0GM9X83qg
/6oxv0I1ak3Min1rFty9WvKufAFzOQHirchOrl2LGsjYZnGedIcOkgXBc2B+xA0b29+hXJRAeCbS
xkjX6QyHtkpYsgrPjZwVs3aXUHXLwo5yo8scjQUZNdDHtd181u9e+9nkCxgMKQBHs7pzquv+No3O
Ooge8SzKbLVk3Cuu4vzccZmrYbtTv0oabXpFSzDZMJXwIWgTidr0QiuQbzWo9zyha+DMJWGynh6T
AHD6KpqaBWePz5hYwXxHGq/vBU2u8NIVprnr/jAKLT3z0L89665mRKAFDePqOrS1qmDPDDrGOHBO
Dn12QilQpnclSP/dQ+2PdMxDneklYoq7EvPviMczafvyzhBuEpDUtQZnAKTlsTNoBKUjaqYbn86V
JX75z61Ve/90SwpP+DIdZhQR9cKDQjYaYej6JscnlyyIW5RKo+RhgCok2aXzWfK9sWvZ2apU1a/m
TMHF0pjA9RXyQjWOMPXMxWCusxhTSBddu3QJzHF3ketRMewK3/57sKSr7VUXPd8vLT1fi5UL9LFK
4vtuhyGqTjcsjWq5fJIuPkREkHJ0Da9EaS0SLvmPDlTQpuk3xwfX8B+U5IIZjhDWDuh3mWHWmCt1
EY2QlvrQuvDQrTdAvOntWAR6I9kHRNN+dmyAwqWR0OVePi7M4Xywwe2jNFdxHjLR+mOiS4nhPXSU
k9MjVfLMgKBPuP+WzF3CfAjgS4j9wnVeDQRfDeOc1Fm/IjpXs9JkENqTNfujMj1DmVpjAx9lOGOu
02uuFmgoPknqZEAXJAoLoSbMYr7b4ZTrRUQ64ytxPIY1F7ER0XxkLDBzMGPJsF4aDGfDQ+IYG6UD
5UOIU+lmvjaw9/kSq1VxHF9FjNXK9DUIUI++3A9IAsbvCLrxNJe8KOSZQ00mW4mk8mbKO29EGOu4
UlG0F4gHIfszOARJHjkpHOjkcAFu++SWbw3kgLKIRA2YD7xCYQLqBB9iEvoHLVV768pIt+YbSlsn
sjIa++VVma9pYSV0sSxwIByT1lRaA2P3hpBBo+4lF22i/6ksjzx1n1jPku6b7CuUi1sKHdP/k0Bo
IK/H+PziJJMRDJ4eY+UfuFXJ/XACV0KsCAk6v0X5ZnktMHZi7kWCr54RxGIDDVpw4xWwJAPRrSuR
jpZFnUmPN4R/yxHagwtBMRXzy0gOxDWvPxrrdhmXQHv5rfC0e0NMijPNkGCaIh9SWwY1KdjkGz6E
LgsTDtix005dm7mpNCDGM5H4n9g/7ZX8QPpZaSXVU+b6ZzaRwnrG55A1kaP4fvZeFYnqT/vdrW2a
bGlJXX8nj5xsWkaYQrQdwXJaoDRmdvBfI5TGh2fuEeI9r5HvF4fxjpwwQznPybnx4xF3somzmvxM
QYtV6hc7HGRACZgJNu5KwRWFlj9UoFnUULPKkseXGw2dAZs1NIg+2QkrGxGlwopUJatrJIxl1ZaW
EydO42kPz5+gRBpc74aRQF701luV9SCPUEFIyfQpjIfHIWO5aIpV3CyouXI/JN/MFtE9oH9P2/mM
4lKtkqHTrtLTfczD2Om3h8VkGGyx31a7/gqT4IITr3bF5854R7LNNXmPDlhnKuXYdkeaKM2NSBx5
DKJjEjHmk3sGf0ynRllGFXcFhRaWGY9ww829tUTgJi+RjjIFhtR85beJ8AFDPe+mITeF9RHTeoKU
OdGxzX1bu3UAWmgTN9GtSpwxxrgbtPJb3HoeSuBsbaOtnKOgPMICnZ7DkC7cLIsBCmNzJtOZkKJ7
vTiHBYVI61fnjrDwysAtgtoqFa1Q9BZUQQmnPiYmWHqWGGmrVJui2kP2hnfI/tKCKa4fZSzHWFEk
J9+uZKCBmGhXvRHfD/xh8PPmTabrRTCLjv+vLszHRj5RgsDHeTj8ff+w73x4kHvzSbSuIqdMEqk1
A3tX1RGl8UFYPuMSQejel7yw6fZiOVjPdPgXtkzxKQ/punfYZZmUWk8m+B3IBQKA4CG3wpW8FWEE
leNReYuu00AC4GBjY610CnHD68Tqhc/5IcEaqke8CnAxoUAUdnSQkXj1WpJInZroiv81jftoULcz
GVMLKcmJk1ed72+9iOekwIdN9O9GB4+rMZMp26NJauH7UAIc1IWYjY/+jGhTk00N7woW3wc8GXEL
GA9PSkSuV1lBWxFNYckf1tDgtdDf2ZLRRVCjEm+Gbo06VYG+e/In5pgYinpdudcpXuoImQjFhmmn
t0nAHzPnkHJhPfEEJJcR6mYImi/2YYbDVbl3kYn8nSFmLf8DXlR9CIzCgeGThZoOScsyh4bGciYN
XyTTWxRjLVF+kanjWVSi6vSVe4cdFLVsGqlB9G2cmS9ypjaHBZ8BczbS7uQyJRcTHezxWnHPraQ8
rRN2xge816c4FHGrL/jOvN1bCIBFJxQH8OlmdUeuP8rojWApBLOyCDtmnsq5ARSoELRN6/S5kfQV
3MHYU0vyYwBn6gYKIdgOjEnbHn22cF3SAQOzC7dlXnmHY721aRdH8bkD4TzYP+m359TQJv6E8IwF
HT4J30UeSkLYPA8gahgqLlyd6pWwsU4gpAciLN1JUCX9TkZ9td9z22u3c3kHqdO12F5fjR4k6ImR
EpnS99BV4PNzQ9nrdSKLDS9AnY8U3pxwrVb11BItiIlwNP96hll3/Bc5AP6MuloVwZo9gU9Ni9ou
DJiPM/msaFPyzq/9eBr29l/ht4LvMN9vUu5Xl+Sjbl46bYesHakXw7QCidJM2O3oHUQrQGwelukL
Nr6xn8F2p1+sIY2tVB1cXnDbboLxMju3Mwa90+8h/SVTnR95t+aLb3EU330NpP4fh6FSA2x+A8rr
/NnwVx+32kzYpHVExSWRnD7IrA+NsZnFPvwrIqSmE0l3poTxKWIk4g4rHZBen/BzI2Iw39kcUm+f
4SQfQK6gRboNWVl/kps+rQgxpDjOEIfeVbqMlZCzpBOaLKF6t49yzDlceWw3Hw7/Kst63o54IqhC
7sXOTu27fmyrMppcgoqf4/X+tijOZ7vUMST1d6fdCZ4prVn0oiFftSqOxScdSBDI+h2jbscQE4EF
CZL+A4OtJ4V78UGKfEtEHyhJixJXBdT+ZOBWPw5s6OELzJXDEkb5ZhNesPkZZgutaM1oNHd9HAlr
V1VlddTOC+p0WY0RLIVHKbYWTNkwjXpHofYtzpssh8SjT3fpyDIZzszLFDQToSgdLJllGnCKJ9mn
EW7aMsG6j4renLIcM/+36soBqwx+9Du9vmgBvEyiLm+OFSI6QeIsvB16AP1IFMW5xAhc4S1mjMY/
pMqguz77t1DkNkY5f2ntrqH62IIWZJ5tvIsf0uEOOnqCt0STLV/pv3rAE3JkZtWnFCGNdO/GEIhJ
z7FFYg+W5azaHfiQgTgqwrxsxp7rM9XOKxmkYg+LHZDrP84OpWQAfBVQfQClRflYRX1fkeOBuLMH
SqzkMA5bRMaNgyZaUdu457lzDlXstI5+IiZb7Nyu2yLIobImtDvaY93BPQDixZg/+k9zAoJF6XHE
Uw/qSkFQ1VCAwGr0uLJ5sgl2YPoYBozeOl5hyWRahgTbq+i8VPRxXvFijSP8vCiuPu+7/wM29XL/
6TqOCDaXmDZ4pnQ0e+3Dte15FWHM2bUPWRqeZbt6z2oIV1ibY1PHL+cPVoHeSAsDGxCEAltvWiHg
Loc/l0XuoqL4hks0B/+lISFh6a/MUg90VE6PE6kC/O7xmZTMefjgpbOtdqickr3xjbpPK3mFgemO
240psdAARwaYaN8gn835DcxGjqt/CU8cPm0oETf+NqKdtz2L799UF3Rn178sk83+Qd1ouDADwKHW
MWR3M5/EQR9YKU3bkBopKMtv6LAD7A9hQBKysQ1aYYZIA8aoTls5+97ne3JlscmqmHlTD57QSePj
KAdxlHWajQgdIHVYs8TWwOFBAj/uTVrLNtjR5doFbCsnHj6/R0bu9/u90z2mK+115v3WDfjDGLfP
+My0l4nKVee/66Cgei2Cb8VeOBlaDXQ/xFClyAknyifdSMB8k+xFG7GRvyyY7hNA55PhTLkGW+rN
G1uHJUMMxdhEZnQywWHIBNAUX1BYADmEWaM9pqHUOA0AdfCYxF3A4t65clmIjix1EbByWS0tiirE
62V/q0q6dPLa5wNNjMgH8CDFZwOwDq7l+nqPE5AocF440xxZO0EgA+ksjuN0jarJQ/mcHhs93jkL
ySsipcOi3rb5/Bi6OH40t0j3K25pkTUYmLmRG2qVlf7ZKX+HjW/v5+sz4PH9JHL+iz5U7X8+Evu2
7bRCvMPtz8UE2NJxqEPHy02fEMlM+jVbUlW25kASBr7V7J7nHs6p9BGmshjQ3IIFz0GzEWP2DS/k
ykmsFYTAl3lhQmQqcETp6yIL5xA2sBoy2pSzSxUIjujcvGi6Y99GykEC2MXb6UkLNZDUvVt5wIvB
eQaov8VArCOTvFIjqw0zOR5QXrk3JQXgc/HgHIiHNjiOt/RF4VTAHbxWnznWqtcF4T+rvXtD4YwW
0QclKwc7xypUNriB0JVDVgolKUoqHhh/cSF3MkzfN1bTDyauenvI8MND23GMMTtsc6RWcRCvcXYy
WWmMLbdQ7gCmbnto09z5/lni3qYXWrUf4BHLEAtY/cK8YCAiy2qQiQcXbO5/ShVXOZtVuGb8dvXd
uLQ2UoQuTgl3I9AzSk7cipbmo2Xn2loU1kPm+KECk2Tokh+h/iWvpO5wLj/WErLYwhTtHWXMgT87
Q1QHj7/MTQxKnFt5L4PSkOcNGD49z9JMtHFINBTRN8zk2RnwvKchwZpx/IuwZ+aT4pdwQLceRDeI
s9QOwdbFmsFT/8Jda4N3MYl7emlbecM+yxUzzJSdeNa0n6XAlNfJqCCFpGBatEivjv4xnu3TbiTV
fbPkqf0oYqZzJJ6FCB76QTEP4oH5wZf/IPmWXAhvolE2dGBMj7xiSre/gC1b6YMLvgROCMHBn5CK
+7JUJDUf0a1EdODV3fsH+XMjl5xMw/8t4/cmdUbDh+VCSGWEA/g+6uT/j+CuAfORLP2GcLWysfmC
2HgspNZZjFI1yGvFMDsWQLfdCggw5f+FoVKeGztKopPRVHjOAiqlctUFlRNiiQ6HL6UiR27OSJbS
oZr+bwpYorerkHpetriP8z8GIB4O4vdR/qQtHfGHFZDMMjHxtDSvLcD6NeUUs96o2UrAIwwgUSo6
+amaSC2tiiWYd/3JkDJgpJv+AH6WS0Fo2PBVBNsi5L/O+g0iL5JOQt6xsCB/omGS65JnH1L/lYOk
LG11V+StFEC/i8qmI1xIrLNtIxQbnZxdWfsA3yXsZiwNVDyDux8euDiamrS1OGkvJ+BFJ/EMEScb
csRTgto7cPNK0rZ449YNup7NmJu9/40zQOb3y8yKXByS1v5RcK4Y46ecq32uWE+FeayKki0MxNWv
Jb1QBdtFxjXzipLuguPpBvAp96g3WphYGLUaTP18LvO0PCYINUZqYfK7hJcZPQTcQiTPWIesHEAy
gb6/V4NSCT6n586ydG2oaJYn+GLCutNfEhH0Mqy9nP0sDEb1SCA9ZFobbO6XAIezjKr5Sd98k2zp
1kV3Hd4qgvk9P3ZxDwi2xtGGo8kwy3RBZUZEK7oZ+LVvlBjbn4V+d1JL5Ps+PSPTgeiK6Zj+HbHv
0aBKNRT7wKVd9n1tSaM2VyDewLCT8Xpn7Sp7gsYf3/xA31WH1mi8ZS9GqlKRnqejk9kNYzmx8pET
J3dRtPjwRYXlEG65YRExUlUiL6yjZqnLNrdG0/xQsYvCqMeiy7rrGHvt8sj6zlE6FPUiCCfIGchc
Az1jDMyqsf63TvefpKYc49e6tjlPkzSEPwvUMYrPHS//NRrqwEceGqSoQ+c9VU02M8/BdEuOm0Er
jBt4apw9V67t9CVcPuPjkqGxJAqXglYQbj2R28c1rgxmSNws8vLdtls3SFGAZT8BJHPwIUaGiHzS
/nHspPbDB+zw5NPCSCpYsuOAut8qNIMxl+DXIiTt3swR9FLKvdFcsi1vXNazapKLRd80/KXFXwIe
OtZGlp4Qq6KbsltUAsy/F4YShMVFq+f4th9tZZ3wCzLyeaFYVmjUaZ5pBnptNoQqVSgRM6TYzPDA
UnqpGXdNLlu+Z+VXBpWYgguLEztlR+tvq2hOc2Itp0Hi2WYAq2Mj5uo8c9AysorXa4WnsobG5NXr
2+UqrDIcxewVWjiEjfMSAjwzh5PxttCAENdBcWFi04tTZt4Gq+UOurFvYpTZCzzybK94K2ZgQnGV
+0ayIEaNJliohUlqxk3SiYiE8emV6uesulD5ijCj6390LRHq80Cus7GPwYNOt4NGfVLqLLZRVv/S
l+xB13iG+DaqnfXycKjr3aFa1r+9lOxq/M/4/SKWvGKe+3qS5cLeqGNabs7EQtWKwV8zWKG8CvrS
eakimZavan+nSR09tNyAjn+GoX68d4tKIfIDQp7OG4vHP090uII4lODwrsQZSMPz3vNax5FQQYRS
Z9eTZPWb4WhJxMLl+dQs2QVJJOAiPG5ZXhfxC+ktAEK27sWeGQA0YsDAzlCRDlaOOtdLRLGq5m5n
dFR4ua0tVdg8OTHmUPTn4cUo3Hs2Ktv0LMlUJLfFW2RzU2Kj2Hw+cKjhhpnYyyPjUY6g0fx5S/+O
m77DFO1c9TvXqlHSQV8rd9bhvQulpSjK098eYthL97St6gMu0ldpkmJmwqN2jXbojhWlolV2EBlc
YQ7xANkoIyN6OzIwY5XGSub6AQeDrF0YZsSMBePwolXc0s4ttr9dVjOuTLsJ06j/Clk53rc7bJBx
XDdJUIyUYyxsbnIx1E6W2KVrLPAS2T8MXj12Dz9O/EsSNKsVXIvRN7+aZvLQjKgGjOImGUQp5o7q
/tVStqeJx3HMmoSQn7dlKyjqmFfzP5xpFn0ar4hEGOxuSFNPaYuJb/6r5QyNqPAm87JRKLvgiGM1
40aGJBrOMegvCJlDualLvnB7qPxRYkK2hZFnF790r9cAOETpq+e5sTj2Cbm0Oian2nS2DaMhTWbl
+/dduA9KrEACZx45XWHzZGg8Iyqn7PKXWvjfT6HjOryNFZBmx5Fb7/SEHQe2RbiRtGS/e0kxFLQe
uVLw4Yc74alJdWMek7vZFEXDwkvf+94LE9aU9FFRYlqxlMRdyYuL+oT0xfpNFk7EXEJfYfnK9GgV
oEPr7jTG0WPydGhfudRHAdWUqQBi1+QISTgcsx+UEUBja3dh4EN4r74S9KMU92lIZvg7NCshFNMR
5ACxUJModTdJP7nhK7CLgVmFP3sFgRFpISH+th4sNO8yD34+cuKN6/hH7JLCE+GfbB3Rdb+CdgOw
Lp1kARg5uCaoTHAtGmGNyE3z3RJq3DLu/zhPn7WIY7I6LorINl3ROmVxZN2rdKfjCSfLhx8Kb5lC
nyCrr2yd8RchL8E0PqcE7b5Z2iZISduzAHX2OByQrSRH1PPIrrcL3FVe1nTPNdCFtppjfXBZyvEe
9uQpHVTAri8cum74ZE7FnW6uJeeYDb9uA5XK5nKm37L622kyx3haAa5wUpTOs4BrPIBebg4QJf3G
+ndPaxjlGwuhjP5EzqHP6QqwPTo1kW2GGL2GZBmL2ABBeKDcVtuU30nr1f3VvLuRoMPPC0Se9tjK
pzsbobSDxHjCLCnr4L036TeNvXiXfko6Zcu5VbknV2hkDDXDuRyxzk5kr6oRpA3jqMG5uhSudFrs
p3QKbKExy6PT2bi4MpTY7LYjqaMZSPRcrKxfXNKuBlwWXVhCt6+ifzEFpwacgnWaIhYzs12jF8bl
gx2w98Dbo7Bngo7021Ogc1NUQPSHFrLdop1TL35rRWduTuqH7y8GlRM/jLdUfWJ1uqzl8UsawH+F
qg/3PXiDGlvVAwK+vJQqsjherSDukVM0KvCKwdTRAsy9eVkFoqAuvlKMAV8Y+Sh1o/syrgXD+VxO
nmgIaoG7DJwR+Mu2XIXez5tayy5mp5YduijFLN43JRTAjI2YhJojCQAk4tzLxmYiUgTlGzaE5YqU
Q8YKVRNffYPJYDlMy0vCJSMFI8myIvHLZSZok/M7aJqtUQr5CxdVHVxabzQx+MyjbE3RDaP5yZud
KPGenHlBjw4Pm5497LvYlwJuS18qvHWtewGJgPxexWakvFPkUXbw15Pqyc8LtJHFYQU43jqsTY6Y
x3dHP0HKQ1jC8sLUIKcnOG78/FxKfFnfOxEA28YGakXe8YoT4bmT7abFX9IXSqw0d7EG0pZfIrFg
NnOJ0xvYNhgv3iqXtN8RVv2du1FCzfotMedsSGDrr+n9H6kYs4vcaNloAALwZN7U0mOkC1Omu79D
20nvAAQj0F1VO/TCvK1cZ7AfC0d+7CSv8K+Rj9tsCR+pwpQ8Dun5mKKPArsEE1emB0pK81HMPYtM
GHvvoOib4me7Lsr0llEmPlKcYxh7mkf79iZ9SOSuPHx3wIo+z3JFIfBMDYN12WVwkvHrIwdnvu3t
f95wU3WNKHvN7zQ/yM2IN47RRCh87Nh64jPU/rOaEoy/KLGGg8Ql9/mVGUjqwgQ9oGMDU5O+PaKV
K5gvI3LDAJYxImP0imaZwM1k2UcINJjQBPAToso6sP+9Gg/43ov3fCjlh24nMufFYGuFOdZKESmT
0+XYiui3t+HE7uk1KwWSFehhGExBhd/j/zSGhcMY7plPuYRiYEBc4gOp7+geZInT9fPbCY5Z48z3
YPvLKw+ltyCogHVaMxojWBOjXvejIYYJaEItIabnK5NVYaEEGfv3snFbdUghdc+E/LoqseS32AEJ
HsgIojJeRdKF08q/zIvnOMatpwC8f+RQwXa8hvuO/Wkiln1o+/cd3J6FCqoM+NELQRALXkrws+jP
dgVPoSU+9wUqS+frTFwPv6bIUB5D38HSzzKWbfYZXtplNDUT30EadvjZmETWbPXD6Pt2dT/15suE
DmMmU54qX1HRhkwGycRRr8K7hdcQho/7SZTpDZ4nngxIjdj4mQ07k+hR/wYSxEButzLwJQIRWSOv
54DYmOlUzEpGzobrjDFEdq1CfbarVZDF4oE5/6SNuMcpcn3ogPNVvz+DR4Cx7rbmGMfM3b36No5X
k5EQJDOCQEtm1vbIkiRLzOIZ795OxpqJPiHyodz5gPBv0/ARSQ85k8Ar/+7iSalFJje/eUSRrQNE
zawDyMoxnVtjnONcfqxxZ4hqk2XoGxt2RvOYBzqiGfxCQnQSi2nSuDky7d/Xr5ceR4MyVcvWcXMK
SyASVZe7QkrmZ2JZ/rN9mdSeektbadkS2tXKxZar+vDcj/CbLJZ/eiwMgMMfyg/AGeYogTEXr1lf
xsBPvyKulWpggDpMqyASxsjWf4tD7PfrkzBl0sFHFZ3BJFabRLcmDZN6pvraWpyuGvwczarFKoPt
R72yM8hemwFt9t+X8FQsSQlr3G5jsbmknSUMkrhAYe+71OubYVuS2V6spZ96wi+RnUKkVM8+DHb6
YADATwAx0kGuZZqJ7PBuGX5dRCjWz1qD6CSGvUbOZXW2YJrWr6T3KXH+cT12LuZXAdlPEaDiLJub
QHg/1S2tG5aSZ8xUB0vRYh9LCX6uC1KGpeBXG4QhU9HxmSKlnuxeA2CvsDrJzFwxFKTfYx+fmnGT
LZ7tCydwANKyoNk+d9vwd96U7cJC7CEH4OJ42WSt1Z3Do9Jcp/nazFXh3bnALIexbW/X+xQNWnZp
XIgB3+JXCXOInUZ/vXwDVsC02J5/ddI1JW3NED4uK+u6VerSIvhAuEcG/NJUdQCpj+PgbDXTQNQp
JSp3DuO5U28aIIysM8rwxP+wkQFeVTNXDUtVtu1/FvB5piBYrgClaPTvFKQ+ox9UnFWl/DDvpnVZ
iG4VqZgPZEmHnT6NEDyyPK5kXrnC0wb1ctNkYHuPpsnrTC7mixg236046M48e27oWeJoTbSEwSFf
7qX7RDL2aWl2y0Nhs3ASiGP3cvfGbwuJGCRgifIc7V9A39WHLMK2OJuUMhTEcU/pbl04lFh/uUpL
bSYdBzy5Yo7gLPdaAAODsidoArRskYdHhJp0PeiOAqKAmvVc8CRF71htwjgSWuUv6IiIpGUiKme9
FPip5m9QzOjYPBwsi9hjI5aLNyCPlWWUk/LrXVlwIiXsjw0lTfSMMUMAvav8LCXz5ybz8pigW270
qXXwMM+LFTDtaza+bbEameWpyJOKcCqR7Eb72AgEMwBA1zfk/lg7S2Y5ax5uVwQCigJEF9DXuFyS
FlDTw/0zTAceMrNUCIo9cO+YhGSik6sSgkRPJIGRX8sFwuomCrS6Cf/aLQggRee+hKmpERtBI1Oi
CHgt5+hnzExc/T5AucfgwURc+mvFSxgotepCvK+sCSJDDO4Q1G52NcqsKqAHnRVc+hXmGft9rCXW
obACMHgnhmH4iJOTWnoABAmnQh3ToBoMgSwVodbLe0zDCaXWiwPtN5MjYByDuGTMNcuWPNxh4eBM
wkjtz2ZAJsU0dQgwE7fUqG3NZHN/Urm4wWGlRPJtBw0TyLoaDfDjE74bzgxFCW4fH/2U2KkxlsLe
rfNdU0BymM8lzed/eDcgZZf8lMD3mWV6izgZQVKkzw3WqEmJ4d4eiMbCyw5BcC1GyciO1raNlMsA
XbEFQgyrByNwab3Yq84yz+IU9qEzhwHcAHjgaM6pD5gHL5dkl4qWUCXcSimf0iZ+Rug166/pPYHW
9dU5aH31XRi19e1dGLkH86osweKNtQaTqKCaYvvP0NmDP6ABq0ssmgexmjzrDL4wpOZKkVXFfmMt
HXF50uyJqdeZNo+hYaCBixWuNjl4qzmFeDhxjwOOb6UpAtO1OggDXxNiFiplr7AwERe7C7QY2rFA
9nricY/MteVKJ0L+eZ03r4+kwmBGvxrhOetvFI/L2ZFLkUehecdXWaYGmwue3QYXjSsWX7DtdYg9
8JaIaTahL428b8xeA7JuZxDxxkwTjCtju4DC9h2fyrR3l87PvZysLLjvqZMDz7Ma+BLIfQA1bH8E
wMr5GUGE/bb3cceXn1s8pWis9lrCwVNVNcKOS7MrYkMGkoeeoiwIBPUUo2xuXSvM6vaSaIktSB55
5LvPFD32Lq1vuRaglFJTBVBUAo6ODzptASW8m5hWYag3o15LNoMSF9z7wOwzKX1CxQ5XSBeU/iJc
rXkvJF4qk9wWhPbxlIasHqAhKyo2Ya/DIV2ZlmX2oW6nUR8vf/uhX0qs1Xip+nFVZosfMmBn2+k9
4f5Y/uVRz69S4dP+gHQL7JEfTjAs5z+NtE8+MEkV9tTvS5pXIagOACBelvVZOWQ6Jf1Kg0gLFjAA
QPvDAOfSrm0degdfzrunRC880VxmcSBOPXL5VtUkmHNyMaT0WHBGCFpyl+UtdjuUSoNyQHgc4dGI
q+8FTuvooYSFI0O083gd4D0fKRziBgdxqxaMjruc6BTMrM7sGHIcolDtmwGSZxfTJ1JRn9WXSKvu
EX0IAbYBO4T0uiQbo+fDh6DjoYvABLIvPWxpj1KQA8ua1arMgrwg+ULu2VmC2i+JQ/7aVhnNaUHy
9ggeI5nIsCXySLrcDoDGuDe3IRUh/a1YU6ZGzDnBdWOHG60EkRwRRKhmCaeetOapDqAuHQaOx9tX
oH8NKPzFQ8llIPWbSKmGW7Iqyia4xhfDl69N4FVhTJtR3aUn+CLzynFvGttP4DWlpVVXdbeBOsa4
BElk+dr4FiI6WPXlsiLVPnVJEdmzpyTAO4W0WFvV5ojBnvEUHPXYybYCThsWhZOLELsxPIfqCu1P
6q9V4r/mzvx2p7yTdslk/JFS0lurvzio5r5iI9z6uRJXQAhPao76nv3ir+1aeSpxxntFhn/Efr2q
oZ1YCIb4tqbOlpr1nSFbHYrUxAw6K1XkC/y0JZHe2EIIp/84Zugdmup8U6jOjIjEHB8Q+XCuxa6/
Bx/9TqeMXs8jd9ji/cOHUipXror1j46C0L6dCLj8b/2rFpK5A1/NPibETElBnnOAIzU0V3DbyYjB
fIpIzQFBgWRlXQZHRrpCUTpop+Jz1L1YVSxWUcBvduqr05vjdEWo2Ei18erX5nmiuOhBND+4JECl
UNza660nUGRCwphIIiMdc5q0IYIdUkbrWYHYcaxCzQ7lrl9mHttDajuST1zJv/9sI27xKVzYFIfU
hPOATcKuZFIFl/FLYYeKa2bXhu9qzHMhw4gge6ashgbPYIYyH4/udr/54yd7Wv0PxCnt8nqRH0Su
sVVLSmDSpg/iAD436g71zeCAW3HIRpbiJygAdNKXOGq+dFWVU8sfwzNBNo8qr/XS+qIwwXg5rgt1
aP5pmzUMNc60pX5GRHnDQ6FjWuQcrHz88AJpRXmrEqb+0JCUFKDYWFicULGLXPFW17r6nA8l6YU7
q7u+sB3mm11GYcSIiS7DDek6LKnrVuFPC9LoRr4YJDml/uTbuGL2xTRiu+VuuhGnjJALJ7w4pVP7
NNzWzmjNH6JECy0o9uCdXpvLu81tqSK4kXyCmPYvWCdLxl8WgwXv9g4YCQ/mp/CFxt0wkPmjQ44z
ALUjwPjF+ZJllk/m6y0lZLDq7/MOMDNzZ4+wiOjHbMOA/eHG3IklEPyKa30LVRPozepcr9jiL/XL
emTFnvlUjyXWWzTlMw7D2YMXZY//J3Kju7bcbdInJo+n5S2hlzagFpU8ukvSBAYzFFd4fgutFLCl
Exw0zxwoKway7Mv9J64vBx15JboN5VIQ60h37tLzWEsr3g0omj19dj4c0eEECvxZM8dpLuWgxeZi
Cvm2zdH27o9dI28p+0MQ75PyPn6jnfI4hkIXQ3+5mXuILvmLX7fn7Z8rAdz73+QV31KtRIu+4rzb
FXGJ6aXFngk31vImX8uVcxY6qHEou2fAjcQGLeqAWANyROoaXvxCVxL45TA9rt/MRVX3pWX9RetO
yTySJA6dHFMsnan6g8DJMfTlsbZEkgLt6kyXqbdUlZWPwQwRuUbqGAY5WVtKG6q+6Rs3ScsqX7rU
2HuiMzMAoRR3Be5rfRbrcHmMcxFp8H1qm+frEAlI2mQ346ui7lFyJuctd7XFkvrWEes0LavNOv5J
NfVZFyxfmtNZH0ApArOvzAiNp4mVR41X9QXK2uBpY6IfTr8mc5gekgGxvH6wvq2xUFODmofKGjOR
VlVtyZ57MMm1YmutuS/TDjuEQZYTxAslQWgMvPKrTmGPwDEshy0Ci5AOnpb6skrlyziGwC+jDut4
ziBed9QIGTRpU9/KUYyOYk+KvTLuJvYb1RpXnSI/GjK1HbifRsuFdecMLfV8cqchEa5a/x2DFp4M
kEIoa/5roMpsQiuKZO8IqiSpvJjGvajN6COd+ggP9uZ9/SaJpJaz1NhDLtui+XM0lB65uVVtO4cj
usBf/UijVOZuD3br5Cip46kq0NncNq5605p05SbKTSWRJ6YhhLgbsK56eOPKsnpJe3B0ncOJs1Xo
2XdZGr4iQmLe1D8bJnKGid3z1EZmd/4rJq/FXWQXFvjjhCR58c8AI7ZpT0/DZRklFVBadn3im/5j
et8QLVjPBkEwe8sn1xbGidnQGGMdhnICrKhhsxDd0IkM9T9cmHlgToNEBo6U00iGVecYrHy0/8FI
fdRkwzh34H+Y8PG4+irxMkbYShc3q/o/KVkyOhANU4Vt9ivyrKBgokjj2mlJRGKl/tHdeqdDBDQE
pLNH3EIoKymH1vYtxmqcZgvCcKPa87uSYsscgbgsk/8ZBJ463h3L7kCrm7oogQQPMoetQH11OJkN
C2yJy7ZFyojji+2XmtPzTw8nsxLO8F90NCP74fBM7vmNhLQbq+IkjSpVU7nOjW6Zn5wj+4kLHGeP
VJgQIDytr6ZU1B1wk48iOH2MH5OBmtobJjajz7VX0sQHULWpYJzj9cgjtclLckKPNBGDkYqL5ZTS
lJUzRHgzg55qvLgeirvg9VQRkxLVCAPnVjb0F4r/RKPkq+IVZM7T4B2m7ysarDJwrJYvAPHa3fSm
2jwr803kg9sbYxU0LmGl8mEWqeOvdzS7rKclHhrVZU3+DdOXXA/3NJQ05+DvsA5oeA2A32Cp2thw
DsGqImOXWU5xsMXL+d5oAk/Phqm6E1nRwYxGvA723KCGz7dWDFUK0yzBqhqVHaiwKse3ygaLx6Kd
662bUchjX5H2g/IrKpr5fkrv5h7Xg2tlH05JMy3uUbi+h7V3PJ7nWAlthE4dgxtB9zlDBS4t8Wzu
TGDJ6PeTMFogkiUHNR8xjg0EN6jGDNS7CoJF8oaY+sUeJjAKWZNLsPM9wHxM2xBlUT8lSVS0/maO
tJKLqUMhzQgsaVw+ov7vl8wkMxPIf3ojNwMMTjHroaOGcqXjfJ6+NJWxaYlWXR2nzoaSVuywUggI
BvhoAE2EUIo07auC0xyjw8o2njXFINnbGYW81eYgzq+QFi9wbu+oLxWYC5gYsID0ynBbzartpFny
u2us8tuflGgxw7zo0pzcIoq196ItjclIPP2Pp9kE4X3wKTgU8QPjDXclfMZUAy4gwj8s/MNpX7Bj
YQlOqEcd/sFJW0r3pPMMsU+OZU+1Po1S1Q0vbOxVjYzwzgdP2Weke1seq8ZaovPlqS9SkYL9mQ0N
lsFOHN9zBCrCCzN83Sw+PjQqfbk5GDWOkBk8qjiRkzxxQO3A6+vWkezo6UOudKHnjaYth4AyQuvT
XEhOQgwcec3sLddWUuQuAWF2Y2N24UahkLFsXB1ndeohtEQuhAOTjkZn6+goA9pTHAClxNhZHSR9
0/Jco8XxrQ8xd6P+7fNEm9iIy5ez4Kp7NDr0knVGekc36mlGHDsSNwyWClfITiu4cJjnDDmFnFtc
YY/XwwwYrhBnYbcJ5dWIIB6JqAJa62An3iBr2/FT9ZAxd5HfjnpeREQKbIcZLai8TsYexkLrtct/
dJUH8xtqNAmJlbckuoHz1PhHqJTnX+JcZdmxiXXxQqrsmdgRNkDotY7Tt4SP9siPABzK8eJz4GH0
HeTgeGT4YLLVjvpfCdYm43zfB2ZqnLGGxGQ4cZSkEqw2VuRmA0PepI//UTYruMKiwVnR6ba1ve0T
CgBfmn7kS4vAB7nlgtWgh99KN/YSGgXtgmdXmHDJL78nDuIdWXByXIYTFkdigLLLPXXlhYk+n0xl
9Df0tZ0eWthFHuTZ7+Lx5Gr+YfaY82knGwYvoWrCqciVP5X/RcJkPBcTqmsQ17pJB7fHGtmramYO
lrSDdqTsUQiY+f0DJaoB6mGOg2GciwQk9dWADt6OkD5cdayRcKRA9i64FvQ4wybfdIedPIN/5rLJ
vrvg7w2mYnm/in33TaAuZ/ImXFV8sqJM9Ss4pOkrdM/ZUZUl86ut2GO0WVScMbVmB+PFxTGFDsxq
G5fbmI69USwDCt3ck/bJy2DJiWuoWuZjm0nj0FcYk56AqGC8/dp/GF3SytIW5XsxDnw04T5qd/nM
700VB6bWA8/XJK8FDytL+VeSmW+msrAeIVEvcq+H8JNd8/rVbfQK5OcKqxlfccy0+qhc2tPVcP8c
IFd81bJtlJlkefEr5HwkqcZuNSW7s4dePy9ZwVGxkGnZeDRc3Kpideb6g+aPeeQXtBKqbSj2MCFD
TzDx5k6b+IfBL8mXJW+woUb4KJAEX9paTDDwCZUe6Ia78E9Bko0sodsFh5KzW2oCeUH3onhBO1vT
s6pwue5Sbn5x/8i4OwHDFhhUMguvxKcMTyK25iCdLl5Cg4sMi5KDJ0xRqDeg2XxQlHZiYx3NIKl0
MN93dk1uZytE6VummNK70c+l0GE3TFKMVh8CO+3XvTG2cNSmcdyhHAj47oKi2G8fPBiY6nIuT6IV
M2lWBTFjSXyIwNmFYPyn7RJ4pKOPphR2qlB65TdLkOQL7zEuEcWE766EcZ3OxNYBtdb/yPngXeCQ
AxKZ8BUxd0tUwJEmm0DRClgMLD3ljn/xHCrAqQyEyJFAeIcDD3ckQzhSTumBU7WtFQTSyhG+Q1lt
u+EcV+N4u01LJMdj4osDInxOBlRZeQXzYxl4y6a5Ou8aMZZ1z13WhOVzivfAl9Rzeaunh3iMEcDO
G0xM3DprhEzRica2j2mv7kEtrEj53yYmMo/EnfzTOOGwLdTMQ3sGcR4GQiJ2tphaRu6KBbHd/1nP
vL1m4SJyCOKvaPsaag4uE5qpIurvWES37DFnMuZGkmSoLzKWG+rtvhDRJjiTzL11/caXmfa/hV2v
BH/nzbB6YNKbDVwi4Ah/1t595/xf0lE6heBC9ChKD2cbJLMnJd+E8MD1LG+bMQTkAK/haaVsICi+
6vkJkPYXWmyrwtX15BULOMkoMLe4Gf8zm6l4EgMmZn80bZtDbmfvbqR6/+Jn0CKbJynvCDHNzmAU
mVIlUCwfW48CnyHPXAAwsfvgTeilmncj3iScwQTboq+P1g/EsVJimrelqBM6aQGN+bSw40mLU+Cm
FHrbJeRius8GRp+MxuWRX3RxLTIrFZPsFKgCT1l+vnhJB/GjJYqBkCIp1zfLWrei76vvC8ps21rf
74+rxPlUNygo4/w1HtMIfByga8UK7eQHyRB3r7YbEa1gNQWF0c/204LJPfV5s4jorX9v2oRnuDma
LiTMNYDtETbdut54fA629Nqp3geL1wG1W3y9utfW9dcLx6wu9CgjiwTbXN30IZBlseNQ1LdC2bYT
S/I7tBSMtSEnG/lOc4r0Gmf7r60AVhyf+9+FdgDL/oG8xR2aU4QBGBIL6vvc3JCBFj3RnOq0ITef
KThgejUO4RKK67FD/0l9FjwRGd4Y63GzcmiFpke50nLSqzLTESVapJOAeSklza4k9s7g4MeryNKq
75+wBY4wkmVUMFPGxb+O5WKJanET7PChoLYjBwXwJsD/HFQE+DabLx5HToaQb9+bj5YUsO3NLs7d
Tjh9zRSdz1WcDgOr6x7mj5H7mNvHu4djWOm2ZzDXJI2vL3gI0Bwb1YfoVWNqOoLMujtXMJHRAHZQ
9pcr1wnF0z2sTnqyTnjV9YR+SsB3Lps1QbKAmxntOBN+RUgboNLu+DPm/f9QHhKk0yAyXysFhBnW
hQ+Jg1nT9l2wbqTTTh32f/icTV8mlPDYNioH81p437NDcavdmO8pJeXxmOj+a7T5/2ME6CbaYmvD
2+qXFg5/1SIiziGPwYjtODmJvgwH9UjKc9Nk0BCqRD8ZW/0vsU4UjkXsw0xV8tvz7CTdfItC/UnO
yvQD3u0U8FquCO0sLYXL5YbGtF+cT75WLXndu6spvob6L4LEvC/VhJ5mgW05/YCJpbFyaR1vIzUK
rzhe7BUhlxrH7xYTH+VrqbwJ6Vkb4c/oas1wIi4U4NunWt5YQHqqWlXH596k0+kP0kStv8ICuBCq
KpOJPP2sSyqmc8VZjDe7KpkpoK9F182fQpBZc907ByUESzGvFuoRnub7FpbQRKk8PXQREK109NVv
XfaIkH+/22BY/KE9jzVgdXxKC74VlBOUsPkjXrixzIJIysYX+DMHK2iaa38s3+tIVEahDC8llE3P
DjHPC3wfDKPIcqXa1h7+P6aM1C3pXDWUHS9rEBrG7W9r37jzPKqBqrwtEYWQypdCsVe7DFrfRL8t
lkFJoYJ04nQuleDJ5qeEjbpm59I18CRxZkxvpLWPErkXAOv1pjxZAHWRpkXdRPmc79Y033adK9k4
GRiZ0ssdzuIlrhPSTW7a1S/Xr9Gn5OVGQntj4/GXFUDQDwVPmdASRHeEi4tyNghIdHP5rqtbDImD
+qETAd/+mGHSW6YMkYo0Ihq8PLh8mVBGJiFjip88Ruor+6VfWr5/+hiOYRme6UVHQyqVyofyODND
HuZMmc2/KANC91YKq8QUA8jskBT4e/f9Py0l2QAhaq39jgag1pg3zURMXnAEpEYXCWGKtvRKDEpJ
EbFLFVM1kUKYPs0SBybvt/jYm6/sdbDamXY0pFNb+/xmgpaBYqjLVHNtqqJZzJtWhQps/wtXv2B6
+5qRCd748Q0Sbhcq/F4l1DqVY6/0j2VlTVK61wYKoLtzZELXdEvhTV5Y/M9HE661Rvgf6tKqgWBT
h5XDZqT9uXtcx+GFQV/4VQO7tx2OG+iD4KeX39gqPgu7cawqTi2VlxH+JIdNOgQS49WXANL7iS/5
Oij05JeNeSjELOsthV9SpwV8nsGFsSfU2qzKX9wZuNMUE/uLgd28nrYxXV9bplCy5qWXYZtXqlS+
HOPEAYsy05BmUBE2HkHXE1Zd+b84+HebCjhR9f+J6VdIxd1Z6A3O9hfrzmqxVPp8EGhV4Js907Lq
8O4vp3mOV9lJKfbgZLxbaTSIbVv/a0onYEAzhZYi6CFxKZkyIxW0F89o2OvNLmWtvlZXycT/81ZS
BrdLzykSJCUm7GFfrY6+SBNZ87bkvB/ehc7lWHXMKz9o9GMSkgZk9ZpfTKMHTZECTTAdNOIP/6iI
HVRP71INHzPhophk6ecz0t6DgouOSOn7xJrdpyWDJ4Kt6JorALlXVLL1SjaMSNS1oGhYiWC3RI7I
uL1kSVJEKiKqEkOVhkZX/TAeEADXSkzMOcQ8ST2z+aBagAs0Pm//J2uvAsfcE5r1LcBa0OoGO31J
T4Qnv50R/Ct0rT6kWeduSl+qG7kioavMznCEHql3e+zgWGaO7rk7NYcP5G3RngkdhhITZ4OYWtWv
qAFyNYAEK8ORq5DWzVwuWxvZa6HvtqSMXwjy0XtsfVhdzGKyqggvbZWwhJ22mBQc191K+nGgwQ8Z
4eIvyalnyJvo2S52oj1KGwLxsj6zbFW0JlV3GYDqvyt/Rd9lgeZYGRs/DrHYXnnhn6bS63OdifLQ
OrS/IRSH5prL0kK7wpd/bODMhl7Wz2SlbcLEpve15iO2ZO9dLgUP2EtFfw0hS2KzCBlro+58u2ry
BNymuQLuCY3riFYtPQgXwjotuErL1gWumHPjbhg8skH3/QRcHYMV4ZHeaI/qa5MFxTjEQWf1/lmp
2dVdBZdLwMd0XJqhaXTPxaiVcVGwLo+w6mTUY49dtKt7RU/kaajffaYBumkHONnpV5ceizj4Fylg
PTpnIcdK+0ZSgZgUfaFJu+FlUt31JFpqUg28gwKKPvc+Rt9M9HBG75EAPRJAeJov6IQ047Oi/6BQ
teWYVp+PqfHd/iS1RzUpj6K/xvoJbIbNN0cHk1NcfUuumCGWS+DirDjf6XIc9zNdB/PsHx4TjCy+
zOPGxLsltdU9jL488Q3RocWoMg81FYn1vD5wnB5NVdovYdtc8UblImY9djlgT3Zy5PtSwwJzgJ8b
gMsaX7gtxdvxPfbCilF/UJnAUVbW2/dc+u13XBhyaeEor2VVQ0WTrZEIh7kCEXT7Pd88UjNvwpKU
SQIOq+6dMsW8uKQM3Y3FLMBT+TtJHsC0U4nFkVj41CtbgZzt1Dqx/jXnSuQxNmzz4jfEKtbvUEzB
hkyAeDp2WCdHTeovoc8Fa6lVuxs6mK0j1AX58vPM4tJu0WzER0i37g2iVqHIlHefhfTcGvgeP4I6
PovCg6tLIHsWN/L9QB1tHrTMMgi0+O1gokgUEMkzOIFRMeUnunLi84I7E5sO+QLfCQKtdnGFqnYQ
MOWEZZQz16nBUvfQjv1eV3YuoPqArJDAXdXdihFs+4DNk7/GhgtE2U/b1jxJtJJQDOdff/f2jBBK
ni5TOrQ725FuCcqYseoyGvkJ59rFFhjIEfkyysFowF0zn1tuMicyoMb9qux/60gmLhbXBrvVzMtI
wWstRBvRdaV5VVOSYZNm5z6ghcav9SjFXH9UenuTYWc95E0480f1C6Wonyr7e3Cj6/yWucoDxxWh
NFk7+OsXWyCeA8dpqhS9xyG3qiEsDm5+uEZU+kgn5fSzWL1vaVR05KqvhdnsnFV4e8mrIN0U7od8
jUd1h7d3F1v0JKnknGXtApsyROX7dLdVJ341OUgdvC+5r5b3UpoL/GVVHBIVekxIjnWpnD8CG6z5
CUAOQEXZ7k/+om4zvyO866nPUb7EM25WuiztcMOlNLcTZHCsBDAEc3J8jkOS4yAYHRzyQYPu4uaJ
RZ5YAeZ1ocNv4Jgv3Rby2Pcz+Z+cTG9A7HzAA8vgchKANXc490orWfRtfalBxcN6nbBfIlBOEcin
HBYiUmn6sKBXV8zja6VFq3iD/ZRPXzPWVMu3m+51yPHPA0ftNyrF7dQFC+6knESIBudI9+W6Nwm3
4xQLwNOz7CuDNnFRfSBQcX2k3MPpifHEWcGA4GgVpV1vzPNmzZDnQ+utBYeWTimw4bqslLvQMGFM
Up2f5LhCjPkS1i/FLvSPpFKll+zOEsVok/jqPrawkJxtpnLRE7AO9jVOzWYYBWJnNqtT4tuJwKO5
UzlwXY2U4lbZdVIuvg9x0Fdz20CzUR8RpJnCkMB2OE0oQgBdtd4kcoOLVBMHgCYq+zIIR+ImP1wg
3tMjpKJnaNJfSOcAReNj+rx7hh+xJHlFXLHlhOVIQCICiejZH6ODW61IzjtPIsviXGwlzYsXEaRu
KFkgfRf+qdZm+XS3Hah/sK1DE4s/XZWYKC1vx9fSJwnQkUIbx51nGEKZLRxs75I2OnyLi9UYZWE7
0BkZEYy3c+JCQRTRGBz6rtKSV6GCtCu/tHZst5Qju5KE/34OqfA/0i29DmnvHU6pVcCdPiWvZUlW
hI2QoGbSJuRGhLvOlmQ5XgRvxCIRaEnARQLxavX3++SL5pdoq8CCRUR7kxEWJBBas7I/C16uqcDs
8TLiNpVUyn1wu8nkoBCtAymhEg9N9v/0XUBALSgYLo3CO9U1fA+EOLb/rAY0AHlZ4u3s04rFLBgl
LnIxuCbMWtJCRw9/n8p+vXsR1QFq4/Ztkvu02XuAcJLFgqFMS+ru/uvuv/Frax+Q8mIV8YOBqE6p
AlFkTUWayUMrpGS2vy2I47jBtzqFex3ao5JAi2SSyEShfZ3+flGjpvgCfTVlc3qBxmM4PJFi2csk
PaWv6amsq/lKQljqqsqw6jn3kbwyV+o3CHLjNw/XQ/PTLSwMOX6M5yxw/MYkfXvkfERH8Dk10tX2
i6v5wt461zSeUj79W/15WaGdVI4EhIHGwG52hjTh9LYRTRuJWP7cyzdh/AoObnQBfNeK+HgF99Qd
HxEDXFK4Cm3FjaVGUAn0ItqlrYgkA8bKxe0aUUhz6uIMghF+ARQVfXsvZNqjumjzSJ+i/LCYVJnX
as0A73PJVM6MnjDDxm19bYSGddzBLvm/0ITWAiGeUlTn+rIDNi5MbIG1j1Tg20KSCuGKoKKRR3gC
aeQ6RvxJ5+/PYDx+fV1MGtT0hOv/PkQDEwhH5uGWn77gtS6JlcTb9C9KNQgnvShPpkDyPCaYN4fH
m8olr5mxvfJgTRCqIJ6S/ESUfKaVCe7hBPkQp9FpySMwWb12zoYBKUIGOPs0/Et1u+Hk1wSq/1d4
k9xO+YG7A2niGLoUilBAiZ6Ge55p2f/KIU1fpu7bt4tqnYnoSi17qpCsWCL13KtCSqQroKG0XRWF
OVDYsnqtRcNh1eMlOKnsCwmgxYfOMr6wzGKj64n91DlEL2g2jCyNf43bmY3FGk1oeGGMqwhPpvdW
KXCKiEPddnS5KiDHeCZPjUwJkShat/EAQ7rvXlAfUjcQ16c1EvchdYd1jZJnBWA82yHcP84Cp2TG
+OtHatkYhIw4rJRGIj6YO8csd02WhMxtyza1mk8pdk0hyJLFeMFhbw34bV8jEqCznbH6cI5OvS6M
iueYazshvxDkMvoNlaN+qGd10T6rqPy0juRTAxSGFzQgxTgJhWcMGuIf8cWhEO596wHxf8GisIa/
9oh8qHNDX/9NxbOJbG/kTMkbyf+FNVGe6ZiHkPDgm1QqjbdBTIO5pOmcE4mW6Q+s+gDYI2+iuDqY
YsFpT/895q4PxJYc2bJ0RgFVfI9IB9HzDIBeRuDgDXrbQ8FSs2impyMQhaVm81xtwkMa/mjFRfse
fBocNAZDs57WWWTrnHv/j8Gmhjc+/nLFohEVi8Kmw0+bNzx2033GsMYMi7wglrXqYnjr2QVW/pWk
oD2J3p0Iuy9N05DlrmJQU6c3NGLqQPHSN/4lK3Z0Q20BibPNQAvqrHNfFTvfXPXeWKs7OcLnMqcc
LMB/LTEIZabFDb0eWR3etJiq3f8UmWH9wdVdzqZS0qkmt9ZtIgbvOTsZMcWtnS6B/GhGo3knnvBb
TVuLXEH1+YasU9Ar74ci3biwpUmswLPIRZsU9lW0AF9dZaxtXXZFtpgxJXxZ+d6w7RWG4ZHHmwlP
nF1/vPnCQp5qfQ+XCbu4MbQA1tKB7mJo+zH4vwt+4YqRTQGBy5X5iZU1UISRL99yisMHnbBhTtuQ
gHdJagN+L7r8fHfmT5RnYhG4wICrbYM3+RzTI3Rllko2c0A0NiYc7OpFqqpJbuDkpd1A+55WuwL6
pDKEElag66o1oCNOoV+EsrQcSfY0Yje+kWTIh5WWnaYvW/zZRdeBjRZe8eH2C3mjS+3zV5ivqvD8
f5W7zFUTaKZ6vIrd0bGshV0e0YBi08xDACdwiH5zIC95v5BuLgQhfr/ZXlWXScit6IY/h6UMmtr4
DkxkG0xQEZGK0WrfH5Cs1HaopAoZP1TG2KEiZgX9+wthkaYHIL7ULzFZmq8hyzAc+leb5YfSdhqu
GPNGbd7jtkqf0+Y8/2IJGuM5dVROxL6KJKP1ZzZYA94maL8wOX9Iduxzl7zexIoOiRwe9QmLUt/P
jzEKvyjrevYlQ9BUd5EIYuXUjnDnd6JMFTEBqbnGPjD8+PY4lq4i+WpkMxfwDKvPid7f3N4fv83R
sKPdaIePbRWWnHLc//2xCQ1HtalkRv4NdFGfhEM1jpMnUYmBhX9a4FOEeVQgGtkzI1w9X5KF+MdL
cbmRk9NRE3gi9JTW7KK4sv2lm2cmAC/MvGdpLTMYEpEPH3Bt+AN9IOF8QZrQuaGEIXzeTRHZhOn5
VmeMv2b72qUmtlhwwUwBAPQGWnAUekqm3rMKbzPUxMDAzjcUDBV7xQ5AvMXsgviJSbvDE+oCjsCl
xkDxWWzONFxek6jTzlisYutWWwrvRkVvl/jP871l7vJSwv7/0BoxGW3niRRIlGU1mH1SHe1Ccerz
TJNr2MmHJ4B19Ig854SLnEzr+R5dqR2spkUn9pNJ0j8Xsv0vdtx5IvAU5qnkzWUolpnjd5CiBEWO
cRrproW7sQuiXn5peIMjFby9VvAp7uq5dvxTGFpdTTg8IR+sEcNxp+J77FejLxWvnk2JNPgTA83e
H9AT+PhMl1gNdVKEkMeu5eiRclb+dZiRzVN3FiTpFs8fn8NvLuW97sGaIKHgoPwNgU4hMJ/1Mugt
Up76hLPJTVk+r0/Ht2Sj2g4XjtfqPR1WIytGks2yeksrofQSZ2hxoqg3kQpk6YCDhkx70CBHDrSs
qKQ0K67UC3fYY+A925rN7K/kRHHc7XIfVGQq0oxyzTut7ik7JabQvtnZDGSEct+Wme/eOIzPh9zT
mqMf/yfspuNVQrqZrTJAsScvSFG1KiagtK2Gs0pbsyGRl49iWFJRjtofMAVTqFVmqEwOJI0yJkjc
dSxRvS/WYWMelkNaBRx6+KqtFnAmLDBJsd6B7JGdODM/PA6PgGDZhxcJ8gAqAQof0KW5ygpwfhUS
RGSJirmqN4uFkfXrDwE3HAJ1dBoOR0FFS8baZmAlSGZeq9fI9yZ9csx/6OgZgUXvKMd2XtFfUMmD
8s6ogv37463RBrXqwHFISKw9RNcxiEM/GWlWT+4sQAtxui2QKWaqeYDyJm1cFEpxNj0G/5bRidya
U1DVkzJ7xieizeXFArgsc/gOvWbMjlNkcvUQQ+qsz8WLB6lCvr1XdLUo75KH2Rc3GHbPnashWdSV
9VZqjDtvExFgbY6GMODHIL84OK/qsd6245V+3mSRnwxEgUmb4ruV+XRdNSIitKxBdyNLfYa3Hr+X
DtOc0ilz69GA9GvRCaWfYO/IWEY6kDrqUayFzxzvTZT1qHcAgd3SmbfpfmwD/Q9womuFLBhvHb3o
JaFWp3aYpDGMZAlRlh0LMYpbLTTs4Dxy9jGVwfzfSIy/uuOl/AA1EZdHFR5duwmHa9xJqWtnt6ru
R9af2NzRftoIYLku/NAZaLPC5ak8JWrp30zQgK1t7oW6t/pyI1QiXqhJX+2agoSm9wYhALt+sy+B
EPnemPAYgZimUMACcrsZ+1GfdSV7jGc9suTLefCnIWnhU78YztWh5bwXHk9Af7ht7IRV6ju1LOWb
TyDdfFT8NZ4DJryfC1FPzRW7gWxeVaGl+/OkzBerJFzewnEYbBHfRnxJebS0GpT+9crrXzrRMAqL
930ePJKl8+e0rNL90D8DhCdMuC4/oskBZYzF18Pgs+wYMdqKUspnDZuJ0FpARDzXeiwEmqodBAEY
qo2JNs62za5h2qSqIEpdZXrDX9m7BIw7tiRV2jmomD5p3mdjbUtacsrQEw5rstHq6lUmP2jMEJif
qHL8guFJiTPt6fVMSilHWrD3bG2qJNV2hPwvGnEoidPp5EPtH1Lwpj3AvZSU21/BCNhXBcEM27bk
Tomy1sjRp7TIqfTt/VeDTfZfwc3NIcHugWJ9faBmhWnPuh0WLuei6g8xAvW54E+Ss8LtCh8Z0xWe
XSJ2CXMAZArKkNSOUXEEoBnANnjcYDF8i7Sh020YAIBtI1pue/F7t3YncP4ClwjadlsNBXNdDX4l
oNdWIFjVIYrGW5YOmu54gHeRttw0ZwfJH/zomJnXjmU263VP6nw+RlJSCCj70YzCjHSxSNDrhrZT
0FtICHECxJWTctaBELW7svkSanY03ciM1Ax58D5ehkaLpGdVxyDSWqXMl9nS6zu5Y1GS8Csl7Pw9
kJHhu9f4PgFzXKMcxOtFVN0Jnlf7maHaqq6DYC089TvBbIa0YCf1NJfhmRoINxEAqwyOL90CMHX3
wpd6KvO9ZwFrQkF/fPOG4BrBEOzEhdOAGMADHu7hSbEsQy/Ur8hmSlxZioUfNco/aOpKWFsy2RsP
Kr4/BgI9C/xAh6hpGhhUXTHZY/UDNhib4ehpf+zshADGAeq4OaXSfk++NQ4eco7rANlE1eAmRmW0
3lMUmlB6Y4Tsf/WzuGsuB7G+X287uAMq4viim0bQWn4ljIs1VvahVv/r8IMz1QwPHZGCgov6EuG9
Sr5TBHME21VsW6FRRcB/ViYRnj2GxI+m/SrubU2nfOqEh0cbW4NNvGN5B2J3DYaEUEhJqeK889WN
jjEt6IhYlbSa7zapjghCS+XswRFx9T3hKygtzSAZ1IOjiaWWaI1uQ8+K8ArW3s9qoI/qEIcg9K6g
0HBU5zbWs5srZ/j98yTLCk5o3aGpDS3AN/SLE+Gvp5TiWubV6jMwAW84At/Jup0U+ENS2tzeCRBk
ShViq17mj/2udS3dtf5YGEhKmskCGqsxG0CSGMMgyAM07K4m9PxXPRthwnEA0d92Yejqriw593Zm
nQtffy4uVUbMvdZK1grk9BhLHJwbgzveGX3wF3KH1b77QvsAfHb7oUMWcVxzbZ7gQbJiJdfEU2yb
noHBnVXlGnA2znisLOyDt1/PsPD+Uw1fJGUrbjK3bQspjoJ6T0/TNN2SB81boSM/pShwC4JfVDpr
w19mK4osYFRBTdJt0BtIWpJPl0g5rPc+H6+1dDXGvXlwcQCti68pD56dNLJd3xHLp1XbKV5w1kez
yY/PQIvzPG/o1I41yaETHLGfQz9nW1OAj+Et6WPZ9I1TgrSdmclg4gKw6epr7a6vsFkplnh5zt5t
ytZKxzOe5YUJVHtjxUR/l2DMSY7i7hjbrY/teEZM9ubaWED36+Th58BngwKtn+OA0/vqKZjQjUu6
bZYf435UQ6NEqOffzidkFU9SgkRpn6f3FNdMvOMaFbcFsOwM/G8NiAvwyAyWgHeP23AbwmlXkgC6
DAp7WehijAzUlQVnBrFX7V0VtCw/4q9gGpHsbvhhnAuMizE6JMe6p3OVpUPNqIap++ZoMBSRZvB9
hYUbdT3mZ+BtXxyZpQKSmnBYgcL+uYsVGP+J612+ZLfYrMzUlj7rF7OGSlQu6PHt6LV4iUtS9Kd9
Ol3o9cWYGm6opQQIw+85bKWXmbb5k8pJ39d8j5svHksghK6l0DzA7wMl+SZY8Y/aAk5pLVsqsHHt
fVAiObGvvUZQ0go2W1ncA2hkiy2QqytdG3vnoUirVU6+FckXVxikzorfP2OWOioMw1jON1FAQKFY
CDtxnvRdZ/DDAVvnEi76MAqtItuxiNgk3/G+y6LhVEtOSP5Jkrm2z8EZhGaH5hY8wujwIxCYmPlX
cjbTFlMfN7rqyZv9y3nFrb1KRNoclBtGEP9a+zhOQGvgc1Ce29VJObyszQf+fGjHhwg6LlnrTlKe
C1XmMzbuUGitTq64i7d+i/5HQzakSVNFgTY4HPLAxjTaZZPSRkcopHEd6QbQDiR/bCSImaXg6uJc
Ed15ERaKTAdaR0bgUvqfl9nWuc2a6ynv8VYDIalpFEj0fv+/iJO9BDCp9KgNX3OcK82ZU0LypPgr
vg6GQnkCMupL95h/LH4blKwkSguBpo78AyYdP0GdU6Xmu8i2xoB+fd8tP3wpp1IIFOpO/8Rw3nka
TtuheNQimSpZSypSJDcnw6y+pU7rKzrY765FgAHaDgoFeek4M2/gEw6Zmz1wVOGe+M6I5vHr1sv8
onbAyoOwKKRcgWENFbdxR2HzebW80urJ4SIzRPUU8Qtkt8ksBzEzXVdoAnqFFowziFJ2E7uw/NKr
LxP/Wughyrb+kkUTd0nTZeeRKDOoMFiDhlovWFy9IstN+N9M0b2N1lGgpz3n0VrprtyyJFd7cMiZ
zWoKLQBJUgvq8jXFDMbGBJxDBQmVnsYrcddkQ2TsJPHFJwNAI91pK6oGpG82C03uBjCl6XLgpoAs
FUqS7kD270E9VMrWEDYOOaKonpS8QuD60Rv1rypa/ViFfRm4eqBI2UcHTCdHf+kkK4vVBnLoBMlQ
i0oH4xn8RZzYXTjPF3Li/rZ//Ys/RNs7O3ESF9Eu/GV4hWWvXs/j7hvJQJt7ZPvcICqBQtF1jh58
reEb4EX2m0zIB3/CIV5USp9OTAPXJq6YhKWkvAHXfv3dY5yBSkcc9VTxvpou1t16wAR13R7UFwWD
h28HA++S9VF9Lf61n9LLL4vjz784KrOhfPC4ht4ziGrXFINgy16QUHsQpfIXpuRj0Fyfp55BtJE2
dxI6D9DxhhVCu99qBgFhD8e40gECbDBy89ea6OcVt43ppTKAegwkRwi+LmFkFJ/h7F4cQPvZMEzX
Nx/YWMf3xJOIb+bMTb/MQ5Rc6D+xNQ7bXr5DjY2aneYAXuG50P+RH3ZgRSTPXSQy5lPse+pN2xLP
u9DvUtDURb4lXFVzLCn9QQ2MqV0Dnu/o5lVGXIEvVibtDngCZUq+5G+sUq7YoLf8Xb+SXExjfvkf
eI1b1ftnwOePz+6KJEtwr0HfmqUutdTaExnDG9T1ofigIDlu1CrEXcJVsP/Q9X9IJYsCPyUlm9cq
UUXvookd7hx1MIiEAuXni0q68NQishx/fBlEb+vMkECTnKiiu8HlClJKFe1o1fTG/zmZ7ulIDrMW
byEAk0Vpt6ne1f+i+bepQxkrD6Wj1tI/iFTHis7Sp4pwlItPW2PdFEjh1Vp3kuoWyWXoQerV2dST
ELGrDzx7nD+x/J+cOt3OC2garrNnYk65A1lZKxNqtOud2iphN5K+PUbFwItblDeKGEPM8oVk/xe+
hl3LJrbfUr8oO5ILeVce1qkDbboMfs2DJlN5vTV/fT666sh+/KwH30qXDuyRqg3ReWYqtJLbdcFY
zuZMvpXxSzgANIq0iGuXVyFVEJsYwjMh3ReHPjU2NaJnLY1+XobzPke79zxSR9gAdc4c/Gdqf3l8
4rWiUgbkPzJlngtW4ghTkAcicREyltotZ2WUjwNo8iHTYhYIx9Rqzku1TOyVj0tHHm+W7VXMC3Ku
nAiaxV5WijOMXOeLP9vrjgpcOMc8CFSyJ1E40VXjS/fgOhF53CtzzbZJKkSHDSvJ4OOuhIZSGRG2
k4CG2h4EXrEXyZs6zFfNUfrLqD38PdhpR2PAjat8ozyNFf5RPTUH0VH1ahAi2cfomK2BP1pl/EWw
04WXnkznNDx9jcUjYaBek5pBRbo0JktEA2BDuzojTTCGP270yDwHdUUcp1zkgBfBE1SVqi+yzplj
hkkra5AA++JzX/LplLafUvygBPIx5b/hGZ7rHtyZSSQ/GrxlPvV9LSExHgXIF65EPhptLlyKSkGo
LJyE0EDqbFgK9BXyWDgpDDHpOBgiTULgjjlMeCg6n/caVgSpNFP+Bpz+VmaIVN/wPYM7MbSxkYPw
YDIDAW1w4HQHWqYlQaQIi7AuVyzkZbK1Py0CAYojuozEx/erWvDsA1m/RYby7xkvQl41E+18fBSQ
tPCi0fh4t5W0Q1xhXe54OmpUUGcuztHnaPcv64YV1qZimMt7Zr/viNSEWuRv7W1NEp32r7EcIvOE
4PBeLIgKtlhXo2Pr7l8VhtBkJz5lymn4C1sxCkJjnaVqGNskX7blt6jLxlPYAIuLhn82ktvFZpQY
4jDiBPlUvJBd/PvSu6ibSh+frQXYl+2IqBz4g9RlBqZc4tIABQ+8VsoA52562MJsuhKfDRcuZ8xD
8IK6wRuTUDeMIvOJd1Gpbahdbnv/5hBBA/j/ldp9cjYjSrFa6zRW0GolJM2dod9K2cUM6NiAShY1
RAqBBgKKZOaGqkY3m9gbYBeTw8QPcaTMxQM7dhJjWfq30DBAOlVN9nbii1aTw0FjiBr22uSjVabt
oXuoHA6lNyIasmTMxPM+Qj5KNipcA4DtyAQSTKCJS2QleWXYcuNpDgFe7Fj8CHwC0epp1XsjgUtM
IY4eUxa2AYymUm8ZuYMuY4W7275Vu7yUhR7eNwBGF+WCscNvZ5EUI6r6RinbQBPMLtY/DCcDXADS
vfNtBJr4sopw4dZARKuNodqCY7bueaSD5YDiUH/lEt88eTv5V7cSaRBDQBEqTbdWzjairIisOfbv
cu8JT9NfIuSzhMvwM6PSX9J8mqSOKamhm1Hfo9ixtsflFZn7Wl7QkB3VcF2xjD+pN8wE1OL8JO6H
lGB4BG/5YyniIsVXiazjxfnXSYyOX2ABDjmFNAJYO7dUURSry/S4H/9ArhL1z8q3QcFeGovOhi5Q
VwjinLdpO3tXuZDxr0MX0b+w2dTk7KBLLYuwgcNFPV3lJZHCkdGibof/Wbbw48pS0+Gh66rVDyXG
eR6/+OdpwtIQJajNlxvJTi53z5kRrGKztNwKYvLbArSty7pHah2mtFD82En67ah7Fa6YNC28zSEL
lMZMaMuy0Cc4u3mJCLsCOKSz9S9mBC+wslmkWgKWOSz2zOq7GTbxWoqKx1M0tpNxBY/07Jw+KBi0
gqxYlVYAdXD1+zqazj5pXOD/LmSYNsiYozB8n6054iusH19APGlUAe6A9h36Vo7mJozgV4Cmklq6
is4DYwMFG/kX2AzyLHaPBAqpK+CAqIxN9hVjvf4zrBBXKIh7LQ4SZNNKzxGUv+7m3xgzU/KVMvg+
ahYozVOjgBYkgL5Cl7G7TZnOSFOtN/9YgLUbv0Duu4wcORJF2q17IQCo7Yqazig+PKYl+IkFV4xR
c2EZDwGvNmVIhzyROq5NIlUzfrB57evU9+lhg6qDBXdqvFbaAxObzK0SacrHFLoPRFBMEkHKzjj3
JQXwZ3GTJv5QjKnzRCp0oM5TOaH5WeQwBFe1SVH3c9r1DJXPC9PVv8IXXKWCl1e1KCO7lf3hYrdP
T/FOQBPfnRHu6ftq8j/F9/c31W2U+Rup8FKkcnIHJGSDWS198rUHfM6RdssDNK9rzWPkqg2mEB0W
5I+domWuBTgbCPhLlqZX+Kymbu4WDfS/UlPIqpO8XgYH/n4FnpkWDvGThdyGvYWFEiqAPZF0Yvym
Ks0Lp6h2Qh11KYbvS49rFGVroRL33If31akWTYSpuR4qV1wtrI/vAabBIDu5/uP16PPwt24JZFo1
DDk+K35bj5IXE9m5SOpnYe7cR/9WcQdcfRtz+kXxKpFAmC3PdeRAUDTnKebq/MEBbHe35F7Uxb8A
pjToUpUIBNRYwfpps3LJb3073cuB4lvTw0N0Owzcuui5U2R+axE/EiFgjkv838S5yp+KU2Wdr0WG
JUQPh0p/nJGJscflJLakJ2ao9ve+K5mRHym/nSuUKduATpwHw5VWuvqHExusinAkjWKQi9K7RZDy
sft6hY5PIsO2tTuJe7pF771uLqXJVtBw1xWdfSQLFWbTztSYZrp5WEDeWWOUPAZCNE/lDgYnBP4D
7P5XGet1YS38ZyjP/EnQTzeNAiMWxSDec8gZ+B52JuZ2nqs7Ty+Jd0VIE01KwKEFaU8rZVozlR9U
L8z0h6evV74wwrf+FTt3ChYbVT4+64MiL257tDvorblZemTNYCAtTBUa47YIb7BWqh0mc/nOUYyQ
1kvsFjxXpp4oRgZIdWEse90T0r82HWNExruxst1U73SsYvvPV7Gu5Wv6F7Sh4FuDmLQDGG2/fZ/d
r93Mxudn12T3qcOjwbW4/4dPQHLo6fuOrIRsTH2wphRKDHZ0zLfZYzSekmWKUZfIiQh3Bs7sU4fq
bn83Um9bfa8otYJg/shnHdCisiy599mxLUCitcQt8B2PWnwcYjnPFjmBi7DFdZPhKTiDssXW2Ux5
lFtJ72q5BKzpDdWMD8RQC/EVtgvWyWSeO+yWD53p0P+Oubd5bWZ+ZQZAiqQHKWfyoTtkEeQ/ImG5
OiVxmrptVi/XaxL7n6deg56hgMlaM8CDrygRkmsH9id1T78u0neXscDmP9VlG12WwQKEeQQ7T/om
x4Jn/SBFkvxKctUesCAjNh8Y3WI5Rw34LRlV6SZBnmaf7e4hKOU34vqFjPtfb9eiEPl0DCh4Yheu
5olMp+J674z2csf4M1tKwg/pDFJiXAGdNyVEBkfqlBPT0ciCWMXmBuADRk55iZsvMhB8a/zmcGi9
1C75BQrK6T2AMri0y+Hp0xkTdVz7PFQd2D+DKo6r1msUj0k5KTRvmMaItSRJmht5R/pofhkqAg4S
JwyGYrGLxdEUIhjsoxmJTT9YXCZeIIA+AyljCdJmTTfFiPs2lTN3fpNc+fsYDRhSum/PiR/gY3Qs
IanPncGPeZtk0R5aBy7GAKLc0VPusyfVoa7XD2LkfxXgve3vGIRzCPFzkk+5LNYmsbJbKaHxKyA3
4FwD8WXsYegLhplWNbpw4G4idaB05hq1W7glRP1ecbxtl7UofFAqFR88LmhfNsyhZXz99UNnRTer
FpzNYyra96kPTdn9Z6DWSpeAYXYqh+/Ji7F+FSdyptHW1SnjBkMx/KkF6hZXMkol/0RRM3hK9T5L
R/TN3FAxL1KF23luHuXxQs2JWeiqrh3viHpsWpLyy6R7yUlCYI3tprFzeMxz1q/Kj8ZmQZywk0aF
G6XU28jDSweYJQDKNlsNw8pg6ZHsBhlp2t8+WQSt5Jsuv8uRYV606dOUMf45yj1N6XXF6sA5SMIQ
ZvjKsZlAE2QEdX7d53S9STRaCdv7pfjoaKuhkyldczvHil0FbSSyFWbrceEPdi6tmLJiu8YjG/Qs
V8y2LakuylBkJyONKmrrL+frvRDbl/JnNh4GgpYrzjJeaDVvyHQXiRDPq8BSY9hAT1g8t9Ae4kan
mMDEGzzgSSUCt996qJAY0l5nEZrqdeNveo1eJIeiC82wpXpphvdV9DGvqS2mqDYMVarg2wHVGVht
AvjKxqyJZWl5K3g2WAXnhB6Py+2elBhFy5zcG4lIxuVzYJwgYRD3fDdTsdKYUVV0u8BnBALWIqZ/
TRBOl3NmyaJrn/pHyxEPdFtDNB2G5a+U4Egeog57pZvClIGT5Y79CdJOB5fMrIlZs3jQ/DlFbzZe
bWa5H4+wUBLlBsQbvrhg14oyiiZ0d7ZPDCw1u41OeUeJGztbWBkVrinfxqM2rRUVi7s/XAUOR71V
QnU0B8HPrFv8RHY1ksXOFm5CPDQw8TgpxRlw5WmlVhQLqjOXdcwHWKdyocIz2DgXxkh/TDkxSRsI
9DFLggvMbQ1KFDDQt/9bqEQFo6OB7q0vjwd7x7HECOM68ohFkaMef0t7ySXNtXxt650pmmYlIEZG
A8BI0N7HMfRW4P8mD3rIVH+B8X1UDFnNQz035LHvuaHm70uzgWtvm9GUpTtQ4n5xWeK58VT3/bZw
JQO1qdOGpnizb9a1c6PsRm75qt6V9A7imT2CCTv00c2+QE2SjXQr6BrVxYi3WL+OQdWVqg+zpbG8
BbGIs4KimxM3ZyPEgLWkArbQPdFe8w+2iMJ3WGM5bRM8xRWb1JGI8mSNBLmmcDHI+fdT//zXWDr9
O+hLgdrM8n3+tbXJkew1l4nfj/iMMSY4sZkn6e27iwSI0ISdMCM5uB8IFxwmReCL7Mms+dznx1KM
gwCxScWMfe/Vv9J0B3DyLsdAjRF6KYU4frjuIa6pB6zqzTiEcl8o0RbI7/jylFYsltgXHR4/pi32
z1x2OGppK/K2qVexTe/vB5nCEHxc3yizx0HpXk8U7uE8QBQmqqwoLK4X54k3jdIo+JTcT5YbH21T
cSxRHhs6gCex3nkhYRiDFqbvAeKYMDBqCB7/Bvh8hgqkVcZQTggyHoy9qhjw6fO0sxc8faL0t7OX
Nease9nOuqsurtYxmgL4Iza/z1kJ2Z1dT7hqk9r3lkfU10eY8V+Pug8R93O0RfNFVrfr/CcgMgSA
CDYa5Xosh2cF2uVIYVK7fnV5qECzhrzkMeMgUp8f0reTXDq/CDTUC2JaYRCvlyVbYWjAZZSfE168
wbHW2/EWa+rQj6SaBY63XEyh7fZK6fyyccABubwlFLHJZs1QWTVBkiJfGXhzbIHAyj1oUWN6+t6p
Mb/NWC83WGZQXfKPjUQ1GuDkFYPA08SSjFSX+PaU5fp658b8bU1HlaXI23poyhTkzsxE5HkZe/ND
W07w3k6uLeMuRt8TbQQc8j7V4Y623O5y0IIfydX9XE8myOQ+K5d5bKMvhw2T0HR+FP1xClJgmC6v
VHM7KiDEOD4CrBOt6DOhuUemdJGHfasDGdQxOPgZuaQU9mR4B9lvA9S1bzXbnYSZXFAY2Gfp88XA
etZdov+q7T5dQp4XVcCtk59ruStj26dXDZ6FhtA+aRl3RPz/gW3rpJ/A2NE2Y5y/kwke6l6BC6/l
2iwTZvJ5N5HjgByPEo83c35SQeSoOR6WHFDy2OsstsWH2c8A9IS1qYH/PDGl1iKT9zom0XbMSaYn
sHQYH7OJ2Ag4ageYRQIreB23i/9PGTuqhV6uaWRM+KJP6cBCwQ4a0xhNEQyh5ZweykCxBTHTkgYT
0Wg3+GUqHipQqvZJd38fvWPiPrER3OyBuftoz9/5FlkVEFyIMsz3AW2HTsD4zkDqG2UyJDTc2d/F
RRrdWP2PJ4VZvJ9hlNJ4ItL5/FsiBhsTotjpetjyEQxix6fdS9WSpEchli1YLZPfA0Onr273zzRS
GhCvJxKG862fwUnA9iH2LG7hFt3yPihEhgIH1lCwpzy7xUlCrGFF1yqxRUFhwjTVdLVDWn60MStA
Q/5BFWfm596MuMVubLvcGQNnIjzzUDaoxalWpfoMzPdSl2BVDQpp6yaT3pcqR1UcrNmIdZCKtXbl
0eCRQjRCI6MPlCBHZFBMK4PwXkVuKt5U2+1OyRwGaWPfSDGz3ARx8E8Sf9ouLaHkHuaQqkiCXO3A
7pj9VRtI6NC8is5aveEAMpArCMYEw+nqKjvaUj1k9G3LR5C14TbszAQV2+la0uRezDZtopjNoUbI
JMRaMqI3dfJjyIohupMZeJUXLCPd6p/PYhxY+DuikxjAQZRJNu423smNhk3gVJdrwzmLSu/XAMBx
OD7SUxeZmCQp8pnsHA39j0EMq+n+QAGGwG7m9sDXw+EihQO/XHEZPpqz55NWGFbckOGPty9ZjK67
VYBuilNJ9+mhRL087/o1TdmOBR07sdJcO4TR7OxdDkouWxBEG5/BTQaV3zKwcssWDbt+kOv6VHSJ
xkfIIkDRonjq6sYJhx1CInRXuZR5NNXXA7cVuPFPGc77YFsMI8PpeflGrpwM81XGiM6ujfbY3MH+
0yow2A2SLHyRwJtk3QNHBqsh7vLFOZY8NA+JGya6jFNDtoVRQlRTLs2YgmZ433sY2Ubjfd5W5RpT
pRS2RaHKpIzs1FsKeKPW9XkRKP38v8nJ3FCCa23sqBeNICuMYtoowsiiuA//GLUHX9HEuXICJqbA
4ohRoWI2/EeZaC+oKhxcOWF0gC+UguAXmaXeacG4bm4VL5JZgHCPT8VvJkoAQ82pUcJXIJpD/LV+
v98HCsEVpO199KvXU1Q+OAD+WexqJ6adfeuiZWoiezP9dEJg1bptVskhiodrZ9sLW8lvdt/0XlP/
wGiVVzPKhYf/HoSuP1xyD7fecyTFQqVwUoALbhhsZruzIFaP5oM4UmdcOlb31FSv+3TImI9EiQAI
f+/xIh5TkRgeOS8Ey5KMAFLFTK7OFPu2LwVcXnFu/hpDkOg/y1b+JmzRnTy6CDfYDV1pXSnbIJ7E
wyR1N8V9zhTVgHAkJGGZ3rtVJ2ku9kcNpkddkVYBcKjmlF60/pxKaRrL78f+DauSMh0maGFAvQH2
861JsrTYr0o+aYrSP7p4rvX7lcfks4uUj1Ci6A76lKxZAsNl+HzQl49cVksrZrIIGlE+3jY091ID
Nxvpc1Nk7ac92FWld2ByDs3yuJjjTuBSfK/KUED4IRdwDFZKmNGr5HOaDjP/VbcWL0e9VwPqa6sN
2ipeDViUYa+Dl60P3urQgsRuaQeVFUd1I9sYiy91zNbEdt3Y4dNzqua+3dtbSWQm3Kx9HYuTyAHi
Rd7OzfZEu19TVb525N+P2cJ3cJJ9ICLkbDeQLYov/apQityRB4daYA9I+mkOz19qmC46zfLdcynB
tdAPsEBOQg7azy1R6ZErkp/XnGyMajoFumeDgCJ5m6cY4JQ//HwI0c2051CFnejLGMTdjIs3KaGy
RrgcEK8MuBhWvJO/jFXO6J7VpQoJh2w8n7gBVudbm2285jKMAhIEcD0eqOhugkSMHCiJXEpIwVi+
52vWVM0rq/OYXNkqz4t8nHxOpqLPHqam4SJ761kKktp8OIaR5c9s1YOvLTKWvoLcSYmQ/wL4UCYO
4DLpWQc+N1Wp60vDE5fbOWEPmdQ9z4K/3RHx15fhLdqQXJJHaF5pPAeLNWJXMFYLvBuKyflD8crs
19P+T3kD/yX2/YgbxrO5b8VvU21a+zwh69msyGg6D+UT0ecO5dLWMQ9NuRczZRD72ZvMjjmd33B0
hfTtXu8dqyFQXXW7/2v3NYW00gfCjjNEa/G0NGkr/UylO8yrWEFjYCqJ2pMF10B3KD2rc+hPDm19
yLD46kxy5n7sTyR8HDK6CCKii0jl3uCrKYfAvqdL2t6c6K2CKNCw3n5JJl9NYjN1uTaGm2HZxSxm
z9UDEVI5uCyuEb67862RK7H7BulXD4yoWjvewfV3byBXQLezpMzL+r6iOdzsNnVzh7WoG7fcQqmT
PMV72qISe52DRR07Rp8zVFX72ViA2r1M00GRlN2oEzrHpQFIXOZJBW1GHd1P4NlRB44zjpgoLrpv
OfYygLDNWh1YtYcubJcmNQGG6TVny/1JepiLrTg2ZFYOuvYKqAEUM3JHcY6embwX/8g/gb+cZDLX
MHUPVj1imgJyIgaLeY1uq6jjv7+k++6oSuqxo96TqkVYq6edtYqFEAMzkKGRjSSYtj2vSV1BS/kH
PTqycx4BKTx+7BszQ8PjE7MOIze/WzZVQ2hBMDCiVhxIhqxsEtVl4IQLzKkjYLC6IF7um3YlQD9C
CmBXO7n1s87AD5nwUHVzQPYW+bEvF4gvagnhI0AMrqgUmLMIp96ptLfS23XrwKnH+6xUBV1xmjcT
rgbX+sm4IUAxbtN5PeNh/aI1l36tY4VbIl0pxa+5jhBocHNlCVu32qPhZxKQfU0HP3fTj/OUHOmP
m03pQIzwYL6Sn1bcDRkevOsAtY2ZeNXJKjZAC2uTr49XW0caG60qcx+SadBUnAggVg+xBYaAAeij
YCh405JBO6Ng/gmsjIxqYgpKJpTGSfcXA03PFzph6MVBYUp+CGMur8vTbQ+zTZMqS9Ip8omi7J+8
FGOHA7dMRO9wv0VTBUMaa18xjCkwkvKTwHAzkwR9XN/iaHXE5SO9eSCqZuCATrkvDjs8puFEzhct
mJgO9gxli7N/+ldSGV5uXeih9OCY6GnvKqrxDWG1CRw18/KK9ZsQX3lPUicEkM4ctgZ3IQFpS0JH
/BHeEvqTWDTHQ/Kw4r3Zt4UEteCxwxsLzd/NQ+OCQ+Tjo6EVYzqq2VLHG/C7jznJtI/LZ4FBu5U+
tY2ICEnCqRB6NoOiL9wOeE2HbInwEyPS+ZtujX+IwzKDFipFBDXXsUXc+TzmgYnguqQybpWR1sDQ
IXAS2AXPik90Ju4GNz4hOKqqHcYT2GtB3+su3MkRSQ6j/GEYGmwEi84+wp18r7Z+dIKc2zVJQRvr
xngOKMpSJTuUM2rYcmk+9cOlV/ne+Gb7UnKktTCmyL6AgmsiQIX6Wy6PSoofMhNT8h57TH2YpVgw
khAVUj4M3qnIIlNjT8ebum6OGgP7xuJRljXEhLPhjNhhbzukC8uQkpao+goMuMnRF3KLs8UBz4UL
5KfO4or19m30aJYbwSZTosc2kSLb7Qh4WbdfxQSfqv91w8ne8L/xnnr+JyGyBbufak2PdQXU2GJ9
xroPD0OBqpVzvonPT0lUbZJuvBCK8qBUkke8siTI2CtlUEmf8iPd6bMR4Sm/9ocOiEWzvyQkvRUX
Nx+ucEjQmqR0ueIu+/GOzI+Pp1RA2jOB4kdekcHbkNmFRpJjStQ0uKLulHmjyf27l0iKFKJJ/gcO
vJiRzctWQHhBtq2QdJAyXhOdN9e0RLcCPdpXzIRAuKoO+kg05l3/rVN77YOAZvcmw4ETb9CEvkvm
HXVEeuZbLu/nUv43MnGBoxBcYpnNG/R2YFhoA/8fBig2ieNGlV4LUuKVBrW7X95Y322HvhqKb8/3
JG7/f360Q/BQOwejtpd/hK/gIr5UfAo130ynM53jgwJ9gtANsv8Effe04NcUz/U35mhhcaj9XV1c
3I0eqvGxgumLQLbA5yuxkGjYqhFshV3YyjPo17AcsfgEKPMGqYirvBv/n/ri1Kd1OIzs6ll3W3XV
WAep3hXtAWc+i6kMSlhTrJo9UmXNwFc7hFiIhfb4KaVo4gO8jwlvDYO9GU4DUvD60fTa8itjL+rM
Qd134B+LQk59T8TumIu2horYbE92AQLWoUHoEVJWO0vYvsSuuezTPemJ7YCyWfysrPYIYe+QOjUt
WTzs4bLl02trK59wAbAVYksldsPQ0u4sVIfDKj6kctZeJA6FmilCXbYkJaQ1krlFYm4KnlVEXlzp
5OkE52HSXlr5sg/yfxA+o34rcRCK3P7V/5P/aFq6By9pjsfjL9wHV6qWxs77m6WrvTZxfedDSUUi
4Fvz8hPOjv0OJXzhI8ogozLCtQxhIRvwuR5fghkfOtP2YEB+vOfyqFbgCTQDLLIoEpsNizbIXi4w
Trnn3t2ZMB6qL1RIFWHM+d4R+CzzOeoOSHa7xWG3suOpEOcJRmtmi6gTIoQJy8nY21eSRcUKDmW9
FJwwS1Fl87f9h8TNmk7eXMSUS0y6iVr+NGQEltxlE1YxzWYFp0LdOy+uXyQm5Zn0Z2Ib0sn5pT7n
DVaQM74Ka1MRUyIkXUdNO2EhDaoxaaSCMrO3OuYhBeENFjDzIVh1QYlseK8Ck43s+SM94edp6Dzm
UJFSJ1O43BhwnLKk+nWvcJOGpRBygW6P30Ht9gEfeGSp1X5ZYBJrMaX1yo8lzOlQn/xGf+aacljx
lKY1vNr3346tz1TYOkHs1ff747FxT7XUvdYaikran0VmbhGsu4GImx0PblWwYAlBMbwAn+jwk42D
GoWkPFNneTS7Q+7tDQl56kMKQku6V/QTrODGPMsQZnyvcNLQKCj82vfcWQdcJpVSSuY/r3Mg2dCn
BHWd3f+3pTUDrBAisFTNdOPDEqd7ElBbkbGA1USrMKpiqi4H0a57CBbyJKqZO1xOhtpPoEkj+nT4
SbZUd6hBO0W29xvRnzc+8lkviLnGsfWBLCSsH0qOlP2RBaGrcGwc48eyiVCChiNu5AXnCZHu78bd
EQFzs2iABKt4QkoWSQLjiNUqJl2LIx9+Xst2vvn+JLEr0XSFipslw9evleDYQcBrz+vBp7/1j+xB
fBGb0ccwW6A+Zal8oKbpUVvoff63CBFcyqutyxwXw40ziYOHAI6maVrq7Mad0zPJQAvIz1we2tA/
i7V3/OLGI9Pcu/Z+BYduW5PtmIrbsTbObjqlifWNqZ4WHbyOg1WAkjvpddUwZIqSozsXSqkzgmus
szdpmPZz+KuHyh1w0aCwuqzyQvycNrLGDsa8zlXxcXOiXS23281nFHzbHCve03szu3k2D1o74TiY
awmhMMiLsdgTYGt18fGrU3BVWqCPg/x2maW4jn6gWkvb/DXKQUBDH20c95hDg8LCsq9LVgHcVtZF
4Girvc3uF9ZBb7vn4gKOZdDpUU1XxPfEpfri5AwBMAMSgwYGnZUE5s/i3tQC5/ndKiS8AdgMRpqX
ETwT6vClXRIHMywMXzwUMU1sIWr2sfPDArguvXb05ruoJmIgrwrZbJ6snTiPUd3LkVwDduO+mGKc
gaNr2zIuF7LQjeXn5Bp9mLt9oKv4GiXwutWptpMXEb09zBISEWTX35zpHZ9mwSWV4WCDVdqML+9t
hCUFiX8QiTSmTgfmA0uu20CS8S484CXml5tNOp9e9mIdvI5V67yb5CzcNQWsUU3f0F8bae7Bbkus
oYUkubC3hKD2RkoALpVN8xEWFIT68kgBxEPqLlf/vvwdUQmY+ZN55M9YynyFP51thrS8+Fa+xVVr
Ap9BSddcr0qbloO2gnemI977UqPAT8vq13Jc/pdAeaIdWHMfbAqzv3R1Y3ldOpOlLeegCgGv81sD
UUFCkiPKYvgklf57lxpevn03xmHrwQfOW6B7+SBixHWYU0WE5dNC+TXjiD7KoAJtzq16hhqwku+U
keZrcDateLQNIdou+LUNj1nGuuzWmnWuGK9sMcHc4OX2gelF7GknpJEwe6sQYN8SjAwkTuvj7hJy
M/LSwCcNzgFtLinOMR9WDaP6b5wzLoTVwU2OybmVJHvTNA6jkvKnJsZ4brQ75OrMMMcU4shDYqjy
g0Bnu2ey0x8g3EP5Ob8OwyF/qKfMMgRAqsUaedhgxq1gsPSmepfUOMiq4zvv+T0AwYXj/xFw3gQr
F0zfepilNik2pfVlqzDc4xnZZeZ0ZvckRW8Inoy4bmqmr1LtRfn4eEIzpsQ+H9tJNx/4FVgd/CzE
8I7SCQYlJ4jF3S/rTviO/n0tO8qePfhS4dcRpTby0474aV2zpmx7Ooqn2XKytig9qQA/ZfU/mlBq
NX/E55rXc9lSBwSzzePjrB93qlT44JqVgDxMzdUcQS1v/2Akn+SPQzbmes02yS5Xnt1Bl+7Xj1vk
oxhGdUHFXfnGybAmmSN7oIgxRBtHtEM+fI4kvVbFFyN+tYfNOk3/b9rYHbRJgLVLBG1CO3HD7Y4d
PP/Id2ZfhFlK4oXT5hliCHvO82bfGaEcFBf6EBTApZ+njzt4CYIK/40b55yIJEggv/H/rh6fOcRX
l2OjO6Qc9NIyI3CJKmX7V/eRPldKEr/XGV8HAXMud4fm4hUdFK4Aos7mzfFcDS+F3uJdHBlOJoGp
3+D2IevKtqkSCoxqqX8jCNjblRqEZ9tioV4cqYyfgzavbhbBSus6i0pVNRPViXN+rVmgVe6l9WMZ
vtCZq3R+A+LaoH2cLqOOeYhDVoRIUkwGtwhWl77V29jeEJFGz6d5CXptsuPU1qaUVK7kC4X3SbNs
utd+6wGy7wNCvWFgIgGhsgmSWS9kz5UjmtXexfyftIowysW30I85KjM1yNlOFuZjnN6hYgUSIdlL
ZtbdUK1P+I5rZR8+MePh8JQ6zylI/al+9WlxZpRHyyO68y4xlUf/k9b7voH/4AxI1vmkZOi9GqYT
pxx9eW3XgiLkQIumSNCXo1Pd1dUPnzPHqx4RXuOCNqMxlMKBg2XCnUYUSJOup4xFH3gPWme7o0zH
Aoat7RP1VmVkYoZ1YtO6gRlKYbNIDIh4EsVqz12J0KW4sOPFiD+V7Sbf8VNnHQJeTyLiRSEiuuPP
lhrZTI90mB5mH/egeiBCklyOA9Pfk5S2gfM0NmuDAQ6HTHs3QzEDTcjcDgfa6uz4ppwuTOEC3ZRp
eKpY/YKgOsRWZJScOpm3wa1UzKUp7CoMPQ1pLTAJsXWamHoR9KuWXgFFIcRJ3i0Y5kC64xYYA5M1
VCw02JofXyuUCrqNBGO1PVgpPOYjBwIe+m/uXDf2XUgloUYYm+e1veLXOrdJ9MUkwH4fCf8U5Zwr
/FKIjBU1DiFGnIqSS7IyxMqjpF8fmsJ7tipcEdxEoeAcjXjaWpPux0uBFUjCuFMg9yi8r58QSrSe
D4nuh9Aa2uwRXSd4yqa5nT+rNi7KotMu4jAcFX0KZmvELfUldolWQKyHC0hBwblMfBpewu6geNoD
M6oNQaKdzjtW7JbPCbtvGk8aU0J69hOPFJa7ybESrGtKP0KBt8+kduYF2QgB+p2dJmpKYWqEyfhJ
3IsLaegKhRVzZiGIkZa4iNUU60JIAFfwJT1XQLKqDkRHmHRERP2Fo5pbVfjEvmFTDXxj8Nk6ZdKJ
lFZ7sC+4hMwHjcjxmW+j6ljm8eyXS0GJ8v1SbMzsWh1ELULeyMJJmyeYBpTAw1+LukLugnxcOfZy
qgUZ+33dQlyMi4gFaq6ggF4Gf+99HvWmeTu47dhIb7/mOf2zCcQW3hiu3YDCQ4W6+CHbC9AR20N3
ouqZut6k/ik5XYJdiHixdf3YRFcV+Gn32m/pkHB2//s56WAPpetqyzvl0A9G58bdMNotHQ9hquUE
h5pnyd8QaIbeZGuqZkGKzg75vrqSpsaruuD75ja42y46dHPMOSliOB6CTYm6CIW6NfqkiNKFSl0W
nOtRy1cVz4kayewc0xd50keR2BT74J/1OYreCXwCwuVWtXJ4fxXzwqiWdqWPnh4bfi8clCXZDmFU
2RpTDH0MxoU2yg5KCNg0NEMa7FnRg7B8lyB6WeOwUYvUsB0iGDfxhvtjMjxxkGklvh8Cswa/Jxdy
IjV9S4Q7y2DhTGi7Pg+1EfJqj0IMBrsnPsux1tHVBPAEoaIXz/IGNh07iNTg30xEWGzI7h/s/VQc
Ak9OnEFmVJbJdLS/q6QcR3VGhObfAVaMqwouT7Btq6fVIJqDIVa+NZcByQOoCzO8t10fbqGbcKcO
VJoObzQ26M9yygWwjlp6H/gjIC8WslYF+3G81AOomNZLF/TA9z13HiHFaKP+CXnYeOJc7aYlr7E3
NomBZ/3lT86LRn49UQ+qs7w7YM1HPnERs+lbD9DgrmJblx1k51UvHzK6UKLtb0t2SyLl7XmyTtNy
0YJfcoaTdlLZfT0uz6resdzKtpcH+sQNeTJswwYsTp3uBytorXyLOMKYDs4schMNMeS/ixg4TzlP
cK3NFpT9fTTkMZHDsPGw+HK3n3QltXmDsJOdwbQgDebgpDOd9cCDNQtRA/Fj9RLunBiUHVS/zWt7
8xIe2Ay6pWOwMuxhqpPhEb6mzTgDYDpSvJ0Orxyb//tAkgULI99xmPnsisY1/PuFnUw1aGFWXLqo
MTH3uhGzIpNjDn4Xct9i4AyQlSkPGrSj/+dTCXlwx/3N15fVM760WpuESPEu8EIdwvUB9Nk+erGj
i8RN7VUTKy+o0W+hMm4dgU4NX/byn2+Grapp+UhcKjSDF1Qw6GAwpbCZdzJunXIV8Ak3pfPRQvaT
GlDDteSdtA4v8hq1yHkaK0NpwrdEtulhNI5l8p9Q8i5cj1RAveMn4JSNnrfbkPT/eUx8Ef4n2KW4
uFKgU4Ct2LdEZC94BXBjMz56+f8SzP5Sld7+xqmd2ZIShz7QU75g5RMK3OVP8v8m/3wp5PYE48Am
qrBe08f728uWxIKkmpL1mjQ1wOvgeyLqvOA6uITKOlZK+g6Psk8RKzX0wjI5d5bYskZwS0Lh32cg
sssjqZZfd/YYtjovP3zHZzuEHyHlA/9UTN8xnl6YQQ5WOEFW/rhCzVxrznKV1gLHy+YsCNyURqHD
sA7tuxfZQczQpNj0cY9J8J8Sdq9fxMRf9Qwog0NVNuKr5Oex+UHOI0gFq8uGjnWMHJzmfwVJNNjC
JVqCdojIW6ae9IjSvI3O8gypT9woNpRwBeqJclYyb75ieF4paiGF9TI0pA1uBK11Oo5/imnB4azc
/PMHjeS5gksk9GYS7EPKBXvMrOVT66gQ6VXLm6rBN/xpCiR0KeKMoGN9tyelkqoJg/Wl4bIzPC01
Fxrx9BMFMH4fuKUzLMvego4gmgEOWUMYNu7PREqiOYQ+ZYFkJvn8TWQw9WHMQ77H8yLEbXRXxjXv
Ef81iWJ8Sb49jrttHRz0siKyowqLbhY4CrQqrcPEOBwGG3iW9Y2aXsMv5fi7gQ/fX9kN+ANnwOfR
bGhQ4gcu/4jcGN6PH6huRggVbQFjNfY+c5ufNuCdxSXKwuzHIEWBTg+bajxUtuOjX+oHXiTV31hL
1PUOamzQXdCKJoYRTFpD9+JH4P38sSAXD0m6EFeBV0ijB5Z/n2PPOaRQjQvo8NPLczvZId7w1DsG
gPy+lF9xS7fQhi3yvX63zjSJHjbidmOyuCwss40DzqGeDSIBe1TEswfs7U038kGj3fFkZw3jvxBQ
TrCw3hBorTQlMw1q8+pdYn4jatlYaDFgP9xmYkfUZSPZEU1aTXfLyW3XVFQvjt+1q8QEttpgABnp
ST968cmGQ8nTtldFD7Gu9e6ZeNHPuCzsCQn5OTYF5RkX1JRXi728V2E1YcbUEVgKwkXnPU4RUA20
84EIXO8Wd4qD3LqXxKDOHoAhWZ8PAIpNYUtcr9Ff/AY7r3LWnDn2HEwv6oWqz0283cfXgia0XSES
1oqgAWWRl6LsR2FsJxyXBEAgQJ6XWaohObFzEFBciAwNuPC55NxUXdQa3fwaScSLjBb+xGxE+dDX
jNZhc1ryi3y5VlLrjMCFPqjFV5wS7/7aLJ3JiOLRIwU7n44X5L/4zTa+Ig7UrT/Ucq1mU+lO07SR
2j0P/njRQJdApHEU3z/PMZVuobheva7aWIfA5Qo6kooNYjD+rlYg/yn5WrI+xZ+wFa6FDyVnG4Rc
rqSC1DpXJ9q7V6g8G+8MjZF7WVHCwDPBge8QXNZfO12DHjKHcjPEtARatYRivzeQ4WJKob8UFgfu
eE6lnVAM5Z0+dX+TUHLjONwb2VYW2SVY1MRGFsUWO3nZPKJ7zEm/TzqxpZLuVCHNpKtI5uvEQmBO
9v8CPk9nGzx93q0Z2Tz7IzLmQxrAeGW55oBZhzGoX/nNB3A9mjkIeOGbOibTYUBwq78OISr9OiGs
5fn84KcMEIEPPRefoIheFI42sq01RJ1412Lk66Pdl/FOxpJoxGGpsxBEoX/bWgeeUM//GAxsKWi0
wQY6FRBLHL5FZZKIf6ajVwOH3nNBbiRur3WHBHtfYCzd2oc2DN2OVDjv4kWM4LVe5CxXtWwJidFe
DPcGpYgSgxpWdbncVkWI5m6yS+F6Q+dF4ataN0ZyacvwnYc42wotfBPnxDlRu+KJ9+2nrD7mA/mQ
Xujao88ck0SWv5zjFw4VwqvuAuPMclskxhUVUeY5biG41Ef4QG2vPvlTKwYVPxtC1SOgX7V2Vgkx
Eb0JF47YZCbzilzFDxHc9MW4kePSVEEKmmpLvjNs2C4/rGq39JJ3eAXqo0YjEsNFZy6mw5W8tiyJ
kNIAzmsT/n40KkNDt3RcteRgJWDeJtkhEKI8/FmHmhXewOAYcVlDBLBeYMMIHP/wZ0Ut7aXfXGM8
U/KdcSbKzEbdFto/kos4wwi/IK2XX6EWZ5O4r2kP4fRhKDb57TKPk0h4Ukx+GLEBVQEm5pKVmMRM
1AIyZBRV+G0SWUspkJOnC1gGGP/H6MoH7D8l67Kq6fKK9kr7e2vIuVI1TLAbD51e0vAo4Nn/Iepi
Lt4md9LBkTvn+1LjlD/jMPNqna2uSLFE2Y834HraUxvcPoiNarpRWjwMmdfaYLizRTsT0h9nwV/G
HpAnIo+GOJL2gnqGUz9itEwwZAep17Yrrte9va2hJ2qC8Pv3LtGDvVTfuZqCEcXj5dXgWTOY/ulL
KzDiRA0G7qiax1fOPXfkhUMS2Stkn8w76m0BLUFhlfrQ9/PLhDJEU0hGwUBGe395fJkKk9YL8+te
etiikUK78fCn0iPoxETOIp272+cP9bTwZRH0B/G5cuOHGeHf5WKY1gST/NX+0NCrtv+U+T7eyNlr
8Zd9aRVyhHDRTaxMbQPLzaXFSV8FnH2pONGjubexwAZeQe91zhpCFfpIWXBAlp0RKSqk7xzHK5BS
WYkWEkA5G0uccJmS1iHRRyDKW+NkhfEEXNSf81qVDWWLpv03+hiuND75LE7WQ+wCl9KpJSjxy8BT
Qc+KB41gQ6r21jqc7paYBwdzeeNjklgh4xLDtawrM4qeDYRkXjuUNA3AhmnroZ1QIgjfLIUhvsWY
9qD3d4tLbHTs40qOrPTNUWFvc1Kj8ShlRBJ3YKCDYtJwROhDO/NDfIeZEFcKaGGaPmOZEa7t73Ni
Hk1Q4GWcfQP3aQ4TLfY/izWQRBR0LIfVT1UAe7577rlKiMIIiju6LLwvVPt4fVMN0YQFpzUEpc3v
DJeM+pUnYPGmU1m35haVoj9nVdnF9OXUKnSyW6X+4o+FlWcbxzAQw06au4sQUbQjighRQ1f6jTOn
e7vmWkmMBgyc9UUgIymYpEMUezMJby8J2I1cDVNA8Wd3e7UBHqeFtiyVWO/OyvaX7BT5Zdolzips
bnNOBaEQVSjzrIx64Y5Z7X39xuX+riPVSBS6oFGTWLovTrsR+5z/jNvHnAKUDNfQ15j7mSGWALPD
OF6P3XSWl9X9FS/mjsueUqgquMX85p9GYpPpTfmg7y/r6z2ekMgV/0RbpW/VmEz0qCtlIbMLfeVt
xL46EiJPmjYKCd42vGRaOBiiWrdKCP681r6nCGsM/qJFhHRcw+yEp5WeMtAe4xQQWDJ9VdZPw9OX
cmQG4UwPWm2SBRZoGSGiitozi83yHkuwGHaxCVZnNb1/O1tLeehYMUaSP2SSalVlqfKWI7ePLTGO
4I6X/zMKYJk4qAh1DvJdSVzA9tDWS+hiL6bQ/uw7HOu9XCRD/OfU0diCgm7PWbsQMs2XyISLjaZC
9tma9NDisQh0qQIOsBdU68U9ST+S7/5HjZI2LQWivuP4UfTNjSUpOm28O25A8AGd7+swsAlvaAu9
1H6Bk4CLx0IlhjSvJ+KhaA7TF+Gfgmwa2g/arxsbCPr+bq5IthWEvxmrTzJ1J815u7GtWTCcMRfX
1a5Gv2ougXY+y8SL366tjsk5DlQvzZJphU7EhMReN/7LndYNTzdMLpnn/jyGxZZJCh24RdFl38Jy
Zzs96ad8pNl6O0b4o26nKYU4m8qvSRlkqWVAOHmc8HPiSx3cm8ucIjCci+9xVUKgi2wiuFjk830G
ibeO2tFYbyLnB+mpaVT6epOyrBlbweQE9N2xCZdcRqOhaXlYXAPpc/fSWmHC7FHtEaRvAB2jI8x3
h/kWn7eOfVEAGDnAvLTFsZq6+tzhGaJcWB4K0/ebaOV85B2u8rli7PFPotcOUAd4A3Ltd2W39SUF
M21Qk0HmDd0XjFrCtJUl7sWcxmmcMTvncILwIK9P0JFf4j7tjm2NXPafJXMggLsQDJ4hEGpPq1Zj
VJ2UjEqACuH1te2sFioykRwlralUznlPPFLMn2YGCtHtzqd1KJA9lTs/oz8wfMdjWsbPmZ+ZCT4n
91bexAWFVhFWVZMiBo0R/l2MDN2go8xwDT8FSdzCOB8biZU2PpL5QjzUa3uSRNJT+aIhPTX4lN8C
paRGj90q8eo6Q/p29h8LtzW2bFNgF0whMf/w5d/oUDgSYWADWzPos5gTeqJ1XR0AFmZT3q2/FcnX
AYLRJhLjueiOYUgyhr1VLfQlvMaFRWRogrlDeEgqkoM78OllppRBTpkjPzrQeJ8TisEtO+Ayj1PW
2MN/0GaArvoirZYtrswmsxwP1AZpbz75xxKJv1CH+oENoFiIdKZdTdN8L1Gi6xJ3w5iR/CBx6p+v
nK+THBPSnckz0259Q1OjkYzdZaFkYu+38q7+r9Zoa0UQss+cfZAZkYQjxo6F7QYmDqWecKSo3SjK
yoaDEFA2GGmyPkpN5e2hTk2Gj/4r21Dq1i6/qrApNglozHN7t9SvjiNeT4/ajOZlvpWsxhhi6Wpq
JLVIOUjJJnUwchhWgf7581JpDnMi12ekzRdI96qUXaZoA89aqCE2cmzVJDgzeekA12MjUZHIWM9D
KQiLlJ0LTC5cng3cYRu3kSntrjTLmA9yf63p/ijxuWzKkXcqpThcE0AkdbkW1SXYreYHzUL473rp
XI06yko+7Iu6JV6EX0sSXc+1NfCzAcaSn9S86IsbPxySb7+F5QL+gW0W36Y7ES/k+OrRzXqMbuw1
pRAX2uZeQ6Os/muZYYNHfFpkIM/vwj10wfz2vGhlFrGYqCiAzcA13ZQUkzL4LmLb8xzYxSsOp7Xi
FBJJYawmlIHNbR/XUOicr824/BZoure5UyDL3/k4uffbDuWxAZ9Q3AabMlC1ajas2XVN4gbGEw1X
BNtcx8aBYhtexHqn2c3mon3nePEcFodem15Hh5w1eAfk1guUDKHj//qSvoEbryh3F9VFrIBLM1cx
mFRBeDYmWc+6ie/517GIidz8k1zDj3sBmhggj7HuZtb3pWKtAOadm74njcgbmoc1fnq/6NPBOcy1
MzjI1Y1xsBclR09KnCfSJmHE5MwFgc46Ja3ZtNJe8jjrOPneTqBDTtRzQLYRwh6KWy7qvNhhSahC
QD8BcsBSVmmls43mhXOOSGES9MyDklpx3XzdgQ9OHS5+40caDKSgTdKYzIiyHgbzM1qsoq0g5yTu
13XI8H19cTsMCTIR67fmNdhAl+g+eNp4K5MjYp38XZ8iTYUrM6LKLKiioL4zK3Hb9JMTlrNl9bo8
trM2jGl8BkhdxO/o0VognDI35ml1LOnVJnHQAuV4qSPKCbso3vEkCjcLz7gb4AOCulM8DNyu1T1N
4vlyHINMiF3UQLTcPD5FAPMe1q7tC8DAZm0MMAS3rxaLPb1OFzGEZYhpHdjwNFDYgNa8h3kQXxpf
o5+IjdM0L1D4GOzqQMd/EW5KGKVr2/mF9rqoHO4kM07yydEQTnD59Y6NwfM0t4JwBcaUkqEM5KeP
E5om9yyMrJYlJWypRtvjmXeepkDTYsP7gyU56PbICkePSyha8mborcooxFai0bZ87T18I9EDebp4
i3Eh/z6+ATSm6C0hitoJTIx7l2usM2gvo9fLbtME9TIXfxFhNhXeYKXYuizwvS27iKQrzRufqwVl
JilikCLWu5epd3J9qNuHnohUzW4x4/mYQHJ1q9eRcYZVnqTNgDsyQm9ilCBlvsYpimVnZqLIYZoC
eEm+ZrSTTm8NGMa4NZbkWkVAZ5F9aDZK1WM1snQS8nObInzXPQyFQsk7UEqujQhIBcIDQ2j/e1Rx
f0AAlN1avf5ko8doweknVMcq4HDzfiW2rjlwgjj6bvdeCMsQjf4NNk3d01mdiEIUZn9zHIUVV1xX
BaRaSW15DpjYT0WTJ7hTeJBDz+hxzMsKmgD6ioEOQJ7udhn090pSBX1Eh6D9+Xab5zk+elvkvPeN
0jA5eBG+ROFLK3KygDy28ibHgFRKpCMQ/r7390WqsYJRekaf3PkqWa7zuSVMov/pxhvYnTJZt6Dt
rFlhbA3JjWNpN6GdKWQwqBoVjXKIDnWr021CboMEzZZSnPJpF/+hSua70FhQqenIxhe5ZC9SDkNm
0U128vHLhjtD3nD+sIhgnYHh5bebPO5/fKSDji8cIiVhiwFVBMvukaiumjpqJjU+J1CTj+fAZkNu
a5b3GJAzyJ355jSKxP5uVka+IDazcxDrho6Lig22sZS0BbIN+GyDGxc4s3+yDffJeHRZzKbyxrJL
2Kdh+w3EGus8ieyS7EuMfx61pGLwzMhD4LCS6pTPb4V/+H+9IIeErGdibUmQdt6NVFAAxstLq88A
isNDLD5SzJZy965AnhBT+uH5JYt9SN7/5QF1m6+8Xj1F7RC0Xzz2rtHLvvgabNoEHSFLlhZNRpZ1
TgWsurfWmj5WmeToLFPwQ4/nteWxcRUlHIjhnFAg665xzArrjCHnwvvlv5//YM5Q/W1kSLj0lgtR
0pIR/mXromH/mHD9NSOkZueVS1uUR9fFrhjDhLsACFXARCB+H886/f660rjQu2i2hjE9xt5FqAdl
rPk2wfuFi3gMCHjXo4tvFKvyOA/zTu0uYNutV/CAu3sUt+Rp9XpZLETSJSEJXliYrKov7k9AoPn1
ftLh+V45LZb01Lk3joFAV4Fl8OzB29u7REvf4P1T4csqVdX0HaRRJarCiZpsuJedS3C+15+65KXs
nWbAbbS+59RQO04bc7YaE4EbSpdvlN/SOLc37/v3MWd84R+WwEhV/QpZZAkIeNK9SQwA4lVgKUhf
0mzgLKLmzZVJ67xEzDADmcNIPME7AiowQqsw1TaihGa+u/WBi5R91DwwGiaKQWI8saoR2/WVJcF6
MKSOdjw55bZSW8Vm5LYgj/O3/cevtW/15wqiJGAdNnPRnjFjFuSWgiLfoHLlT7nSxX4nJYgWNkFh
ccPQBnxIUT4p+vIoy5YDZLkhDGl6cHHxKRxk16D9bs5ammQinG4W+0uygue7MuRhBIHbHws3Y6Ag
kZAX+ZbbDkw7duTJZxBa1Gz1w5zpEgsH/urYKHGTrmiq9hbJ3+KcBfQoWA8lUWlgm6rjgO07S2bm
LUJV5tgBy48NQDQh4vaIPlmxheM0dS7bjwaOSXpOD+U7Emzlhh3CTRTVXnoy3EEEMNZgTcxckv4o
y/Or56HWxasG/jqEt8KpXfs1SuusKlJLECn/PtdwvjKIDLet68AZ+cNnCctne3kYAxPdd2a4THGx
7hsj5T6rabYct8vr78yTpAm+99kF4zsQkPmLlE3K89alKnPjavZOyW7Iu+rma04ttKKNbrh3KKiE
35WdPUB2UcVPt4L2NOk4jNKbXrAKwhyDmEw7yfDvpceuNK0PQBnpSGXKd0QdeeIVWNQ6ri2/GyHC
mypEjpzVjT2P/FFML+FXBrDXfYNdPlxgucq02fVcKa6QKU4l6U5M9rTCvepkeoSDfXfqT5WGclrP
8nXiXkLG5C1MDk56wc5H455X8XmUJq+TPNWzEFhXUDHConn6RypB28jeQ/BSIN/7RDagM/QboxYC
HKFeTdx+ZwbZzlaWRiKniuvfY3L5pczspG4ODXUZjhKO17Pma1+dA966/plKHrwxTmB/sOXuVTf2
X8aAks14tSMs+GakgtPJlgSAOKePQaHOSNjln/r3zchd8QlfvoOoFD8MakqIrCZ8aysybwMHXd+h
vL/NBNkZnGJxpHGfH4CxQuv6F+1vsBqGtAPRFpyDCNonQI17kS2KeOfI41ZAmjiFPI6TsEb4sQl/
UN/oF3baEDpC+SvmxBjZSifKvT7/BYkTsjt1wIUR5NH/RpJC63RtwpB9DHG3KzfNoK7grw2Q1xta
jkcyHudKy+jpknbwbPEtjLuKCYuDIpopxKLXPU6wSVPspLGXoY7oDt2mAOqKBby5ia31iFh0vb+Y
a3DfbsTxOM+bXoNxu/pfkSgHHJvzPcadszf/UZxtTOggtJuIeCtRzLorWqT3qEYnDdYcy8qf3ORm
R62uCrcfIiVhqrAip9RPDaNBGARinDJ7kBbu909OeYqC/6EDdDptjS0oKgNscWhYxQCqYBgC9BTa
eoWwtCVpMOCvsu2eZVPDtR995YHNL2bsm8xP0fEkUqyQbieUOVT52ptRz/EPOCjl/grQhaqUKglb
fa1iNVTo0l81l33vTrBNLgjB6j4nbP9XgDu81XkdQ92p9UyRzLRvxokcagilhPhGNNHcqbKUSOeg
EKncYnDkT3LeU7YQ1hDECSTliYgOGq57DSOOXb2Ffb5waMSm+UCTLP3nxjfE5GxeeJ4ex1vNAEV9
cg7wzU68fk0aG99FAUmgpyE72/dXJBjbp9Iq95Ju1GqoWNWE3P5XFh8B1IJyUig7dIrMJ8LWdhuj
dMd8EmL361qQ1/1Jai1NCnNSPklBGDhWRVqBFLFXHpE2W2DZZfEvWIzKOvSwS4w7hTQXd6KNsfCi
dRBLaQFPGKF09nHv62hKHJIZp3wRMQbduDutpaBEuACzmqa3OCYbWpBMaNptQUcLcu+UtJPyvodA
Pyi+ka8Oid5mSwXJvYYuKqzOE+i9/cLFpHkkL+q/nYKUtmy40JCI2HSBPHzjgxq34SCR9onpTp2C
gNXBo4PSIOyh7GTfJeMkP5qjHktYh6Vglg+esivGG91clU3PEFRcbWJBgc5gIdYm8nyAcb02Qsva
uIokvM2r1Q8+SdM/HWXcj9RbcLxFk9c3tQzlEWolmrtKPnNIjyCmgsm5iC3WPCtuC5Sb4ascapXU
O6jTj6IKKn/VnyXwigIcXj5AM/3rTRBqyKohMudSJODP6fum3Ncl/8dKwvcVnlgfvLIvmzrX6uQg
IpMLh7kmDOTz5+ULePg3lYeA5crf7mHrmMJ+kgWvhXf2GoCIT5n/zmftTpug+VMYM6qobRNaS+8M
1apF9ix5ie7GIOA6jpEgXg00sV3f4uEu6rnhdSsc7OLG/HR+HHbMOxsnS/TresPFFOjKP9HMfy19
bp3J2KiytbwiWw147GkutCalmWua8ySoxC+Wpjid/UR3VH9rPf7c6Rodb0oLzPkofyBnslL1F16G
fPgW1Smbtuwf6KZNcRQzbrwBxIWyVjbWu4yCxjJInJCgTi8uJdW6Z33bZTsOqUdLJr97DtfgRd+N
gVL72cXbyNatxbRMGgqk+VNO8xgJHn9Nq5EdutrExew7rsLBu506VRV76pd+EUYRDxaHiaK0cLLC
Hnzfnu9G47aVwN13KkOQmNbdLqromY4S5GibzCujz3IjIV6WYC6RJooBM0vPCxGxLJ0HeCLUpsWU
QJow2XhCiGIYzMwFQNBL0DzVI05EL4eZiisvaT4GP2LIdSaIw30evE/Ie0y/8mbHvxbrlREBd/gC
sFA0lpLOppzlQ8NqfMMg1bbCY1csalvng9cRCeFjbrP7SqTxajfiRJBQE9W38gm6ibn6si+s8AZP
Qf23IvgWs95+rdDPNtjCJo0bQ39ViybGgb8cnKh9GBHks5yrhNxKXQCDIyEatoE0PnSq9vmGlqpf
O7bpj22xuZnim4aotfCYVYrkGdxQKOmd/MrTNcoS2YYvACzsqu4k0SFmvu3cCfbTb/tSrhx0DXJN
Ba0ks0IflEiLAHwzuWxttGxo2ZWez5Jj0x8Mrdol615l6GQSFTxXe1vmYURP7g0M9GGaCg0t2FWW
tiMIBTF1WAUfxuMyJ+AIxzTcfgh1oQels8Ks2+IgiHWaJu7VOIwsM6sz7BtjbsdoqeDOJtMp0GO7
0Dvq/benjpsTLVwazJz/XqZWecmbv5lFzhgSJtYM4/ivfhDEEiod73Dfs2WwWcN5LmhNxtpGWMXe
+QBW0EQ4otPeKLbo7HdsMxBZ2Q1Uv6ohEOU81NKUizgBlx8a7SSzt+h8+Z0klIMVqauv3Z+ST99c
klyHPOxnX6ee+1KJTW96sHDoM8xIpvn6DhjeulNl6sH12YhvGRqewkkQaoFUcYVZKa0ep8jpFSx3
iEKOA1TPN8sBBGiuXtSjYU2myKAMhMHKsfxtXpu7KSOdY+LlP/czP/L++Ib4wFz3h4QByrmhKeGR
qYf/KhTAKMAUNWlcgKTgr3aN7nAZxbogb3qyMN0SS9SDu+iqD5rF+aHctTG+kf6iNGymERHIFBE5
feE/CEitoyn79Q35m1fFV7Buo/A82ZelDjcKruVFMzkhNCZohy4mqdDLZRcdQwuSW9PLeHeNNLCs
0xSjITmxtpoB7jDWOUGWH0QyQoBHDNLyVOLLs7M4lxS8xU1YjD8VmNoM4qn7co7t02NlCLw0WMJC
jUQEECoji9VFRIycEZgD+fOWQsyWWxHwv3ccQGW2py+nGd/vJ5GN4LtK7SMGvRNNzTY5HQUIUBY5
8qDjJggMa+R1q0kBkjBp0ex0vP7sithskCag8L+DhSHJJKE99plgqYgS64Y2Uk2yPbX/5D3vyFGh
A+k+bLUalfIoAIjWZRrlkxCyp/MYy3VEYzU7vVg/rTlTJsixe5wTBiP+3NLV1I6r5XA8pt4m6gqZ
vMcROjdZnEye6fZWMqbKZhqkiwGaXYno7BbxY/skMgdjXBOAadj3im/Gpqav+hBcFKUs9NxGsls8
C+QSx41sFphqdA0lGgXTT0uNuoB5TasmXuVmM13NobfIwoYnw9l5R2HRlPMJuolFkVbjHDYzbX/C
yCYAx8n/lK0gwNEcC0kEnl+Z+LfrW5zUyhQy8fUaaXToftCTNkHqvdEqCFEgBsaFXm6Hmotz6czT
MZMS7nW/ImJz5IIZOoxrvCmh3LJUIS+2KzEAx+f0HEdsJxvEC6u12sGKyS/C0INdRio60dZ2c1g7
l5+kA3RFcI2y63Ih3tgMeNDjUZh38rc2+6Nm0lZ430aZVFzdbLde0RoM30vP9tc+adYMzpPNpo9n
uCFtpYLBsvDyCvqj+UZgP/Y2ZvDbctJeDbG076eeclOd/e8pHdaB2Dax30++r2fTFixiG6YE2M2e
oZI5GcXxpNEi2ECXq+rSq6+QMzrjB11Z0nimsAo2hAgYBufF5e6TUonTvkqL+7iet70yzWJlI/IO
uxeHyABfJaj/56+P9P1XSIbWyNku7Ub2hqd9XD13R3GgkYyOxnegUd0PuaEVeLEesCvcsy6wYNvv
8Hp8SN7mD3d2/DuHINGlcW1l/7my/bAKdDdcde8TQqCnWU89E/1ZWMWTMNQb1JrvFGNmsxhKj2zj
1e5IidrrbZt2ZQfyq0T8AW0foUCxlSC6DxI5xbC0qJ/AXYSe+D6huGcMxmjb6i7qn7Ndhn6aZx+B
ct+CdqycYZydgpfU3P3hKD/PxVD8exMyYDEnJ2B2hyNtSRTpqhX2eay+iTjwXwhQEiOwhisR6axk
kHsctoTMfOgNAdY2WXk/EmxVfI9fJHwNqDXE6iwHH3wCvllmjUPXZSz7ZqQTxwrlzFTuNIA6dHC2
8SYFEPXNxquyQ8yXMZSxhoDdM9hnAc4GKO9yMRWqkP5YNk4RjlCMWhiesgXlES3H4TVUPMvK0HOR
ZuShGl5bPGpblYL8+KUXaYxUz9goCkGn+Jzt6n8btRxwac2vU6iUzwOJpDSpd3z9xGP1vreYR3az
Ll6mTtaTguK3AzAVi7toHfIoAEQEGIixJ3DXYxj0i4YTmv2nTDERDvPEyLC+aycHER2UMutm/lI2
wwDAjtgoIrQgqiwOgxuGax5MKPcN+CNdsMLvte8u5xq7s/haXN6g+SWc1VcgK3EDSgu9BrZ4VaF7
u18AHFkN90MAU5XZPb5LPCZZ+pMKr7cAGkMqcB8ig0ZRlJee5UAUHGspjXjNQwwsg+QWFqh9R/5M
GbyYB3db/oqWhnfYY0r9XKVfbzM8TcRVmo7tPBxCXgtfMDQr0cNAr8nNYVO+ghhZ5ntQTz08W22s
00q7Uy0BPY7J8Jc8z31xCAoRYRrTYaFsDyd/UvZ/Kp4jQJWbkS5IBzc1pEZ65ft1qhMfjexWPyNn
NrBdQYkMJ1Q1rjxBBxVovWDpPC1P30xO78L3qMY06GGrrH6kalkeyRIBpIxnPhfNGEmqD/Hx8+jk
Ko4n1HONamaAXg8OrgacITUpkDGccnE6f1VIln+llktldS2yfItoUedUGUruVDMpFE5n0jWtFeCs
Qsa9mlsdBPyCYSau+htxolWTJ3u4Bi/eFLKNxsO72EzY/Dg0dhotP/dItQWxOOTTmdWgp+wvYvt6
UoqXKMHI1a0Cnwtag0CCo3mvO30uLHwzNnvdGPiRVmZoRbCsBOoLHOqcBxbbySerj/7BeDyqy4UQ
PUr8Z0yczi9BApwsd/DK8OPJeKJHkyQaE3n+1/0ZEjKjZMeqbhUoSeo1uhudV/VqPe0t8Rkkc47t
RyN7DpWuHJBWo2qkN9nnqbR88GTG3+D05uxf/tfwBLaeJdTT9F4eq/XbXirIzhs+1vHVgn3nnJ/H
kUEF0B8C8jKzMI8mN2B+I92F7KSYihA8RPE27lQDQkH58takoXyMw2sYdbBSXVfkoV4kxIB4EwxA
SXkVmOFj9Nmd2AX4LTrnEFcqpxJk0o9Ne72ZDuAF4z+EIltdr5OwSqB99TftkMB+NQIdvKw9yUgU
nHhEIK4ndkMfODg+c/2nU20Ekj/k3SfwhjTWV/b38QXVAdZyTxnzv9z8al3L4itZJ0cSmHDbwFE4
TrLRN8RH/ef/bE20PfVJY/h1QUjig3ukLfWeJttSbwL+hf87l7xGvhDLlyeajOvGkY3eeUTRTD6i
aNsvVF0lcSfmTJ4PlIJn7nYSO32GY//hf0fFsV0xkzBNnPmi5exR9R64GMxlLZqZdIDp+dnhXcNo
GjvdrihpNL0LFgxAFYpX9CFV+ybrbwTLktAZbZX/ZF/dpy+jYea92IXStDW0K3BY/eKHlex0vfSu
5MK3848OHVX2NZRsr/6FRe2ea7hEInVy8ZrZ+U5MJA6aWr6eZjIw3U+ABIWbfuW/S5B+QYC/Lyl1
soaUJH6pBbKsLOoBnYwwXBXp7VNEtM0pbwN1i1Qct+EFqUIdo9IVfiJSAGlK4p7Dzc7zIOYsPr99
uEQmuXw+IjCv0bB+E4ypVfg5ki3jEBcuNW3ZWX1+4cHYMOJza2vs+aXCx4HeJjc3Du+oG7VB1DLT
vcyHeC/7uHEUDRv4wWIw+/jM6x+KLAtVpuH0KcLtlnlsO0ItAYC6fv9G0B1rsdp7gbVJyykjsJKO
afN4QBUtsHo/Sz+9ud0ZH7updVcunxz7tgK1xWkmANdc0ZMPdIzw0iMizDLWdaP+BUBSYOYB9mGw
KEiypVS2XhCmPD1KqUePZMRgyWsU0EgZTYEcNUg3Q+G6c7MDJlMgU7oX0rwpxP1TZAtlK0hJaHhX
td0PtZjO7cjAQvfR0B0p6ImQGL5Rc8zWgLuDqBwAQpnhTzFriwbNxjcO79DetBHZ6z2cuDPG1ouV
w+Xm7JKv30XT/+VvGU0N/o7JuUgen05DBQEm/u2MyRnYDY77+pvjy6ONzVRYFI5oVnGdt30W7pOV
wzbGzU6SeBu2JoXV94YJoN0/a4yttgsf4w55eVxDVlLmuu3R2ZWhleQllPTOtTqIYT4QY6y79XES
Ybc3Gh39hKmXrH5ZZsQ8Aih/1ydAyD0zPVaJj54rOOnLv53IBEhW0cGwefTuRPF/1Ws3AyFXNZG2
N5IU0MtIWNcVXWylTiDHR1T57GBnjPqyiXN4JRrv6fJKr/zl3vW4btMKp6eNdFNtGx7TJGXmW8KN
xiGM85ekBIU3d9dmWKSv76Q/UxcH8qC0j0/royRUg+iOWP0UNs8qSLeo2qo5sojVJDGWr4RDpaP6
N4/k5cKEG8l6/bvIQroaOZx7BUfXB3HtzZLUMb1fBWy4e2gY+uZWO59hw4iw/Y9ercbf5wBveThX
elKThREJSoZNf3DTpLK2Khqrz+VJVpdAGIRj6dTDiZjwajcNpcxItZmhj+d0hqYWTnBiYoE84hd9
r0YGjBrcZrh1s7eZi55ZJmOB+/jixiEBPvt/Q6hpTQE1O36SwpUm/acbnU5a2JSE1lJszzXl/0K2
nCHkhOplkl6cZdtki0A2AsN0Quo55yn5bYmQGnUlScSlZ7M+m1aQ2SazoNdyQ4WGlgzdLmkkdL4F
YC/iRMNyqXADR23F4pIY5AAOFs8T1VbmEABPPvOH/G580LabCiWPFm8djf2TfHSERIQVDoi8p2MC
6v6qxuD4KAnIiGmj1DdD9cv2L5ZnOr3rUVQmhcmohuaBluKQI08NbtJeCrwuo5o7k47ecE5O1qvk
9q3KUTI/5aWQ7exClIIW4A6KHr+pFaqG7Ct76GHttlK7TGLtPgRtbypEt+IIiY70YYBejh6SecQj
5694+1EI3Gu/F4dlamLnGVyvHDJr5WTwAOjiqgOnM+59QwmPH/yv3XRVqlkCoXxEoWO0c0QZaKtp
bhTvnXL7Nl8QVRfqZ2ByvWV/jfQLCypw2UPBKB/zoj8xxDrw05TfEItdiYG2MxIxKo5KhfdijY6p
Bkrt8uEMFcrVJOFG0vuqrXs2b9cdOa8IXVseSftPO+OsIyw3Ve1fx0TVrZGTMxWf9Q4wOr0Ik5yM
fdFvxREoUmM/ctB8UJVwGc25oOioe7A3MM2GXHAZmT/NAYo9IU90jelZiGV/7aCnmseFnbN4jf+p
Xz+/L38BQ9F2zlQ4U2BJlSPN+DsdkgRmwh3KiISfiMOmmxs9KwChWXy0RPtCyC5L+cbRQys9aqMB
tGRUEE6fI4TSnMdwrjMjAd7n4aOMcxIiODjGPd4EcUczYEU6oe8OkAXjVpDjgqUZmHK6KUnnu6Mx
OUdEhgve3HNJ7Iod0DIvEYXX7KOsmGW6yHcgdfSvcYIYmdmNpXmx05epJP0X3jnpe8Mmw+RdWMGx
Qm4feXNi3gYzSuS+5aIU5GrSmxEiTOooMWRYA6l4nCZhY/pBwjfifLCZIEOS3Bmn7w8zAL11NYnX
D+DZ9gfKKenEWd6oY66Fqzb3OtZs4yrExyOjNl5XqGTcTbob2BYOKaa0eHmzKASUaOyPUUBUINx8
wMlRlGrNHl2CRoSPfLo8P2VR5IyJ0hStYSBZP2yiE95Uwt7AtKkTICN2E5xuAE/VLWG5r62SFl/u
rMPzYs94ZTyHq4WCBK67Cmhrd8cEH+kVzl7p8kFBgeD5rMD+kUcdO/OySGF+dU/w/1eAD4G1R+Y2
j03QeMe/aJy0hxm47Fsv9YVxBWNX35YAxgEfuUl+sB2OE/RuCLj1ywIFK4B2KMl5ejdUMSoKFzbA
jGeSxH/4iNrna7DcRqCDSXGaZJb9rGTj9RuLyfnp063P74G4QXiigHFe2KunoqDR/X5/KU9Y7C8v
PQHoWLDOGACHBIzyALVPIT90061I53UsIVAcdXx/5yfeMUimuJuByX+yszyXoEzWFdROHTLTqjJK
w8JxvYx44CRtkSsSJNvXmZrtQIx8BdbPLFpGTdfLCH1u2M30RxxDXMm2hzTyRC9h8wiojapBj1VE
pkKLLIXhGhrT+Us4/Uf1ZK5CRZCvVJWm8x8hywmo0+oaE8+rwGvKUM42CZVBVeNVzqgwg4kWiuWZ
bYtQC5Y5scTnMXS0KDtMzb21DnFQnEZunr23XX/33AAEzn/LkqhGtuobuE3MJUFMcvHwoyhcNa9P
hQxnLOh/MYufPUgA4anx1gndyB4fheXwYXb22jkxXsFZ/wUakdHKI1ntkm3P5m8aSyJIkaZPJ3v1
cq+2j6q/VbE2V7ovS97PVqdY09NARHxwz4jlXuYvHkhc/ZP4OAPqab162YEZ/sdAXepOyul8m+LE
EJbOYiA129QPyZjD/lRcIwYrloJcwsTky8q4lw/AyY0zwhVi0s7paRw51FACRv829b2J9H3v0K1C
lwyk+tLH2+bwRZAxcV5oio1pzV8VF9eblwOsPtGOxrzW8Ry5ow3PSCtkWD3LGo3LDj8XYpKJpCfi
QyXM/L6AdA0dFVNHvtM+uj3niliv5SYwIbVP2tXZoH2PnZM3QEr6mc7RASCCmAPVXPhkL1W2m+eD
Giz9dGD/GX46+zDY/N6homhEkxmUt57Wpuc0GEuYGRrjMwKDfMQqMzd09DRECIrDmqH0EaUeHVTB
e9yPUCNvjnYLvRkZEBuW7Jh76sXsc/BGoH70+H73YcHUWhBQnLGSYRrDG/2rd+n9FGlD3TE2rIuh
58HDgxJ1uarzxptH+ZfQFXeNlKIFK0bJ9SLwsvjicfHj0TKRAe1S1SN9oBfCQgRpPfXEXvJtaW+Q
DtNU0f+N+Z5Pg0WHlSWjmUwKbfdpugAvjspHWm9wmvFumDGObGU7YsiA1cFwiz1yhNbMUQtbEpfs
jXMWNkTGiqnUbeIBi0h2iPx/5lhRGgPhlAxyjCXuE2KcAsVbgUVTUOkJt9WDiGMxnvlWwof2D4ED
ient3vy9pBjTTPUrC5Bx1SZv3jKKkA0FoLhOL6ep+2FeIh5+c1m0KQd7SYJHgpUb59cNiaSectAf
00cbSAmGZ1wi70Ze8PV3p6uPii3U2nODTvBYrJjosgCZ8dAJ+cUtzhiBS0Dywzc+cNT0fOvbkEJE
81wc8/kN+qrTA4ua3aFhDe22LgeSKF2sAFXfnF6JEvy4mX1xJLVyVqXLTo3Ea/OeyBqnmxTbeWBY
HySR7NpFffOgbRvrKWzkJKI4C2uCXT1p+uQ68CV4cac2sorEY9HbPwCeHhZtrOEuUc+f0Ldzov+i
01rZaCf/tk7VY44Y1h3wrhfurOwotnilwBc5v6b6BFjd2w/89T6uMpmFY6m2ksN8JWi5/4ZlNm/m
vjcPGq/8ilb2AalOlVo/eZp4BV4g7GJEOQrmMhbS8A1vbtQOhUgkAvVeb7L/UY65pAMtoqPiI2oS
pMR6RQPikR4uuVTxCnxPhrC6GZW/s4yOXuEBv8lfuq8dNBiulsZJqOjZb/JBStBd/aBAIheLf4SU
mMm1iIj+8/fx4Z2Js+OD7u5rYxZ6zvG38DvLBA29DY0jBmBMYT/Tc63isK6O1myfAYv2Mu8rsvYO
I6JDemkZwIBpWXthPOLywp2rGOniNVMejwSena06Q6BJo5SZCdJWf9Ar6HJ5E8xAUGlNmwRdrH5i
Cg8EMlvZWjX3OzK6msvQNN2DMYhZX0jXzyvsuep/AE9hXsfZcZhX1xj4vXKTWiiAVUczGWR6d4CN
1eNUfHD83SJDbZytrv70kUTQTKlAO/nkAeg+6g7zxVkP0UiEhITdedAn5I5+9r829UXDiavOCfIv
d0t2lEE1sJRJicpJm6XfqejCvN6m7cvbj7je9TP7oSH9rPUu7Y7QkC3+DjcRUXkFg0Zuu6L9HeoS
20csha5EpsfeRBLkEfQVGzjaiIK8z6nJXi7JEMpNYUleLwOuP7SPzS+6b2JjwpkuY1itqTV5kewm
vVDW3aAjMgNEvdV7AQOCjZIOo6icFPtRt6BMz2H9VdAhD1L1ModL6TPpwppb5NmH0XoDAu4Is4vb
Ypfuwmpihvz4EjVapVxLhSGRCnmlK/o6iM5tDNFrK/QQgsDYs/0VNp7leb+D8EsF5Ac5GjN8kElP
wIf1Ih7Hosv3zIP8bWnl/DyvZX9/g8W+dx7m9n6/A3dMZL8nJk2XepwEhOtb2B6Cj34nWh4yO6RA
JFpY8atVm7r71Ft0LF3fxG04GADRqtlIEOI3x1RVILFlow5+K9n7PN30UFCcB98cPW/kKbtB1i1w
7Kw2tGYvsRIumVTBs7HBerU+PnqsnP9aF+sZR7Qh6k68WpM/g0YNMVTrrgSwKTAWekGZWJOWOBxP
QHaMMc0V8ImIgxhWD6E8Fa7JSRdWdkDzeZ3P2Z77MkMaWbx8yyjA3Eitp7Du9AI2GjbtWmVLx5et
vosbKNm2srq95C5o5aTSg2iWIp8sP69eblnI18094SvBqtHJajkKwQwtg2OSSeFfDT7eU+0DX4r8
tiPbENB5aTXezsrHSpgH3QjSG4cQMIXUqNjTBS6xa4UOuGuXRBX4nk0mHpb39bEOwrRPRcfMI1pB
6aWqwNvNwrIZrxJwe9YNkpMFbljrT211d1OoKwrwNN/ubrIuphppGTFgFLuo+qop2qraGKqbLNS/
ahZSTBoWt3KQxJWGVSoa/dqmEkW0MEpeLrqX7vB/8MvJWh2tw31yTdHPrW/+Pn+6I7vQy4OzdDiZ
5SP0QpHWGrOO/cxg3tVICZHjPoO7BMdl07IDUjoUZG/yhywBiLVkaicR3MICoGsS9/+Dysx+zgya
3KfAkS++HxQKxhUNaFLMitcPiDW2JzoKdFwJe8lU2NzPm3lIhSgN4CsxGRrz1rrdfupQCLlsvFNr
tEXaHi8Oi6CFwX682778MfPqDqmheWXvhz7bjMBqUB7IJl++AWVs3JwZVMWESFPEayyXGmHAVLP5
6ePotYtfmNz6Jb8YjFd9IeUROIDr1kbZC2zZpo4uAvq5ByWyj0cvGzLRpjW7NdjxX1pT6m7Zekts
1SbQXbTqBBeuoeO9rxPZBubXIpcvi9HLTMvR/yp/fhBtIF33ZVf1yN6HcmbOmhY0USa9qHfqt3uK
46T0pwjiVHiWaI1dkXKePFHUIPfLI/X4jpqgFlTzlfgMNMHLgzYCBRkpz9iKiPyVoAHh9d1vyfkB
p4qeeeGgW+rPA+0E/yuwtJIy7vzLvKTWS5I+VbutIk8PmoK6MD8Fwo83hVkYVe/Ah7JzlQLAB6y+
ntNnFdeCcJ69Y/PLKCFcdyWvwlgYFVAVDfjMYGYAUMRoLg9yF/riSXgUO5Ry6XbBGRNAvYJhPSsF
XVIVpfkZixWIt1ImPp9Tjqfsi5KYIL+PoyRBzT2xUWXRRlAyQtTS5sa+AGSHxLADlO5Z+1OT+wwu
99frvfULFYyQZ9jA7Z/ral/ifndDjvDDR0RTH6sJ9c97jgLqRs2RtYIf0UMDS/WszNXhIS2BwF0N
6zVpHaIOCHnACPfiY5/jXXdFWkqn142QosfPqi8n9RG6tmfEuJX9OHUlL6gldeasdvfz6D5dPnWw
PB7JJviYfaRgrH9McRCRyV17Un+AoYwEa2OhmDUD36rYY/J6ipMhFw5OlRqEjw2KSMC0sptDCLR2
9U/cK7PNoSQ/ktFAWyqsERMQI1mkqy1vuABrC1Mxqz65G3oi842Dzg6mJi2c1re2VZmpR4QvE64T
dsYd96DFXKmlVEWXTLAw1MkrCzPCKhNZ+pHKL3ACXdRKHKBDZv4pef3jtPKaL4irobVfDcA7vFHt
QAKEluRjdwLxwngMzHABbAKXzdRx+v/Eeg3WofkTHCtC7B1fBwxoBUUzgMBb5pdYWcQeNeuR5Uqu
B9TQKk0LMyHFXob2RMvNi2a9OZ+lkCI7rVGH5VnF4FMYr/ZbC+Ycf1xkHW5TSUo/+NbE5W8Ve/Xw
SgbFPr64niACwR0VJk/fMqenjYugxWVsjcxi9ch21pd9wdl9yCOWtoUpPpXpAHCe5TBE6R8VCsYa
DDcmw8NmlmoRsacIeMFYkY0LPlJVCcoK+Zg5g7F6OU6BErjip292bxA3RnQvmL2HZZxY7MyvAh3b
GIoqfHXy+BrDxL0r1d0MIU9iYQ+NTTQrVEBh/5aZ3Kq8/ApdKjHdtBq9qeywMwS+mKZdDf1f2132
xQZ5K1dtll4u6l7F/SNkt5YByQhBf6R+PiiyYLuwQIi+p2r5Pou814l5rrNVA/NX+Pno/qxmSlzn
8vky6QjT7QRJZR9kiA9oL5/3pWYG32+ps+Y3pi0Oqhm6L2TvVIlAFcbD+Md+c1K+1UtD3wAlxhYU
tDkuK0wNvLfcL400mW8Ruty+AZ9CBGnC1YWOKN2WjtSMNN/814WLQ4DKJjrux3Jvwgz5omXB2bED
qGv+RSDO7JLd8e/3n3BMPeMomUz/6CZf+TtAmUNEd5VpXh6ykvKyZmMBwaRJXSpUbcMNwt6bPIPD
T/txwlWQVK3sc6rBt/TmY23QPxWOOD/bWZJzwGqb3T6mr7ooqpRnzVv9+pPwH9C/+1Z6qtMw3n2h
hGW3l8qSfeStD1err3FQKA7NS6d+TXn3nl3Hpc/ZI4MtbvPB3tg1y0pNV067OQZxp+4O87EqRFrX
M3PALl/kaG/Dyn7u63PK1uzACzNeKdCoAxEswh+P+mms784wkpzGlKiXkeDv/tWkT23CpR/Van8Y
78zX+abKdovhvCE9Ccb+lLg402KE1zfkh6b5dwCHVjlM7Ej5O8eHdx6bBMTp3sbLUkanhHIDS6a8
W0FUVs4aPH2fIzMk+MR56n9eeZaFDaLf4JX7UbppOyOylA96TDI+9aWDbCctQLQzOYvxZRjExvlU
nRR24sSb+h09pGVoFCsf9r1LYm1GZOc7xEX5Oz7XVZlm1K+CNg0Z24lVIzB+a7dapSYRbLBPAIFZ
CfbAFql1gMB+tIUMnCmgTVFKGeWGkEIMEaXksLKQRtiKvf3PY8IB7DDpqVUsujBL1KW/ezxWc7eS
6nmkencQ5MHk1UB5+Zt0kzFfRbjaZemVM561iHYPJXl9LLCyWaaOHvBRUX2beZXL5CdkxfNabl83
S0ekDnlf0rdxJfiqRKzbZHCZpZIR0GL1rIv4qI4dVssxcWoWuTuW4JbEYqLnYMhCI3jhjcem4V/q
tpcc9QdV0b/aPm+1hdZYYY+dpPTK1bLfGqzZVqkPWeNq1CH4zKwm7u5Lyg05qifLcC6vd44C8q0S
JtxPCzdyBCciiKzTdMRKbRF/3hYhRhli6cIcpc1ygEbxLEl+/GeA8jvoPn1Pf04OyLlNv8FYBPBU
5uECxvI8tiZ3/XHW+AZRHDRMp7g9j9fm1TD3jOIcsocjN/mQ9qomo8r1t19myS5TKmsgBSiWMNg/
yg3N8INB4OlWDP6C9g13eqaM+dj35Kg85zyCEPGLZMYssDp6+x4zUNioQbYdpRRO97fOT4ofbf/1
4h0c0LQy1vwsPEPC/+lTg3av5q8G5KCYkFO12c4mo+XIrJh49qnRLN4NVFvpXzC9UrAzwc83cSB2
ETyldDDFwEOZYdqEafDspx+6HM1Vzdbw5jgre3weRFq1VDNPqTo9/mXOtRE1eigJPiOjX4VCmnBG
p9Mr+4iTN+xLTp7A2d/kAfiWDKV4ms1c/JQKUSbZmcjZWm8TVSDheSS/OxqNSBxi8riC9gOs70V7
E5F4z7w42jXWYQPn3X/g+1cQBNYUYWjmQZATvs3bIGyYiVUwOy5ZCwRGGyJrTVX+didDdGARHguW
R0KcBhUm4SjCw94JU/f7W5IRYhyx5/Ta2FgsKBA9Tmic8UbnRt8xQZjU70aYcEFZ0+4Zb7428C6R
71f09/OXmhqjeSeKoft58kE/baQRddUN+fofioGXhTRKH7ItUYY+CUfbXqZW9XYNg+oemcYDSr3l
zcIRJ5dMYEkFeDWMCrgs9mWRb16pUi8BDhRlO5JuhxbJxy9iFsMzLTPQcdQQRL0iZZu4AA5Tl5Kf
8Mo4FmzwEcJlGRJSLArbdrjYHsZ4YVGNb+GV6wIa5XwByuVYC0K/SIhAb+GoNyO7/uNj1+d0wI53
ki2t3vHXNOkoe7tPJ2zaPTVcGYeUvwDKWlYGNFzYyIkCyHb3cQ4aI8LdvmjilP11F/SgXq4fGLGr
UoGgf565+MwhK8M+sxFnfUXF4WqErIZ7pe775QZkYQtGEeP9iQro9P3ezikSilqQy3Tz40Troblg
GF+rMg0rs73KzhQVb/1eYTHwfnGFJgcG8xrupFSMK+1gvM3Xpxg4EfVhL2f09N7dfF9hXFAcgQOf
d/P7eDlyNblmOmzuFYd/jCtCUCWgHtyyzueHlKakVuloG/O3GBOqmghCctdkBbuJaJxRCbMrGQj+
AAq273GYK0ocMHOQiIWtkp3rRGExuvxbNnIu4gIdYIc8535hOrJy90LKEGSwWideBAZvvDPhxHmj
y8TR5/YiovmJbqd1XBK4QvQB5aGboNw0zMFG7ThoGniOuTf8kikzTQyCjkv097EmpaPEubw2/uHQ
uqQuUJhytj4SbJ98hTuENMQrXCPg92+DcEom93mM9fNT2nLY83QxJx4e4IGZrB8t8/fFSTopjDTH
A1oNLxfoa/akEBKqSx4DZ8JyqUOc9N2Yg1jmD0YkcKOBTLCY1r8byRK+r2Woe6WImt77hgve+3U/
oa5/lsbE1yNyrl+/mb++B8FdmxIQOlK3anwR0znHZqnUVR4TQMndDkPG/T/dnjjy9EtOBwEOxmrl
AiZHvUSaPA03O1xPpRLDd5IJ+VJ2K9H2IArD6lwb6Vo1bna+HYzBczV2WGoAkVjeoRdBp12Zb7DP
0Xp7o7spij+RMoLIRBACDHFHe2i9XrvxmviV2fL3iwvkb+TAh+wpszjyA49iBDVbvmMjzJaMOPlE
l1Qxz1Hra9eCkA8iKpZKvcO+3KmuAiATLnwncAwd+LaU1tuxS+6vi/RIxBWnmp0E3la1K1vHhdWG
ueY/eeDGUadV7Lc1I81ftRZs13EZZaJZKe7qkitTCwJi1pd+TgRbn/HaXY69RmqngBO3IPz8OF7g
rxzQDvlpnt5AjJk4zHqr1yL+k1MdWFtmmNEHqvtcfLO2mWtNILCADVEaFEqT3R82uvrmQyyjUkEz
59Zh0S1OuaUKIUVJ7t6cjHT43fGihZC/hUIxHz+sBLxBLDvpHvz/B06SBJbe6xORhvkHLs7syJrx
lzyq+hG2tCNyKDianm7UUWYH3a9rgNxTyJ1fn4lGLOuYmGoMC3KlBBa8kS7J+VIzWI48HG6Ezaeo
BNrEGj3LWSvkWAIhA0edeh+ry5SGHhmBwTC8NOA3V+qXtFQ6sotkOqWKt6PnsL82sdmZIvcAIQdb
FpymfgkpSr855rkwnTEp7R3jMapSHdoKDYAtZ1SpkVe3wuEfgodeqRgaz0h6mBw0Fc/TKDxjWOq4
Pb7S/dI79OTcWeJ4kbLUZmxHVGUNWVFpMc+IX1szyxvM1TVY9ZsVHMonmZq6WmsdvyLJX1lbSFl8
/o9XrsqFZIE3XEknKBvgAdivQTP7pT1EnrYkub4e9KhFNvk/7uHDxzu6Ufx0DDPBsogvSpBdr/ZR
Qm0x4kdNjTfknk8xZm1NYARpteyb6beQaEIlFOnWYVbZjL97oGugHI8KWP3Kum+hG+lLxvRurSkz
S1wVqtuu6O4LKL6DHjk8GChR2yrEk8w0qGfiK0CHZZZ8DNPzfBbdqCOHoH0r8cAOk+o352Zx38Pb
UFKfBPXiaxKHgfjlHm6s21HcJnfyWKRRIyygCQot0Sn13LC0tvTFtRtkd5apd1uSoAf3lqMrH4Tq
p1eADbYsWYGphVsMoLt+RI3GTDtXW03s66fACa1LCA2HXY9SfH8oN5xU6CmiHUWQpc0eHf0pqtqS
75kygngDgGpgCsDEQEreVWAzRe8nN4sX/h+FLAIGbEIIZxa7GcTEBQQtu+XDcY85/YZ4qKxnJF6W
bIvTbtPyGrffZYMPM3PEYtwAgC6V+x4L3ppuVrDP/2HBeoK6vc+q+uK2e/06vdm0Kw4M6tUUBT3B
kcJVhmcO52O9KSkAv3l0ShFScTbrcHx5dhOHXNU6LnrHzuqmke4LiQA8MWKqxdjPqrEElnjQffIW
mjfPQ21U3u5XwhdJpZIMKdzpNlDRmHQMtpXKCw2ap3cAtxt9gzMJGrg5P5t7dI4eVA3USydOLbD6
JbSkg6gT3KW77hMJuUM+5qYbJzJC8EFnM0DvfboHQRtKioFCnJx4x58yrNfEpuqER0cIZK0YAonf
hpl4CsImStZjkQJksXOapMDLV+Xs1sIxEFZqOMtK5OU0nT47D3/QZdL6H1JPMd+mYaRaIh524K06
Zx4U0yJ+EY7dZaSY0owe687ZKPUzr+RCTnC4dsp2asxiejcSibqzJwd+ikMfs/J6Qa3KPrFk4OFL
nfAtU3AN405TFR0fVLRpDVs3QqvXrpATX3cnfw4JYO3KWqiNFfYRbGQHcay3BpL7AqOMnYl04P3b
Msy/QVj6VVl3xzmx5Bm3b+yCHvcJVanazK4Xyxj536Jpf+nfGuyAHRHEhwprVnUz42iI7cvVPjj/
XviXRPKnw8UOdmoQiBg076nOtQ8btml7gJtj0U/KhBz4WFTtxNSXimg4aQWmvDwv6/NfvM4meZ4H
71N0GDeyGO3mNtYZriepUjnYjGDpncIe5hRT/a7CxwSH4XzDPzNXgru5nzwVslLvhod9B2QEFTL/
BZKbGpeJvihRNvLedIWKnkjF6VvvGI/9tpXKi0WqebN75ydHCbGcsFxQeKe93uouR9rYFMWP/WoF
l4G8cnlQDOG2RzI7VcUkF10U/aoKEw9OiWphGH/yFBkveF3HqYCQtn4Pdf5JEWWfzgfPX9YHl7Py
9MtWsnSQLF5cNquLV+88hvq+QXsZRHCQeIcEDG0aQjGGfgB/v5FOZo6nIv24WGlCRTOs0MpHH1OR
ldVwYcmCtmRg3Eo7kuX2+eHs5lj/xj46rcx3L526q33L7fRpDgxLqv4ri0UWVAZjhqvMAqvx6coL
BXIauBtW7O2TziktukCDM7NAKqNfy2m3cdnQA0iN48LL4yxLA+5nNYmVjnfhYxMBC5Gdlye0W6q7
gpIZq02WcHZuajoDGGYAlcgEImx5V6QbKTJO+hZcLGii6wtCyvmsyZrW2AZveAeZD+cAgI+pOWES
ozQlvAZtptw1DXpo7/Q9au/Apd/SOqfAqMVAp9Hd3K3mx/8qNvLd07SRMPasRkEsC8L2m59AIog8
FLGbLWQds0bxgd+INYqh+4C2NFPrzZdaq3lggaJ302hZLIhSDbMcsAI4omPexL4953o9KjF19eoU
3x9HFUysSFvrlgv+F4JvRYQxuERBSAkurd1KywhUrndmWInCH0/YtiXyz/+noEXCUmZFwNyfAcWm
0PPEi3tbf4tgW4/vlkwcHeSuRvaljwnl/oGCZHLjcr2FfQ2unMX74FBvpyWKl6ZgViAeIl3jL8hz
af6OP07zdp+bkKN4WtQYZP8qrwyNshBhMCPRmSxzuBOODiN1EbRnkPau68sFvDZ7h2Mzp/0UjR90
i13yHwdx/dAJkyfOsP1/iFrJvEm1YX38fU7UvN7clDrwBDuFxnWezFIPhnrxicV39u3KNFaR/Kv+
pYPLhQDSa6lnnKZwXJ8TT1LeK2X3mwmQ2Hd4kv57Eijf4gEQ8jMm/IB+zw7VkS2fx7yzqzRC+O9a
6LJz3aPlY84jbqXz14ZfOByUMN788FBKm/oe7uMEoRPXbDyCgB9tZ1HPGQSVvVyWMVfOPD7kQIgn
DtajkJc7QzHfZQvsdJ+B0YNKmIBO4KIY6tG7xHoqZ/zmzZDK/5Unnf96gWSc5lUd2l3Mu3Z/sph7
knhjq8CugNlvbN3BuC0bg0/NdOOf4GCBQjM/YC8hf77ma5/tQBgStA76Lx+k2QEcHoiK64Brg5mb
BRSJ0pHNFV/P4XgWjQAWOXpXkWK7VsEfngpWWJQXe3vYHhpOQ8dUWZSWyd1WdH6mGBX4pbwwSXSF
YCNrZiRV3DLJQqmAqG/J4x0DRuUcS/N5HuFbI3lfEXp7CLNB3P2WCCcaGIE1ySDjpa5LKXYkBapm
+Src9ZHmPBDX4T0opdjlTaZBn6YSl90pvUaAD8OPhrcbvz5GkVY66XnoGZ3ub6DW9o1q7uAN3xql
vVWF8zSeeX1e5SKWJ8fEzFLObmzP8Io6fDC4sLnjE+XCKJyuuU7P90tzO0amV2xF1B2FEP/eZ43Y
7the4MVdQ4Qy6gPG+AGG6L89qlY4/Yqn3NJU7Xul5JkOwtg987J6g6voA8BmqueIw0LpyP3eNZAJ
HfnTz/mIG7cF67TLyWmdyi1xoBJetQNkQOTWJ1NSVaHw+Ph3BRVPKyRhs5YIu+StDtMirUWF7EqO
N1n9w3dP7IDVclDtS7IKh24D/Ax5aO3ndeQ7hXcjdGa619shtZye18FKQ0TkQztmwUBEnv29lLSZ
E1ttiBrBK3bRPGSezmazoEQ/59o8PJ6Am3FDHjyOYviOsuhNi7FzYuFZ3AnygmEI/9INM2yGC31h
FJtoBXh+TVvec4E4RoAcOtH203BFOTHrVIQbJuML9Sc2pSJgCEp5uwQjfg+z98IKyuntPjNHRTWL
52gRJRzYsITHVQw+0AiIu3fCuisp/snYOIXHginQk2Vig+u+dvApIPQLIC/kRHRlIWTl0ee2vg0C
b4JbAKP9jfacob+3/UxdhHd5/Xdt8+D6zikiSnqB7JhyP6swMx/lHpppbPBHNiBqagLNo78e9PLh
t2brc1F70orLIgmFnY9oV3nJfnlICsgbCsyfo9nPRAEyNCj1XY0fylR4/pMsyQPAUn6wF1SjJl9L
BWGskzBmShUxLYDB6Hztl/Jwt4a/XBUSqI/ON2BAIYU+h/4CGlOSlioz7Y2g3uRyA1qrQMbd6Mrm
XKJsu2ZP+/ZYS6IctmrFRpQYScPVeHkMqW0ceyEeLMw/kAMnULujA8ov6S1iXA681s6mkARq5goo
NKIwHSAypZ/LnxjlTZlgerZ9lSQ/dP3MUNN1uYxI2XK3lPycgPmvX80mW/4KX79pDwmwCju4Dn66
3QnLFpVryWvUaVumoDRI7d3594nur3lqogN3xhX83FnW9iB907amvAfE56PFtjPJkImjccmOe5mI
23yOpfxGKQgFHacgrwsWVPV0GkpQMN9zIsuNsY9w1Wctc6MvUj4X3oNEl5JVGKamVcaQXk85xMm+
P/tmSIBJhUH9BIIT5ZVPSstwMtUxxJgrRPNKwgvpQU8dRfQcZ8zQJTj7Rd1btUw/Ynfc+aX6NCGq
T5aV9P6E02bgpie+XPjqvA5hjbd1+MJNzTaFuPpbZwnQPHM3IxPtUCSiUZs1nFjMu+RjjCTZlKy/
Co3ItMYJnT48YE336l7X1pZoXHVoRoF5W4p90hHUK1jZyoVnVLytT6/8aqyKprSWqPaJJbv3WfSD
P7DWZnUfOVuoGoHdDnv77xVnw23p8QL4V0SfkobT7pEbZsG3zJl8U/Tttuv7jU+NLUxbHyCY7rw7
pfWZAbdwz+casEaiasodYqy7X0C80vKHbqK15tUHjcFiLWeuBGvNAhAkhWwYS5z55+d/AbbF3hEN
5XGwVxhqMeuddI3TwVy3+ORgzVDIVEbCDV7cKk4ERZesu32psa2UrXpyPwnZkQj3g2Dz2Dn4CWqj
bIwXVtjTbehOyNKM6BtFjSlMfDjB6+i21SOGLfv6TeiDUA4F5FUv93+Tm2Tk6PvO3ugDKhpIz1qI
8vgCrSpqZw+3pK6gQwFpo9biNgyYtWdKn2Da5T7ZjrlSYwu5ffRZHamnVqEEbJo1Ku2lBwpSdbML
m6G0GCMW4u89QKQYOdP5VyeCMuZyyEurLyna8HlXDJxMTXzh+N8FAqB2y/R9XvI1BZaynRJ/z4GZ
PssApNTh3RRemdB3Qy4+H4koMQmm9l48kG1cjGmb2dEVWZCKDhEdo17dEkuEiAmTn9nAPsuiTYL6
UrkSDPr7wcGj2Cx2d9FmDqn1sOslHBe9oY/PTdDB/4z+S4fXEsPFuBLqJl5KaRk83YadSvPylv02
xH7QPSiLpGJpOwFCkyxXnIuWyiQhOeRuBVO3UQ904LBEKjnY7H90pZ1o8aORbn7qC3NxJvtvEMUA
1b2XW7A+aUBZkmtF7hHmPBFsYDSpaP+NP1f3HAd3mx1cqRTXXCfarLC77uURBZHhDospgwzbPAHx
IqgknzFVQSw8z9EAAzJWcLSEOQ0NMdtvF9pDgu3rrbc+ffdosc6OaRn3TagV7Kso/Q4uOvl93NUO
PcKJxe9+HeJ+qNMNHI6scaJym7jeHcdVDALV1GyRXngz5hXp/zyEkBa+p9QJ14rIfdsufE+SLnWi
BucXuAk24vYnMZ5NkOPPyKNegbchKVKd5fbnfWncOmfeiiHtbmzY/8w76nLWoYM3gZErFXeF2JAy
OQCF9cjza5uQynLXyegp1uNdnjoauRUXw4q96xe0QaZy6JG7+zwyswqQmE1UBv7pTKa9nnQC851h
pzJ3eMILdXDEpLvTBR/vODceLCxF+KKx9tt/Ove74+MJwYgU19r80gX2hVmbB81KAorV32gPCBvA
FrKJrsNx7859KHfDELzMLTA/3sgNRnHX0dsy8w8OHH69MYiAFLMOuHHwsGavI8H5DdsLTCMl962G
JT7htRqU0UW3YcNJmnAEUQrbQopoBQVMiL1fb1ivZEE1235uiLslpy5MvDaE2UU38Rkc/HO3W7zB
DS5ba6Vs1t73joeMah8L5hUR4sVxMYrngvrTAfL6G1PO9uwP4P1CJ2sM4wOt89hQBRPE0fdV18v2
3Qu7EkSXezorYI2qmetPTzrxhEliJfLmFRe2uGuatrvx661h/E19fpZqGsLhLJNbz4Whb6ff0aaS
bTF4ep8vS4f3HTc0BEcwyVNeDErsHY8jp5Z9U/f8edEHen7NCVQ6g3He3Kdqmv4zTz184QrPgi6j
U/VGCo/xqfE5XdyoUbXgAd3kJe3hWw1QJCpwJUPwGos6byWh9bQLTIXlZU+wnAvBorZahBcDrdCi
0aVP2TRjhpEuCvqzUWogdTzpTmNO47cbwvXwdvhzO2GMPGBPkZCBj8H9pTjrxEO4w8VkzWXgR1RI
QOY4UrR/AhC+xzXTsZlmIao4OESu5j8sEUm+7it6CWcovIpX2VKCAaAYA4kB9ojvnw8UkTHeKABG
Gm8Yd4UG6N+TseMXiZDflq61Mtg03yZuTmPKpCRCYEmn5ymyVvK7/0dWE4YhPRT1vGZFwbcbJMAD
18g1FFa2aG6J3N/LOBtBNULKZMjNCrjvk0ECh0MBKBKAj+E+Q57RKAlCpE8WazB+pGV5C+3xEth7
TTjs4sLixWzhNwq6Utt66PBnrL9jnltHY0GqSynKTNbxrv/PN+Y95CuNwWJhD+JD3K9vq/eY+5UI
EhPb8zKPtLulf7Jf5LRR1jQRQOYEKtMTl2DdQf3O76w0iNVrYMMh4whby4+Pgc1ARMBZzY/Mx+/5
/hXXcjd8dhzwNUUvxYnz+kXbxUjR3Yq108redkpg2zZwnnd4wJQjblG+wsqKcjCvPxkyO2xV1Xvo
8IBJwwzwa2IzJk883fbmfc0HcGiRMP9oyFf2EmwIlnTY5XegcBxKFgm3kDQxL8V4sUs/ceCFLYzN
OZgohdgBqHol6dWNsemmLsBPpQOktD6eD5WY+zl5XshRuAIFld4MXqi+QfCtnHhagfLVrqpjsEmA
BKJ+QuZf/F7kGNgIacIKBDq3DJM98B6RJC6XYOYqY6WdP960a4h4gQOYe0tti6p3smKquPoIerrT
vXkNDbnwK6wclM/NWzofgx4ZJt+ax7GQkJyvy6dGh5z981FQbZODRQaZFrTHwfPGzzZ8LVFOo1nw
PXsM5Slx2eg5VvYZFICFI/DrUlY9cM6BMHXGW04o7SNd6J2lfg+B+o9v81o+5ZyeKySWBo1le7nN
D2+/SFCcUpKWk2mHSCZf24FC4C4yfqpPzk2icxOqkv8J3WKBUIyIJ1oUqyBrqamzSKhde0mAeoNX
QdTy5j9dSkBlHKnIlGG26j3iOYxjIKtF24yQNPAlmAqVPAM/kXTqFSXsP5484nhMDQgJHRgad6YX
lMYKJwLksX/9NNv5TbYhYC4ZMkw0o2OhD/Z0An1NtitqsCt+LmrsuaVHQ1OuNq5n90cfVrAe2Jqg
H3wydFr/e2AyETA3qOa429AqxILY1oS9szO8wbarkDw+LRT8EvnZ1INmRAjTTpSUGwVqkSudxpFb
KrcjIb3XhEdvtMmHqIB3KrBPCsCzIZtyEc7hpoqlTmB1EjjzxtUqtRXm+cf/k0vS57RI8NouWXd0
1SDUs1uTUjx/O4OMdIFt5ZqlZrenKJZtc4r23zwP8npuow/+EtLGRo5ImbVwvYRrkOBDm8LTRLqb
SMt955t9I+bI4IGooI+YF9WngOXWUEE8+ocyMev3BlVY0w5SLmIyFkwuhPGhDzM4A7aNWJDVICgi
LfibetClbgWIvVK37o2bi9gRKUrM94kHfH/gAyUpEshWSnLZNJu/8KsFb/mvO3opKEvDCiTk+WP2
kYyRV/hP2/cgZ+EB50x/nYDmsEhTDTshkWWjISVX0SH5QB2lgzA9jtbpnu6kT9QA1UNomg9BNIc5
KD2ntts/LtDEzveqkwQhIVa0FNynVBXQ4pgLk9dfjub9TzFAwdgZtREq4acftX45b0T1xT2EYAx0
jGBSfDsqOKfv7yeIAjMkSxyQhwWimx8TgwEfalyyip8+ka+wQrnR+pIPtf5C33NHmaa9nMZWWL5Z
VkhEgx9PKcK1tsqsSGL8pH3PO3jMJfB1FwLs55vr97BJ65xldXrSeq6sTbO6KRO0coEqPIcp5QUU
8yboIsk6QhBRsbdvUrnKAFUqyOSTxCz/nUAKF5mQm2icZRHqGSpnxt07uyqP+O//iJ5T08Q6yC+z
r+CCSawP4TYvPXbeG/UmGg7oHRNYBsWjeNA535/obKTAXDG+V2lAGbvhGA1JmoqOqbS28fCR35Kt
Y6ilG2+UnWSgR5WAEWdkwCCHpt04bDVEMzOoH4F0j497fTQrYwbM4y/OwKAAAGd2oufe/DxYNiRA
p8dDPDTXW/+wDzuPd6FGqo3yOeU6F3eBLc48Whwc4I5ZEhVg0zUOBKu7ZxxcmEJJ8cLJ0ZtSUQTL
V1JwZBj2atILQD74C3zJUITsKSflWCO/BHuy4VcItW/ysneGTd3jcyqFU4Hd7y77Asph1H8HLzgi
pJRckd0yEeodVwxyLJjIORGVAvjjCyt0ZGUDzaPuU8QxT3yCA9lVRsdg7qFtkoXHhOO8fTricBsh
+autHQ/4/sPdm6jwVGKa9M3tmycJS+gsgrERbMAwP0+ELZ+UdZYmEB9UMHKV8UbfDsFhjFHzqaIM
p5thFgJxEgu4LA5y8Ou9KU6QB+++uSleqVyCw/qZYwxRGujyErTX+KzB/1eFRskJW3ANFhV+SYEa
3FOP/2BN1Wjj9O+3IGZTwBroQwPsjRjjDuTdtG45eiU+l+o+MTRpBxbXsP3Lc5hvHfHqqu/Iv78s
LU20XG6jrsRNl/7h3pQC/huIz+8GLPRFqvKrThKs0+7t307TIj1IPur/qzKFqGpAQbxK4CoY45PS
pOC1N6+zqRPwinhCz9H01vsWCZu2qJjWXONO3JHbT7hDYNgbiDdPdOBcVhVmPO+cer3BDX01uOUS
sfiE+XXRMpVMpi4oGq5PNXD4byZz59j9s9TJZrJWoxpJdIJA+pRdd0s6hylONWUcxrd5lf6dzOCd
WbXlZLUjl9m2vxBFEH2lpj37XleAyREoTzphzhuJwkZMAhbsiqGQJ040AojnUy3VF1RhZg3oMljY
wkxc7dmmy4E1ZSiZ+IqopfSpvf0en3j2XXtBK82vnU29v1zBsJ4ZRYiWZ7mPlAz9jWszj1Oz1VS0
aCTv+0jeWwFBvY0IeMpDKULM4RBjKWKot16HkS33szmgS/8SByduaSYJKRjXaSPOTUfxANAJPmmk
AHAaokEmoURS+zoyeQAJ2xABi/+c1M9Ye+1Wlk2VJiGg8GcN2v12ktb0lOv9CmR2olf62E7/GzVR
Mz1f8uEwleoeShAXPWGLUFTl8gMyT7Udhi8XwfrZrhSFiHHKXbS9EeggdefmV2hgbwGx7Df5JCoa
hJNdG+JC8CmdQq2AooCPrBXyVyPvAZ4PjHXXNCseTw6NaB509GHub+/JWIuY4l6L8fUnYywBhUT9
h6N49nxxkA6ZBJAdavV2zbw7CYLDLAMw+rr2onp1i6/hM0S66+LU/ehLV8kgkrDeIUDoGHn2mmpF
pq2TE0sU/j2Rk6c4shMO2+nmfD7aQM1uaZiITc2NNRs2JWhy1BeVZzce8eRwLhQp2zCfYKEqrPT2
EhhIMtZ0Qh2V8XbNY+fi05Lm/P1LagXLY5iwiz5jHS4fYvfu9bNrIgeNx9+mcc4rvDQJc5eOSsWy
b9F0IRdpvMr7vSr+49NZpM84Rfo1Oi+G2iMJ+/TrgKTzkf7mGfFzMfGF2Md5wzCZPEQCHw/kX5IL
YzGVypKsXsNy5fsj8Rc9p5/RXVPzvBqMPcNR1JlADxdlpyTihN2yiXi3Vb6JlntN+49equTvnVCb
SIxNzQ1oEzchSKFyq2mjORx3NEX978Ceesw30yC2+ytZm9A0wby/wWDJb9sdTOy+VuORkrrCTewm
skZ/Faw0MtPLZfoqH6RsOp0TYErhakOZ2NjSCISS/PIK9zHZEfKsQntJtBXTCVJZjLTGOjm2by/A
qCpgGhKhm9rW7wL/KOswmrORRYtMIVizGTBt09jnl5S2rEcPEsoSMIhD2QlUJxBMG2MkW9FjA9Di
Hdg5JItkFPQalchgCnim1hDDuQpPLR2+V20CgsQRjMcXr0RNW9mtRRQBTg0OSv782mpE+uJi56zw
6gc/nF/XnWFO7o6BjTS/kWIhozBTs3nzXiNRPhll/bgqAJktBjrrmWBuPYdp105FHbz6bAvnCS0L
zS40EcVbr1Ii6JlmL6/E6rBF2kVh+9TY2nuD5inMOuUbkYDQe5FPzC9le1MPAnNfXhGx97up93TL
bPiejy/zcJafYXVJi1tfTqbq04R/Ovbhu6r6qovp71qH47huxJsw32ZMCqCuANqJzIx+MN80ZHBq
I+pvrOI41eZOLI8gfcQrQkFaLehORG0ZKvbjvQy96iZauJ7joa8VdTuPjDLJwp1gEb+df8SNjonp
61OVjhfmS6fPOIERqqyR4FicPzKWnRUBxDcjrTLLQtpoaO7wGUo4Ps44xa3Ad6YdniULO9bjUOMZ
7Up57s9mxQar/jFbL51F6dLK9xFr4xFTHRmJCQvAoeoy/tvoyB6gmNo9MdY3n3AsbFuoNvhCfX2a
GGuCwWmnNe0O7MnQBWHAj72oAQYLFlu8MJOHB2RjXTdSebSExuNV8YFMZhARbxI1ygIWbpTwDON5
sinxU3ml1gAvkUqmSV4IYtBG+Asm5PpKX02Lp4YZv9mi/t6e3dalJUAyZuRbyZHKj0PuJaXPozdW
JT5u8V4ogtqOrYHTXrngBmgyy7ZmxvamoEPjpAEC7yPYEzOvLGTPLR1ox/EXTOM3P0QyEgeN1mYk
ePFBlVyWHdjPFycn7LY95H8PeNhDkS31I6d0jwafE5jrjeApBQktGY0tGtDhyPpVBRG7mbZowNvz
aoCISbm4uEBzKkvUOwHAJv349ZRVgcTDz7R/YG9Z/zMlFOWDlrsFbWvEJ9tuNA3GPV8MIlXUw6cA
FD8g1uCgl5YPs2WUibOf6pTvud8bDMJN2QWM0AIq4Pp6WxKpJ2Fb9o+71fmfMnj7+4sYZnsLKFSz
AoCCJZ+c3ixIXEQnVkJBtpx6xjiDYfSib6PAL0Yyx9blhefTbSfYJrUqw4xFoZTrQqbmZWi9rWgk
Sxo7IBYbHf5OBMm9YnQuWQoRhFC81oGqwnfOQMGP4mm1NlYFoAnaaLFXrDBPwi8qQun/NbcEU5Dj
cTgyBLLRDqDkPVikf79p6bwlrm1EVWtdZKpl1867N18TyWbtyU4Um86CgBVLcAqaatRd5VDRCjEf
/u2zQxrp4J7d5awwDxe/Il3FTyhco1NR5DPKf1NCaPneuKml/j0vAHetSMaHyRErdiv1pVGmIyCe
i5LyQmH7JfJHcF+OkW/h0iluhZ+46TJk77C3OUfLizeC5wzl1B9iPGPIhjx+8G2tA3uwxR1z60TZ
zOocNPZNM7tgbuFV0CiqQpe0nIFoJ7wv6pqWW//cx7lbKHoB/PUG9czLu0lQyooaHMVhTCQlk522
rqZXK5tA82jzIMSegR9G17Lk4er7tQiZ1ly65LHFrMIwxaAb2XDVy3eDTKLX/AezEgBtu0WwAG1d
FzDWZ+PPsaCtqzGy1Di3tq59JslSWcBunydgXyVyiIvcFv5uVR+vCr+F5fsyWKKZB7Y7v4FBp2c7
AeH5h+jVj9Iy20hcKqfYGcTt2j6pTPNp3x8+366VUtepFgEb8NAtnVh1muADXOso5to/Ud8VYANe
cQT+A6rdlEq0rlkX5KMSnU3nUaiCtX9bhbe+xwed9ca+DWBeVjL8hrVDZNkW7Rk/90ZcZJzzbLpZ
xumjOQKdsuvh1OLqfIyLCsKc+wpOVqTN/T/iQTnmuun4I1bly2mcJzYIzqsk3IxkZQc8wMWN0t/a
qBVvhhenScR6IXeqcd7nqbT3978TbzdKd6Uwx7pYpn9AaQGrao05rQvGSpYpc3wEk0Z3CotysI3j
5Tv7mdCuYXFOtx8HGVA0FpyPs0nury0U4gQ+eQGo3VKsjHauXwk+Cg6o0aIFcL9noYchMdcxsLOS
UEiGRToBgJg1a92mQjOrxB8irMvMHgPRMUGxf79uVc9/MAod05icUkaeEcGjf0qSG7cvOubW/Wys
dXKF4bIT6rRfo/Gnwu3Ef4EwEFhqSXr8XyhhXPalaO27L9JO1tsg2cdc8GACr9JqBR5IgvFw6Ads
nimjRpl8z9Cv+YjzLghA0pOfYMRi8EM+Qn+7MkHa3TLYXP9eI9tLPDgnelFd7lzy0mDxCzBP7D48
5O/DqThGFn+427ctU5l4B02pmBA1Wqjm9qqKDMUjAa/qLGS91+dXeEq6V6Fsf+bEdjJqVZQ4a5af
bkyOqtdGbLfO/ZwqILAGx+MG/rAR8RzlZZ699cj0iDKdQL9olq047TtqnSHzmzCxI7EZ+BVEnESH
51JkARlD7KYTbPXbtCIVanjmqL7TgT7Ff6LNK31/cGm0K0hXnU6hi5V82IIl+BjW5wDOsMiKVIs0
/tEDCemYYS1T4VzCrro3Tsf4GqiB/JLqeD4+LX7Y2dc/Z40L/mc1WiNE5+6l4aUwI2IpHhlD4Jy1
W6FhulbFmzt/454TQtXhtZ5dsPUEi2eyQuXEZp/aUO+QEF60i2qK0QrA0ex7cNPyYKM2iyt6kY/F
Y2YczQw803zvBQs4c2Yn4wHkvGUd9u8zwb/N240lP2DovQidYTGa9Edy4658SaC7Hg7Z4rjgOds4
azlvGV2gpaadn/TDCcsJJ0N24FkfcD97wuzihW2++JVh19WCuGXfZWOTxMXuvf3rMxtXFaSFpSs2
dKBFYPs6gLcbliFn4c7u085krqxPAIlDlK+RFlQ+cc5oXBbxyH7pcWRTi5tV+v01MKkj9pZQ/I7L
ZbqyUnoCJarxh97HYNjpuHVgaL/BsgzbFQGQ0OS+SjlKaLFUDW//Hc9GKzr5oeCoHw1xTmSJvkjl
IYOXMyi1tU/HK2ge+KAx4lJ/IOqTszz+P6/DN+GLs8OhEUs9GVn1V2iq9J5YoDsMbwHXH7JwQZAz
qHfFtM1NnLZBakKAjpMd2P2aqZhH/+VKtGaoydYoo1jskvwjskba6UjYO73JIBbrEdmVVSdgRuER
pxSdXDgHjMNg0/U0hdu3Y/SNKNzw3XSHcoGyVdgkeZwUfzUisd0O363CWi1M+hlJByB+43H54B/V
WUWOI0Pw6EmIhOTImbrsj5qQ7Mzt2YkhJKK9qcHwYLGk69VAktKB5agcyRqFHDLmEtoMpvKEwHRk
2163qB1zdzQaamPMDQjhb3ZWvFgskPz0SZ5B/G5rx2lJTMjRBzIyzQKxnuYNehhcVYysUiAvamtR
Bh5X7gnwO/GZ87tVCwXs1PBKeMEIxBBD/WoiKcyZKR82zTNktwbXEQT0/WkoI6i7Bfsbc+XxT11M
CEYbiLE++svQjTqlfP1NBbY1TNgVMS3E9vtAaU9sDvHt3Fmm62dukeVDW2dodIKVEFzZAkRL50E9
fmYV0dgCt++HYxMJqDoeZbP/6umMcyPsq73gAC8JQEH16kIgfL+qygaK5nnXLP9fmj3+F2GAZxvg
tl8IU8Ea4JC81VjJFiGNHCItCUg+Yrc/FLyyvEeYcowb0XVlFuYLk72WMerQy2JT8rxONMsOJga4
lloZRtODmGm/t+tKziGY1Y0Ee7yug8bkHmrdsq6K9ro1yTgv3xeG2ImqMliAb0MUCpVorYmdbluU
amDwVy0GgGc8wWikqlERVWe26okGL0tc4N+dDxR6JBz6o9OwAmpQVPKIzrvPyXuKsLuiZj2QqL4d
c8goti85VeXGNM3TgPX+udNDWmJZ4JbUw913epq4eZjQ00+JgY6ia3OEqrxOqYNiRP4mmbywhZTT
y9twEp7qkuwGCKb+O0qy0xccRcRGwVW1s7Q/1xbP8jC48ju/74Tz4welMFLDUeAaJhUg+EP7Ddo4
U5MbML4FiXH7YFYuWYniLnsXf9o6GAdMrHcoX6Z/IUaeyGzFBpPMktSCm1XzWzUx9+aaiRwoqwUy
72CVJAZcO1etIYMNRyh/ME2O8EKq3YOdhDciDRrYbUJtY8DHXSxr1ivRS6aG+1METGNPChMRDusL
khUf3QNixlQknFYAdEjJQOMU67/Zf6BiHauosyyVJFfiUwaKfsIlcg3+sJrlfjnu+Zg2xZfnfvpi
txmBd0DkyjkQ38IjcTvelwkfd/wP38kHeHorxStlkYAoL7oe/YwLOGdbxFbtxtj6UEgUcWtrY7+C
rFeKor/co7PQk6KTC9DgtpdP9okWNEPcG6U5zTsFNwu5LH+HXJkxckHreYLrpclNMLJwq4s5uqq3
tzAUnpwg6rBCujb19783e9bbuiXu9ckHYiIVE+0X6EkCzmUJ5OI3aXjmC8JM/xvsHxMAf7O0WHcW
NzYsyPuxU05q2O9VZnDvi1/3HyFejOWX0SWUaJtRiSdGfyR8MnWH+hUsWRc1gqS6MNV6rDuwoVo3
+cGiKMYO01hnyhF9zoy8GpIeiFUY++Cvy/OlPLtnbQXDk6GTsnw4QBNTVaoKXsWW5V8hZ9Q2eTCe
1oRl2Or4YTtL7ooDTNI4/9UvqZgNZfm3HA4+Ioq8PYCpOEEzlTYyEP/ePiz+t8ar1D3uQduB7Xsr
kuH9OPYwMRNoxTm65uJY1aXIjj8tNgmyoDEXm7xYObtlnlE1ikiv0LZ7XFD53WlCRqdH84AZWURn
IQKnScX5G/HsRNDFDcVoaRsgq8pCPOypWuW8xneUSzLvz7h3NIJN8HTwzUlDOd/mBrUNBsK0V7au
BJb/wR1ST0Wve73+p7byP5/VtaSbpdnqDimBJYYgNYYACm1PXlnNP28oKAGuF+X6arQORqaENquv
m0YJRdYujNqHqO/TRp/im/NzxyW+/G0k10fP8wbupXDz/vp+1D7I/a4vsEx3V7N4dHyynibILGGe
sgn6plYD44qbmlmUE9GXV3cMVn3f/d2+AaukGEQLkzRfe6NQp/s8Vo91K4awcdicosv4MjOEOuHW
l4iQZMWghCNEffDq46T1wGLHMCsKfcQIL5geeWbSVMswRNV7dqK2Ik3gSFzaLdeo4FEWnPlbBNFI
Hb9lTvBHCkAQdSaFGOVDl1PR7/AvDkrmj3ta4L/jow+PH3LY3H8PHDwiEVyOAMIERQhaDSeNN31L
bP4L1KqIIyjh1wkNFBjvqSfydaqcN+4OKkPie3DjSYUWScqAnGwyt66vn7zfHlq40Wuy6xolNdRO
fDq5Xo/aW9Iz3Mtk5QTxZFHiAlyAMlFlW0lMwXEYYgbPiMlU6WmmTqu/2Q1iN9iWiDUexHeZA2D8
X+ax9M/dBWUbLwG2d0jyQC2yLOV361x7hAkKkqfA1PikNN+ZWCiKaRu41+bI5uLPXqt1ZAB/yRTv
O4DvY0ovVP/DZDmBn3evLY15NczwhdCTEYr4AmVDyJvIhLBN1jBPk7MqrmG0DXBFwGSAn5RKKwfo
zulRXg4BpDE/rRNqBq32Ch5mTE+hICr7P1OxXZnD1dkoZpxSjD72AYBTTxCwofIbp9S7Vmq6b+zm
yjHYM4RrcTmme/eYQJj7jNfFnhAuVqd1l6S/zI9PTHOrvFDXhX3mKdTHek+fy//SUYvLasFLUCt3
3VbDqVIgTgGMrjccpNMolqrg+WJWOvs8XzBX8eZnWTBgoQHtri5pUOsAnG7Rf3yYIl/PbGrvVgot
g5fkF3Xckp0zU2P5qohY/KEXnetdeRHsyM3lo3KP1es5cQdKQfKLJDxlH2BS6Jkde33A32GjoQWI
ou9avGaW7f9G9ZnWphfsrh5i55kVzlsNfznOElfJYeCIDrYv75vBXc5KT7+/0GOj1uJdeX6ol9FY
GounqJGWlahZ9CWAS5sQiAuZU7xydlOeNiT44XaEpH6XtvIKtNcn/FsNGEILjhjvzYR0GlmTcx2R
t64IZycXHh6JcsinrIdLvITMYyoJropYJVX20gKFkKTEAfG7OAPeWxwCxKl8QZYYd9MG9AcIhc6m
irszsZ02xWMN03/XkPMA1TQfJLSM3wM7B7yc4StBVgsKSuvI98+1+XdF8GjfPPXyw7eZys1eNEQt
g6XP1dQqqVzFlNclpxhS2gjnQVetiFF+TlLR+3WmCZHkg3G/UNhmCOtFiBn168138jSJu4p1OzbJ
890nZvI8nEq0CwlEZXCi9g1SqGacWFYdAq7zEj+u+2Kgr/BPEniQm2avpRlcKQJkId6SxaPQnPLu
GCVo+SHKcBRRGG92MQPJ7wycGdyIiXNGyWS5uW9cGZq3N4XHCyTAoeiZsKhxEa6CR0jzieZkKbg5
7QmeZbg7nAKK7wKUVp2Xt3epHPRSedy/H2iafLoJCMCNlmrwKSXDE/uf1kmmEIjzHCc4gtkX/CNZ
k0XNt4hxHA+BGSo6eSDc5JO97n2MAEMr1LrduHQ0Kpn6JOqaEi4xcrUHrCnatZHAF9GChKlpXiBe
CuVNWLOT/kZ7k/wCTB845BXh1/JLxoWFd43CT22psvKy80jL4icteKg/NlBOaSWN0qDvbZzyGTrc
qrCWG73nl2/GRSSXUCJvAjWGhqTerYKcPFSoSNmqkayX/x7HTW4FqZ6cWel4LrHRgrtfCeE/pYae
gWr4wfWt8tZTt2WgMfaWM7/Dp8xt1tIpkSQ5Mq4OD/R+oNKg/sAcfBuuaFMwH+T6QZ1OprtAfCfV
szO+ETD+OOUnGEZp6ydRB6iMcQNNV0Htrp3fiTaonXh/e66mDoXMK80JOAmn8WSK5CVQOQ7HLU+H
q+oZwErNrPwF/LwYgMZ3k3sQISnN2jUDJtqbN1UfT54Rm2tIWhlPsiIE5uaR61ze7R+szdWtDABj
LqoSM3hnuHOgJ0urtah3N/QZE/caML0VhvUAZhz813n55QErpbxXigWCfu/GlmMcobG4J2w1aYKb
O4mxxmod3aj9JKLVbxsAr4w6ExsuBnEuWeM+4pP6kxyDqZ6DQYOFNUuqxWXT3EgHKVoBwBbp4Azc
Rod7tzhRkDOyYyZQlH2Q/pJddW55GWqNeJh3kHnsLakQ2JCWGvJa3MOpRDDpALmRV9aRosH/htmZ
7p90aWq0mtmY7Y/peXq4R5SLprUWYp9cwUlPOHCnX9rclMkh3fhxhd2p0kvuBCWP912cx2jVYnVV
QU9WQ5FGKKUjogqRh3OprDjlgWu3plYv9xgyB8yzkJwkTfEH1wSoaQtQ41pF3E3Kvb/xKzVekEOj
CekiGfcUeTLXIawWjcf0jDoljhAm9LlxcPcIn/vWfQvdTuTLewhhb3Ye1crW6nk7rxBCeB1PrNa3
E/RIBQMg8zr5L4wu2fPIWI7OB3c5kMK4N11zERbsw+iZvaB+td93EhscTO4W6hrmLoddk2P1H8Q6
hYQcVS9uZvpNZFTHzZ5bwAraE0K6hu1MEljoQS5JcJcjBLHxgS+ex9fGUpzUurq1KL2jsQ9lsZcN
BaBPoYqApb/dYFVA5RbbxJCwYj60JviqGJVdKDv5M2Ri8F8o9n2v9Y4WuWUenL28awQDuCn3oQtK
fMHLOW1RAd+ZGQRe82FHFB37uWp0ua3K/FEZ+uGXJ0qJuAu1mcXzmp+l4SRJ7n+WtuTJ+yj1FuTy
rJXv4wC2dA0Isd9xzhEqw7HP+CoV4rQhDeQkkE+qpGTySZQQuwetyLcl2h26/zglD0COUGkdDBUD
b9ETPlbA4qlM8iDIlwMQMnUmrjPxiB8bP2lunVxZWkiubFSqVOpmEyMtbF6LfeV2Z9J5TBwiAqKc
kfkVa0iRipSkIq/jHWZwmpSGqyrsIGDtqQHz/0N6vCuaEUqCH5veXWkAUT6Xq3Yg73JYJ6liVjm5
6y5GEbW2mMesWPKND7bdXw2xi/7hDd01a/wP+hfSLmDTlST2o0XVf5qarnXeEkHagKrkPRSnkRx9
Sri4d028CcSwYuDmoKbwt5a/1Bat2rdDMG+uCzd1fSs3aGbTmlUFZxWY4vLy6JhaEMIzaOoXNdqc
HQuHp5PENKRryFD2QvVaH+CkNyYydqtms07AovaXdeiClMQQF3j7urN6kN5nQ9Anvs/xKPOrM1YW
j1a9+af/COFfdLBHW2rrANpPEtvdm+kg3vQHogEsjYuiOCTJT/ewpbErK9XAyiKkai4Lx51yr3fD
hgCHxf5lOIi6mobAI8J8byt45kDHqzBV90NMCsVq3/Yy7avZAp+o2mLTMcHWmuBguE3iU9ruBTcu
oR0wN6pgRg1BRfoZRs7a1UPzgnrgsOYqcheaDcs1R6/xRBYgUHR41BGxRfxYnWxli3cRxCWIsWHJ
PNq4gU7M/wALFi+mOzIRUfI7BymIb6ND/xZWhY48sn6alb8Dt0A9ZiEltqcCJ0ww+MyqWusBfF4x
e4lzrN+etaxz9X4FK2qnweuI/HDEMakOJUHJLQo2g/bYlslTCbuAzfmA3qwSpE1S3y+8HJk05G6w
Qhwn/V53OKVqHT+PUwlcDxX05hw9Oxa5/KPiGmli7Q2B4QfzVM3IpT+91EBJ7s7h4KON3KUFVSgL
AmSaVNV1Gcig4jbaAiGOVsQLgHQCVHt2TgbIG69+T9nFBah1tyIsEDZQIgQRuwvYBrMWDCOeI7es
bqkGLdkZe4td+Z3kJZ+PFmqLEODrTuO0ZFWtYpMJVLyH2BwkPg+Zxzr7bwDXeHvAJKtVUkaJKYkb
M/WhmVtve6esE+yPi1VRJeA/FlEo8vTx0Uec47iueaq8EDabOZoYtN/CzzoBdi1agGCWelnsp71e
zWVimJPkEXaXaDba8E7YejRHec5CR73d6Yab5/z3ZVCp2o5p0nTRoHeDpMOZEucminC+1Ec2vAIz
/QfWdS85AAbSMPZSZB2SFQH0kpo9i6fMEzFn1jOQXVnvmHHE1Ctmo0tHwXG3o+gpgstwcjXnBFEY
AwCUVEQZrYW9sOe8hjfu0q9GaIGdgkTZM8S5byH/tZV83WSbGXhQFrP476DVXIbMjsCBIXDzlKQg
0+s0k8tbaiC5FLPCDKG+PafhWRUEMP0dY5u3M0A52nsyDwzza7o8lQVn4RYGC9pH9Jt4Adaz4mVQ
Y6vtdqt2egKSyWsQ2DsSZBwHDh6FckabiOhVbItYwaNgJG69tWHSJn8pueOFGLYINxDAGxbaCrLR
h/WFDimRh2BsQOSuLDUIhvTsb3N6MEffkgiQCD4l+xpJ/629aTesbCs2LC2lLt4NNWj0bKHcMLVv
IgRfo3jeqxz6vx86SwRrJO7LXF54ENYM2oIrWMydeqdTblUWfzLXhcf6CMj2Ih/Lz1e9sEEueV8n
mesA8wZ5u8TaI+DmCiQe3doniup8gJHvlGEjSHTaOiBIctu1MjPMLs89vGoIQYuBQPEneZLIPyw/
zSNKiV2CXiI4k03nRdSdWIfOYxzobmcqOn9icBuocGL/o4oWFuYTnlluMDmphh4TXq2FM0o4D/g7
QUBRHwO7RjqCZIpOrdenDaPmoNUng66ZrxaRNVfCtYUnoOU8/gv0AsDPnSX8hYfoGcCIHstkA46F
UJkP6I82XVV5hkcipRdy98rHq9FtFuClDe+6fpwxkesfAHCr1La058fnkLOclDECJpDOLH/Pbcka
yxVXS91xIUnyuMGYJXpF0rufQXAcrAQ1FZ8EyqVC4/l5FhPJWpv9J/goEsYjUrGJvBNxJPzC9RVm
oliYLliodVUUE7yk/UPFuXV5YrEXoIgJKr24umUKpFmqtWYAnU5vdyKmKtaCJUuJo7bodAJg+dxP
Hmtdva+IHI5Xoi9yCIwf2QohTfRthgJmqL+O200KDZKYqawr0Ep2fgM28aVY3zZH1Tg5UQ7PyqwH
tY5aqTA3NhGitRnyQwIjWVgoV4nn/hrWj/xAEdPywPA//xKZrkK74EivMig9S3qNjZZn7d2d4Irg
DrVNa7tXbU7XdmSDwYmklWCjOmPKOy9PPQUm7MapmKtPkIrG4ZkihuYVwKYBh3d7OXSvRTugHqH2
pcf4025g9ISW9yCHTYC3SsQMVQX7y8FL01iWWMgkKKpYrZB2y8pyFOmdVn4y3xo4mt6j3ZqrKLrC
yySj9Uwh6VTAx/OxO+BtIqOtP93nmiObUXIv7dsmcbQlGqaiGxzaD1fSf+CUDFCOqNXkfY5abri6
ktoHquhKbFrV8ccg5FW6OrGremAmCEy5xPmjKKJDxGvqrGIyIPqX9BJtr2tj05xFcrUkMakOww9x
IflqmWtgAJCsi9topTwDxh+cl4NGZP3+NcWpzNwYrxy07FoVWQakCmAoljBfJ/1fdGBHt48rKKXV
I8c2GuSoK9QmqICml/dQQSOrAfWEgD1vUZybiNIXllNaHAesSdccYxgNQTLIggrwybYGxDLcwJZh
eo19rn2ykJ0bzc1oMI5jRfd4hj+TwkiG+V6DVosL9U5VOLRHxnCtmd0zY6/9qgpMWl175whgzBck
H3y4v8EYlhBd2XHQ1/Drw3gIUKqrq+eE7P1ZvntzkZQK6ZOlc/egKp3E4LUzbcpq1/ov0L0Np+hN
83FwM/ItpYEtywVz0uOgrfGAWgnIghvCOkaUoMC3rRXB+vqR0ZmhHiypaAyq/wHD1cKHYkTgAUSd
9WsXuLEQ46FL//phdcfBTDImgYed4WwbGfQ48tFpgTtAH2Dd4ARkNL8eAkSjDoRuPs02RzVC5ZT4
N1ypTtwSb5RAE4nDRSUXNbszp+H20IY90eSWcIGvana7QLG4Xg5L+xOLvRydRe6CLifXLh4N/nnW
qX5Mf57tgepSti++svOytF7igEs2+IeFMMeRYi8R6eQYOAAePPTMXxgefbCSoa6g3DeJyEHTdiH3
U3pIhfhk22snXfmhmUJIl0deIZqV1VA4JwTLHRTh2ce7rzEdM1lnrtbZbvJIt/+Cli6JIkk1XLQv
us0xZPUbwPQ2ANYwbUseIuFAH3DFgvpysDxmtQciSMqr2XeJS6H83Hp6LHb1U7rDeG1/pT2hnRd8
xg3pQt44TXNNL0Rve1LqedJSDUzzvh2VoQ8z92Ig6uahXMExSbHqjdis6qUC9dLWidt3mjLOxajj
jWQqw9qBk3Ib8I+W+DVj+MmkKCY+ogj26NL289L37yi8HtS9mrMY724KppxCCWATbJCnWkbvQtbs
DLubEWzltVGo+FwOHTLGdgQbqISLYljbLBIRQzVEnbSyawFXmW/qZlVu5GN3nZD5s7rYXEKfIkLZ
ysrXvT3eOoPN6sLmqlXQrAseau3yk9GE4qkzrjmEXdrShRY+H2iaJeVcVNKl6CXe1XxbKdpqunBI
chj0jJcg5qIodwfhT2NveM0blbPrzg1/Mfh+EDx95N5W3UbvNiYM0nCH6OcBPULrv8SREO/wl/Yl
V5IlgqpxYZbSZ5hF07bvX9htxjDjsXZxkzZd5kaWw4BiKJGcB6l9of3UtZNe9yGO/dxIsG08tjiH
B/az0y8Y3iv8r9b5ABzdF4nrTnZU1nqK0q4bHEssNn+ovv0vf2ek0epCateDKEk2V4xKX9ekFHMQ
FYKGku4KqlNPhWbIiEMXtdJbrkpSc+TRJfRUrqyuaNwwUrwYBRzNzcP8fgNM7+KFIBgOTlw5z/bA
DLP98jaFUc+y554Wd4lqLxP3rxseGNTZOalaNUATAH4CnxmGv7BNNVXTQCBvxcBHyNNi0DFyyyyW
rwzqGaoOFNODYjuhDuJfjY/qVf8nO+SlHQhI2Tb0AVV62ox3I4HMVwllhmwXxlAuaBupBwbw8bpk
b0kymAOIjils3CSHZH5vltF2nuamBvsSrg08wil4H0w0eLYL6TuTX+ZjYSmdPhiOcEyUcSOcm6c/
FbYokWVrBc13L5R9Ar3uOlb2dSXPb06hg/WXph7foaGje+tTPV78kWPLkkH1jukzMAJrUWq9LQnO
Htn3z8e2K/vw6lCScgGDriY4+8Kun8Wv4Lkg4teTe9omA4BSRBgw5kWZZC4LeMe6/KG6+sZXe597
zGdrU2WfAZtWrvUfOqc4eslGnoOaXO9Jy5mwcVHNbu741c6Du3rzs3ltS30Tfwq6NP2xKYwRxCfD
Wg0BCdOG7XqwNgEKC+Cl3upIoeFitom0ZnjMWfuZa3FGIa0gOKwXA84nYZwuvt1VbHg6dsDY8m3Q
cYmcW4d1HbjoqPaPFhamwmXl9U3J0DWOB2ylhDHgfY2RWU1FXzT6ovllTVeX+/3AGRMIThMU2E0W
7fZYL/UyvKa73JOXec2R5PZgTyrKweE4XLF82qKXqui6oTkjcZOboHvQqDb5vDQiHACJBseBv+uM
Y7InXsDuiPtK9bUozsSwWqqRdNNcDf+nwYG/nF5FKVkGYixUO0yC2Zo4kc/uj8JS6CAnGnw9NTrt
jbKCIp2xUZlIkWXS3V5NBTy+ooiHS/tk0kJI5fKg3/Y/tLf68xtU+NG+hrc37b3b633x1wzp41Rm
R4xRCLFAOM2ArNI/Bh0u3uG3Y9XNtYO6n4eSy9cVRCjjWRt8jpqsLul5vBBZMx+GNVJDm5zQtgrc
sSt4g/oWIpS8IqpPjW/k0X29vmNa1kMfjnHe5+k3nwVK9u98fUYf9wDb9eqy2zIkBxp4pWO/vbd6
+pe5EQHFjcH1+oD0gjGHgJC0ek9dSBNpqk97xYaed+d6q/kAW1Yt/jsW/QSZP3uanLyS7HEW+j+n
GQkhXwOswYL52OFuT2tXFPICK//m/KUpxkG/MVAQ7+v+RXAKJfuHJq1I8rp3xJWv2PaaN7Ch7FyA
KYCxW5+y31JtjsmPomhoUcD65GWmt14M3TmmQbkRQuq/J2qEoLva7sUXcvidAbUmtHiQWmZlxbHO
ACDoX4xsr+sQ8qMhEPlvIkgs46x9mi2Vkbbq3vLOnKhAFy9LsRcCBGE5BtLgh5+31wr4opqAD3Mb
uBvJ/rgJTPS6lTCekzc5OoKJ6CvArsx3rh1mVB6iUM7pKvQDHbpJI3M07BlzGjfW5lxbcbGmQCgN
5cA31znJwjCnRDB6MaIXzUUXohHczMtsv+F3IyfMVgCgjw6T7H3BkYL3IWlhlEIoGjnGuB+gKojL
mPFmlImRa0OgIA+ZwohS3koHEc4QfkC120KPx17uaE08q1zynRSehwz/OrULd/YkYprwnf3OwEAW
Tq4D5bMUqijxJGT7v3gst4SkFyWFH2eFx3LlJeBpznGUyK+iUGmBy2hPNjN7m2rtYWQNdc7KNlI8
RBXahqKzKDOqHZdT/q/chgc8Fvx1qLU0Qc0rwwN7c30Sa24XwpGlfLzdblF7NvroRWDGGy7CN7D0
B+IXuOW6mFwBxW5IyCQZDbAjzi2qTmGuH7/4VZwEZKp9qfSztBGyHM63zKvxorUiYumyEFBWLKNA
F5eB7eAeUDm2HKJR9W78eomlVT23Y0R5eFRPiBl0HpBoAGqMQHXAeXuYQPeAk6w5PJiXpxR0cHT2
UpFPZH4OP++bojA7Rbq1tUtXqXgg7CdYAZKKfe8/QeYEm3QIvVJ0L6bdzGRZz/KLGWZ/a+puMneJ
oqjwmqiwF6bSrtLFBSNEm7JJXGtdspEcFEfYAXYyOz8PFtf+YFwCnNe+WX8D9DCTiw038+yeQ/A7
AhTR5Yo63iUdLmx7g8z4tn7n/Sa16KcEC+n1chqo7bVKaZyVeet/Yvhh/LX3cIeqHZC19BT5pdx/
cuMsBMR4O7eDDbVOhhR/P+Mtc2zET+lmKQBlyWuIdJnyTBOn/MRT5T0R4GXHtGUosa30kpb7Y2+o
l7p65k5wji/V0D1bYRqxc2xxdJkwOAagVJ03SpV/5qsMtUQwvrqctdHk2AE6oFVa0Me0iZBD3I4X
wa4soakT64LBFDvmB0J/5Ria4gkugmaYXyzNty/8wiccKaFyhZLqnDphoPJMimRlpnM+GuNLspzI
SDvo22ZEzU+Z49LT2FPOm3Dn7VSO0uNutyPAG18M1GfBQ12Hja1AZ54cXBXJieXNp15q3iA4ZxAm
qOy3dwKk7xlpJYAA1Wc5vDUQcDojPWd68ixt06l6iStDy+Q+HTvLqTxJiyZKJDbiHN9Gg/lwK62u
QzsYvBfeDjLWZFfWxJm3Q9jXwV3hslkYv8adRvtg84KeXPgK7DApFhHCVuOiCWzd0FAsPl1CzOsw
srgg9n6wnjT4CC8HCq3fFdAJzTt9r7oO/dequ+C2N7z4NYz8PIWsmkxG4vZCo401tmSCROBd8gzu
FoASxAbfUSuEaSoRlJvnchfDy6LqUNIftzwnVOAbJTrZct6XMuJLjId4OofllnC/g4KbI9wvHX/6
eEzGl8VduzG3QANOXPsveejwaJU5hrSMHmIjP4NUcWgRi9zktShADZO25b1aQgNgzWKBuDKBwsJs
X10LtRjLip5MagUk8fhWdaVZjQqKDn1+tMdmRomEsvQiUmaoYnlOYUpOo5jcD0rfRInLi1y4djQv
P3hp1u+/qYEhIrvdZRWfJSPIu6XLeGK8YOXWE9lz0Q+B19OBY8zlQRfbMwzLERsiXV2OMQL+tJKD
xDgXfB+MYtwln6RXqr/lMWDDt43Cs5U3wbT/L/A4/0Jb/MLchsWCZxVMvE7/UeedVl6mwps+lDJ2
ykgmMX445mnaEsR+YMHraM0pdFI04qTpLlLtTioRHkP4sRzNhc8rKnPG/VzfCPXbnOeLyHmVeerW
MQx6eyn5BFyPamrpKgA8B3QwBPQB8V25kchfJWeNtfPF9bJrnqsZaWTKSDObmN68n1kRNmjG7agX
VN5zF+xxi6dbCQd/W2PftTzUe9daWJsKI+2bf4M9HGXYGTNWvGEnPNk8Yi3YEDqv2iOIhvepE3dD
RIPoOjo8p0FsaOrOLw9aMLiD3QvTWKu3OKmimt4z8X0KIkXxTv732pl5x4kHNguq0e5KAr5UVKhQ
DncLoRJ+ILqIqjhxUG6TD6MhuHaRiN2I3wcEavbtqgapAyEpPrdslRvtWL4u5nP5Qe/Kr2yShVY2
Mmkg5TvpKItXgRfIYFDnwkXUic/1jYge+08HdLaTZmdYB7QtNn0mVSiWcdcby60TF89UYOd6T/7a
XrmYQZN3TpywqhUGGr0XSgXzNbOKJrzsts9JphfNdsQ46lR+Ou8f9Xdw4FfmZzSVatVxUAgf9t3g
5rrsvO1xofYfHSXvCG1FpSAxs+6G1FVjtDHrGOfLy1a95l9dcm6HlZJpEjm7/6knsWS0l1beU9pj
+uEHfkG6exub6AzwsRccrEwsl1VL3Mr14u2QcfTDiQs1TrFHMuVc7Y2t4Zb+V7+naiDN4BTDhkYS
kMLgqIqRAXjgRkFQ2DEIHfeTApoWeqSVG4ro8+kb36JoVv9NtZa5Izf8Z3UWFLO8ZytY72f801Sm
oET8LpV+ZDhQavis5VwSuMLstWSvJ7Crcd4ikTxXUZqOpMXui7EGSS0lpLLHoiBaLdBCN9N/uZ4Y
/Dc+2SHuldS8ZB+GL2PQUNc5cT9epFWD4F1V18tUDMZGlg3cSSNZ/0BsaQ+rCbwBHbVpXuXM+tio
l+EQ3UNyWYmzhdOCHua6w77xcW++qHdNMBeIn1vlKDO34J2IlV5niMI71XfmUynpeZFuxSQmxN/v
ndgB39Ul7pccePip3pvw6BIlLxjs357KfSAij07fGpTla3KnW3pvCN88hCtLoXobkGnkjvzmACZu
QknF7Ce6X+bOjtnUhVOE4ISeRBn8UTKtGU6879xy6CI5HVPNlgELZAEkeQhNY3KG66xcXcWty/cP
lCg/YgPuWcsDxjKrKZt9Wtz8PECQB2s7M55mfx6zFVU0S2uWff3k5Txabe3Y25gZ9vno/cyI4l5q
MmRI2fKDUfp1RDMbEre7YSVarirCKBlSxCAUNQWsJ7w+FDeMDYMcRnmHUBLIJyLNaGE1Ipw1gXqe
wbN4YL0opZBKFfktx7T1JctYLJRe2qj6GLWayVi4fAr5panzusNcdy3tDoqtUdXFBcR4KUd/Vd+v
2IFQ2l3Sc7l12EXmG98U6tqeMKu1vrIvCJ0Ow2j/UAcKqysiD7kfom9JP0HGs7yxF6ctHJ1i9Enb
/eEDw/Mk3GKfFLTT0j8A00NFRdzvtfcK9a6h6V+vCw1Gt9vBxK+dKFPbKMQ/kPd9BWkI+ppKDJ0E
Vz7xCvO3Z9K8AfSe6c9v691J0V4JjA+E9O2ETDwqt82+PPkkckxcD6V3U8+wpCfT0ppzJkaOQpnF
sZw9zeouv8CTEdKGta6jI/Wt8FrRbwz/BW7XL8mclIgjzKmkqzMK3Q7DZK7Z5BNtmZRlsPXPE5IQ
s9QNXQMXhPUfLc4Mz3cyPw5ZybGauG/xvzWc3vwNP006DhuT8BX67p5Xp3ie/4PZ4Qn8wdMoPTJb
jMDdBE1vs3ogTwceRMqcn2WSlK7mm4u45F4EzDJEVNzaEhJF0s32/R1vk5k3/lUwepdzcV/czOBL
BbrfSEvgRxB8Js+RW1ILHEvqD9hmW9qGValHsMhbLt36n1uOUdq5bre1IbpWY0ZUkxCTv93aha8y
kcvFJVf2u/5JHUSxpQgOeEL0VsgjYEKZ7pcSiXUcOBHZOdL1kwGawNQ8nUxv8BNrhyG/ZTZ1T+Qy
Zhz4jkLi37i2h3BotDAY1lUYT555abdSNpjcYYfWfbw8U1CQoqTBscbsbS+eDawZtE9OQD32dxYy
ss2InZiE7dq+tqJJr+6l/24ESrgdxTbcxMDBloc+wIBwSHw2BSKenT/xQccudB8YZYtGmQBWTMJb
zU+09ZZxTswXFGgGIPH5yB2bSnW9zdjPgwaWoB8RuDefkWTfyjIA12e+8ncgD1VhxvYR59/tFy6U
axMOgdgIQKes6k42uBF6U7wVn5fOzD0FZhlRYWGWRr9qxlh6pIrjtWQh99+lIVOcOCU1WmjJS7k3
lL2Ql6xsWoHFxmsPQrNtvowFlLkQXDXaWUouSw1RRmG4Zxh9lNLC/jfKw35a6fkkvwfLQrzzAEVw
HV52l0EIHBMLA5Pfskt7TkWOriI+wdmztY4UCZn/WCepUGwBLlPoH9w/nW6xX8o++X/oeZoMJUkv
hfDTl52To3eJLz83lRkcempmlhPG9MH3guqskQYF7PKY/FB+HqTUhAOb6tFc/V3NKYdiwdQ1cpor
GuraIAOqAy+5DUp/xoIIgZf1CZC7hfJ3Qic43bu+NStlppnlb7FGCs4R6Tfj608SJ8gGj1EvC0wR
ZTSvQNLh3jdX06DRSYauduHd3+v4MuarWU2NUPRWGtP61/uerPmof0prPGVuPPz6tzXzLp+esiIC
pwppdDCgz22rdIXtGu/aNeDkawcTS9t5uORd0TGYUIhkVbhQAueP9AsKhn4SAlxzsoSj4iaW0CLW
zdcTiDVnL0smE8zxs4GT0uuOrmXjEbGCBdVczM9rr7aWwKyrepm23PvJp5ukjVPA49zskMv8o8i2
ECaiHDoXXzQPLOLX1HaB8cYYmS2Ts4KQQC15cMSHgQpiSouKuJliGLFC9wyEpX/Rzvt1jeFQrYGo
Jb4fv8y/HfdgZqNM+2dl0v1vYRc2UekEiCOZw/ho6f703BzJfVQq0hdsDmzHZ/zdKJhTZGvBqino
wpzdg5gtQAMFjvQi4qu3Bf6/BpdUf7uPyFp7TKvD4WwZAi+Trb+l6RImDSLwE9rRAjcC6pFGPkb2
/TzZa6gJqig0NrsZp2avPzizNfblzp3ODlIhfJFeTMrPRoY57QvFwKtgCk5Uw4DQVMu7tu0jn4o1
dcXExHjF8a5DlNP4+wz9nOSF35B37lObfMy7aT2lIEm+BBR5x9GYizq6Hh7Rw68WznwtngQAncdw
hs6Trjjss5zBB4H3l2ZVnibcCU/FwcA2c+RfA7wNArk4spWYG173O3RS7rT+dQkgYqlNew+h/zFK
YnJMniwKZgwr1l3xwXf2p9mYlLlr7htPFW1Xz1iCPaPDGOhFkzeKr01qnOmKBsQHc55GQvlAE5rz
5IKhx78YBKsrp42FGHm9nG4KxerX/WxRYm5usBTPxeRIceu3l0UR5Bo0p7a8lGshCpX5YAm3L46u
XeJRPEQHPj89sDg1wcMTbmpmBz7nJfYw0/JcaFgVrRON94u0/Me7k4+58SKxHQ3ZpoH5qxPyTJGy
pPAWH9WrsF4Ygmb6C1fW7uCyD7wYTO0YEDwlYG9tjtA/06T53iCs2EWa9cA7bEDCrsBEkKx2RHI9
S4cK3/w4cbR2DIWLjDFFHBK9Mi+bOwF446BRa9mHRc34Za7XKOPD4IgAToZN+62ODf5Xh3i4vHpu
JFJArJpXX7hRq9Vlc/Q5k7ZqS1hZAFmjvTsS/80ib6X2bMZBHMHOjR2Yj3rR3HZIpaOHWuoncsq6
pzIFL0FaYCuEJtvnAFwLYO+EWf+w/VZASU6IZ0dHMrDKCCmNboWvHfNG3at2T04SyppGAJURei1P
oXi9oi2Y90KuIuiGoX9LE47di9iADQtDoGbKoy1n4fLLUxEpD5dk3adEIgUuKskEKBDzQMWLqfex
na+tNObv/fw/uxR3o1RCEV/Jo0PAsO+aWbMOQIBCRXFSz+tJidPvuhmg9accidjDL/JChk5vnZqh
jnq78tEkVlXv52QINdJaabr/hW6snRnMwk4phOm9NYFjcsSfMiViSXSQHAguaDUMawFzQhNJZDql
KuAoDdekDx8zK9frSFeYt/T4LENwNLwyhjAkdPgHiRcmEa1d6imf8iL9egxsD+Y0V+XM4S6Ljm9s
xda7u8PuyZ8xNml+MD+w3HsSWfr0F1oUgopqcXTQcJ8ZQbrxC5CqDmjUWSkq29A6MYQsGSwZ7Lq3
ORfquoE9rNc+kNUmQNKQwvfd+25lKyK12fs2dTY6uOvZenkAiVszIfqPQ3/PUcBe45DLE5WIUe/c
vd3BLOpPuHrYmJObSEkwLO11+XcF1FLzWZwHy3Sd4mu/Rm5rQ2l8NcZsbzvAynQlufRQeEHR45pj
RB12XZ4Rbpf/G97oJTC50GxkzoiMVYQXQHw38aTEtVWvmHBKHQmNb7BOVzaqBFZ6xD9LRV36VD4O
rSzGnIeP/5ax+ZCea0S0w/2oh4v5/vqHUcJHO3pm9fnZWcQzapZAUnczXhefCZWDlXoHJrKvzPIZ
do3mpBOuClu6+MZ5nNm3RPYHYCVlypYScFSWoRe8peEDdJ/RefoIup/HAljOM7UiJlupNJ1baaYK
drsSrXRVJ6vA5wtWOX/qYWprdh/InKnjwdpRrJhQ6AtOSRZoQxu6fg1+sLz/Vkd7d1Wjj98ynQcI
Ee7vInqQ0GlNEaUXH+3JevH/FnPBezQGsQhrEzdHxyh13EFqLvCvA1gpOwtSXE/RORg1PJnc3S5x
YgRkyrB1yNQ91BaTtn58b4YGqrSnYoRQD8nWVFN7zEFKlz89vUJK2Pdx7kxl7uU33OWz3/Cbbjmi
4WS362g9bZsBgDfSBcIxiAeOa6Puc3HE0bPI+L1GPZ71pwX++7Flxgxob68DHLX+uDzzPwcV6H3/
O5DTf/3Sgue/E8pbVnt1+AfWkA2nndQn7U7RT2jgL4mzjmYI9B7c2IPCX/iyyrPjeARRxMyiXoYp
KIMXbTUFLs/n0v8bDaErhY0GWlRSR8EI80UwZjgdpVsJXmdYQc06plrhftPcZh6uDEr0s2wzsQ0J
Fw212S2zHVE55oaepg5tMp00rsQkxZxBwbAW7QSo6+KtpeYjRnnNjHg5X2dDw0NoV7Y5g7ZLD4y4
aq9IeofjddA1lNaZFG7FJWXPtSh+8SDCSeLRRhWtIEiC8no4gU3h6Er9pC1gcLKKJ9qTuPNHKDvg
4B3x1X+gvr/o1xjgOkdHPS3vmsi1Uwjn0eYwlKZpCbzW2tPlQ67FRH5Ot16NGiGDtqCOe2m6Afhe
/v1+b8ORg+OixlFYa6U/cS9eXUqSoQIHKLvJahUrDI1/fKMf1DQZQ1lklXpFE1HD/H3d8rMPrcYU
8K8qxOU+RbIFAJdJwr76Z5CHUQZ0cNrtwpbytYCuxQcUd/1jtlXs23oYQ+DvlAZ/vRBLkss7obSd
H3OYfT6b5FxB8ct1Q1vNIN+U4wC4SfonqT6Zia4lq9hWYT/0gVzgeyMZSfek/7O/It6NCKMYPMLh
hjZn1p+7GRy/LEQWbI/9uInneDpi9RkGF7L0QvDORegJKgJXvJAopGAJSnGBkw8WWRVB70e+TmTs
7v9qmbnBPK8P4Y4XoNUi2I7jWiSwJwel6z/+FzYWJOwfX5GvGNmb3v285l0P/xUc/+AfX0gkg35Z
Tt7XDXFiuuet4Z/mrVbu+HhFulIUV/k0PX+k8NRh+VSehMBE9LGWjCDgB7Z65J3cl+IOGsBwKTft
2plmUqI6n6PZvx4sn8MjBc2ebIPejth2p6S3oDHbRM423C3tw88I8cJZXm2enT2WT+su0l/1s+IN
tY3K8FLaUsYT54OSlyhkZFXa/I46H5cvV8PixP4vHAhzyRiZqUwIFinLTxMs7l785c3lyvMnfNqN
9xSEuKlVcy4UmUlPs70JzWbpljIM8FgAi8wVuRmJrWcxl5EacBMX/zv/9RKDxPyrymhwSD3jh3KX
B3t5+i2Q8TKVvwpe7QXSbpTBacPPgmjd524xtz/i7c44WWRvDwjwto59+tOT4ARBVWcO+9ssjQf+
P1CfCpYoR6WJk3bXS+BaNUgd4lT4bNeqJeT35Gv8h4rtLx5vXf8EJnGtExkt/5E4RJs5/tS2r2ak
8V7HGyP5a249TWjZ7tzZ+oH2+QZfVpv4QJcKJXwNJIsyPwNKJawWjHl15X5fWzMT+UAluULuFvWh
Qhk6Fl7Mapyo/0uJJ9tL9q5MVsr9fBVUtHfIFjiKuvce3WGkQan+fzlZa3wLm9k+GgA/ezy92uZL
2YVHbZcqdIUgQ55DYCwHnClvHRmIs1Otfo5V3LPitl40PWBdY9wFNa/fW0wh5/XxA5AY3bfW2QS/
Z/+epYjhiH8ktDjx7TLDuAZr7oPVISVH7IkJ5qxDODLpRlyqk9Uj2v2YJhRAu+n5m9eOX+9CfhCL
uRjNGjCFB2NqFIVc7cJ6B4/y+Ec3GcwC+MvzAqYU0LKZM2XIHea7R0M/w5yL5MQYudx1dqJIg0qr
MgWUdvD/ydpB/208Burc7ABdrP4NoRy7hZtKgOL5oOQe5JU1xrexv4+DvVYA+5TP6FNFSj+fcVfW
uuVn0S+Na7q1epcGMsB9tEXoUOW00SYKp9aALgx4wHUILolPfTnzSVwOB0dpQS2G/PXZ4LVWwzLv
WoJEhjVsuqDdr2y4VVubLLnF2Ba+UlQ/sDeMNxPHLCMf51PGuGGmS7gKbnjqpc2eyyPjtr21EjwY
q62PXTJreqA0DuJT0GTqDr8bR38xAybDj71kqB6JPxZaKrYaTgGYL8NSv0BXDF/cM7mhDT97Jx74
7pgi+X2sDjmq8jY75ijWgLJE9un6Hs/NyiCtKAuWSuj3waXx1vmlo4YFx8tQkuulidMK7VZm7Lhz
JAGKFim7IBTBHSqyXuI9pPh39QAkwX3nOX7bdvK28/brqqQnX1hOlSQxRz0epXo5mMQW3uzXdW7u
iTOcItEX6KUfeCLijGOkEliCd0ZcwWkta0BpO6QI2gFLTGNYiSE/XdfoS1rBVN2Omrn9Exxo8TVo
N8cJQtinNYdNq6G6QyKR2di9+CNM8dVF5cXXVOY58qloi74KusyeZkpRaGwmHLL30gjmJKArfDvx
LHONzlXEDQxzrXrsGHffTzP8iVZFxJ2NdZ5HC8KUN8fekmWLyN9Xl2BGQpqjLvfX85pJdozm8Dbp
/JkeN0sUZ99tc38nUak2Dt0/0IHPBmMx9Ls5WN2EnEHUTspf2gxYQriufCx87NnbMwK86qouNcPH
WajsMHvZAaWLC827nBEFVUYcIcXd6HGKlIx6+yQXtC8dFp0lU1pTuEa0Pf+IJo63h0uPvlQuiXHX
zWuPJDVe/1YB3HTIV1VoogwzKrIkdTs8Z7NVIDYfP5iKcUE13sdnRATn5UlHmyubz7IACfaGzkqi
cz6KIG1yhh034ZUzvP9U6ZKyi5Cp5xz6MD2701wtac5HTAXv6RFEn0UIoX0YTt9iAxOowLnxefJT
+Aw0SVi+6xjS2Ceg4mHWYQE7h5V94pH8GRfXGp5f5ug2jsdldF7QVsJF/HoLBJwhps0wHTb8Kqey
E6lLugYWtuimKzbWavMb4R7AYLq3/LYC2rRkbO83tFvemr1z2uiED5z4DdwGuopAmvGnYRl0lt/w
2Cxyl9xSOZ6+YZGAl/kg9BwzbfvZrv5W9HN6Z2s/03B+0WwvuQPWVBctmK2INO3D7+A0jZCEGNlo
aCPxJaf4esY/DuK0BXaOwcAjG88KkLVV2k+PRIDCYwYGupVjdLGNW8fsdnLT+Q3Jc/qRGObzAopv
fUtz5HOyfaoy3CEgq1E3NivdtP+OkHg6fNcCeOhtDKjNh+NTAlS1iqPE8S2Aipdja9W4usAufZMn
z2sYBNq9M0ER4oUg659xCPeav7AhxjHtAMMMDmPWl0dIupK5sowdW6cBc3YzaJLq4dA1fnRovgl7
BUZenjTyN3A/iNDRI75QkFGx2PHIZ1n8BNd/UMc41Sgd6wjiVEJBzMGbURib2VN0TzLvDEgkmhbA
HxdOZTqULKcRDTL9F9+tuLuhC/zr7XgCBY86qgJ8r/lm5Z7+LtcUUbOccwmZHdzL6L2fSOA3KsV6
WQ92+3mTQToEXarXPrO0xpKk1/wtqB38vKDQ804NLLuYU98CT0yI+cY/MqgZmFM5eM5G37/MRqZJ
HqXwEI7k796dnh4prDksShfra651OjKfuoB9Ulmah81rijPxsND8QqshBaZ8JuMt2gI6bUrQKOvy
hdHY9dz6rs5v1H94KkrD0J+4OKaGjvmQwbs4hfB0rPsH3rxnIL8R6R6vrHcUG25ANBdOZvbcV6nz
dNSZCGkkS6mGA7AOwd2yw9Vdy/XZJxVCiueoxT73m3BoerHWZFmBgg9sNQfCmwlXQxMdDsRdX51f
o9hVDw9bG+UEBvZw7V8OY63+rpC0SKvCois8zcyY3ciOHw1t8SATZ7bQlo7m2z5IhySxyO1mmrxA
5y4R2uGvECmus5UrfwfMQ7rxObILab9Hay2YaTzF9iHf45BVHYxLIIEs0IsA81X1ftsia+QXD5Hb
STidcnaVO7lZBJ1erVz/03GVayv7g1JAMB5IAl88PSS/SY7qQfSFLzdNQgmMBZjdkOHWlR6aQFh1
kO5izyL/IsaJRTyRLPKV2cM3p10QCFs0XhBifirLUtnoX46Apq0msWjtgmiQnyi1ROXoINM1EDRx
/I6pBZSBuiLtLIwBdwcwUQILI/7dCuRoa7t7KTvCQBKsyv3Ze8VfJihb4HICeD9XU2j6iHuTDEV/
5NU4m08zE2wz03ki5BnREH+bt+012Cu/Yc05a5gcYf7dJXWv03qfH9jKTg/y5Q3+P6CHgBAb62KA
Bo/siOfbyl4fu336VQLuZMJM4sN7n/hElD1rD7bNnPVnVeZXeTnINFGvo2YpAvgjDV2zv2Q9Gi8h
+nDAXI53lJOofmvLhBRp7rAq8Hmz0NPneZhNo45haaHw8yuwhRx2wgrLhyQLeM8zx20/wt6QedT3
QHxgTbD9/54UucpRyts9kghYiZ/hlH87prqMFPb3y4ux9UJ52tRF5gCGAEKkaMQ2NH76i4koGJzx
YZIV8qCDfg2Tz75IgpnxTep4PjM8xZHLhmGL8zn/VYqjsFG2pUrclWTMuFNOr+6yRqb0aCFS3pB4
lLFSYUpiMs98bH6fhaWALdNrm3FsgULVpr6UOXXr0Z4jlT3XzpU+tZrWBjTJUcfN1SMUEhmOC8jG
JvnAU7kpAux5LbhyFvIQ4QLDU1G/AuhCGj1q96o3ERKx2oXVSoA8I49AKc+SPdbrL/li21QtEzVI
Kc9aRFp13L6BPIpavse02WjCU9q4WJnDxnIPDDDbeybteQXcr1UYU1hgbvdsG6/zlPqNiMFAkuWJ
yCuwAAaOHdNIDJr85h/pvDQIDigWK67001yYBP0AD3FunlaJFdSDWwKvkSLV8RmTXT9hb4jJ3PFJ
QZIuipVv6Rb7akp4JUgcLMLQeo4ynAJvV+8wNCusbQcG7jILJLKBYAL0dKZjzY0w9yqRcJOucIaw
TWRyPRA2P84yxxnbl2wVeYRkZklXCZV4EgvmfzzCqHyeQkkqcRwtcSLsqSAtspgpjvAQFTm+U4Lx
OeSxUUolyIs3ZyTI1NvfvBKhLWuHmXWIDC+fnzeQ4OFjOcZpNSkRZlveaLjgmCxHZaa06VzooWWE
YHy2uwK9nW4zNsl4h2VcnOMdzNW8hdRX9l758TSYoYovjKwnWxkqlqo+dVJu64sMRxudCF0KsbYR
ZWWIUThJ/KBJvpDoRUNHAOQHGVxsYmf1VfSQl313ueK/My9F43deyrXu7EcE1b0HjeTXJwRHryD9
xZ9PXti5PUKeVtLntqks50U4HvwqzhcqFwjHu9TPfhmp0sqoDoPkx6KqID4Ti6GRVEGfdJl8pnF9
kRMjHXA/qtU7nZ4aCKPUhJIZ0q3t/G6/Mx/vq0gU6pwX+UWf4BwInUqdfhztlLoJSKuqgLuhbU7i
1noIO4x3RBR2pfOGFnJZ+YZaO1xnta5R81n5VHO4AsYU09km6p8uPto5PwhRdnt7TPFWOY6BB32O
FiKSh1589RlKOL8MFX4LB7utee2DZ9C5CHR5F59bAu2LchXYDsd85sCcSWdBoY67VQ5w9KNz78m8
Hge8pN/CTU8rv/PNybsAgjw0qpYrjjgAoW9J3/iU+pg6Zw+B9H+QCxxMjuC7wl8t6SeXGnpjLpfR
FQCwYa+vXmX/LfFBLTJkl92FF3ApyjSq9W1H590iHe62Uk9mxLOxV1TuJDSqIE86KQ9O1z7MhzFq
ECxDuz5U6DODwZ5A790AcVOxLoMu8le09yipLT4bGa53XABVTOI4oL4mFWzuEGt+UOgGEimmKKdN
hfAK2bVVvXnpHbiUGpGSnfHkN3trJv6zSxGlM1Y01/a1/lhwSlRsVYpYBdg+saFtyj9GEfGpK9D6
1h6EYGwAe6bm8gLGpUZ4wm+9XV0CfH71YSmucMPwXUyQwC1gCnhXnzfC2cnR8UksfJ3fQTVizZDz
1hT21T7bRHDosXCWnxyCtvWST231WgzhzEXpfHbEN/iTD6Y91WJuhOmn+ag7MEIkoZ8szGjANp6u
wyclE8+JpAmdIA8u1f6u2pYWUp+b03riGOFxT+zTtILzwiRsSWZMHa01QzmS7moxTG78eUbglVWq
yrOvGWJfIsbbd2Q0CwVgxv0yg7Szz5iqHPZfOw+uhXst/PnisGmIJiOcOp/2I0C5fFa9vxJ4IY81
bSQrJ63fUQ2s02KKxDsodbCsjtYfTlyMd2r7RL75s3hsBiaEiZKkfSoeieEBbC6gZH4h0m39e16h
STObp4AlWhm6mz0Mysfv2BJVr+RGsTYRvt89oYfuI+I8rGQLZZIiLGaa1seCTV1C7zqRkVZ+67v9
nCLH1KoamNzU5ve5uJ5JzYRCx/065g2e7bjKBa8T1ZwCvtnYXK4CEaWMHUKqHUMYujPxtt0TKOCm
dHHPGfOOx6K7Gd4S6krykB6qNcFDCBHTMLVcFO3c7NYNLw9f+IgS8HC+cysLNdgfBEKFm40Jk0/F
8XICthXbrdYHsgwFWOTRQkxZm8pEd2vHMd8V9Zo3EmMENDs3psiCF3mTXL8GhBg0zQuL9tzYlJx/
7yiRmnWm6y/rtsP0I1pcm+Rh8BOdTDbR/Ed3JM8fkxg4EJnt+miHbMUVnlMdYY6FMEOy2+lIyaVx
UE+cBjbos9tQsEvkYmPuFl2tSIyZUdeFkvLXHyt746L7g2dEjEdF0BOGvbiMX/hjvYvUCCx7bCB2
w3bOBjyCbbEgD1ThYJCanHk0nJlNuSUZCUpxYluwQd4lRpRNs3n9PnZZ4qS2YdgJ/GW5NX1+6Ver
sEIeIeNmW2oI/z3lpEsGwIPVO9vB9CaikQ2c9mv+PMhLdBwXqVLYC1LIs16eSHgN9ib1ZWn5Xx8P
GSUV0WIxwqfGoToVkI8TuTXZSYZ5hYfLWcH/ITXMjo3Ae/BH1Sobi/nmMP4V9ljDVeIQdaT8DLda
lbflPuZZffU3Nj8tk3M10wL6Scj47kY1X3pkMbOCBHJX4QI6S2SxVAzjZPiyoQFxpl6U+Xqbnmpu
RVu3R/I6+nWIySXLUG2HEaNTcKC9CbWSuKM4+UF/DRH8YbMmiBx4HvyGkGf8l7K0nY/2RofGfpCS
rzM6i9YtKVFYj24XGpddrzPjJZb/Gkk9Jfs/R7q2lQ15bWq1HVxfZLeDhviUIZyaCqycNh3v7c3w
xalKY3BCaANppYpCqax8NUI02oOJIjc1WQkSEegF1nU0dDi+q8oPf0k8Na0ZE3NFlwLnrQPNxR43
5GwSX/XgZFle8YEu2FBi64+dqwV2nlVP2sV0SFtMti3VDE06CuoG56e3t/Ec0js0VA/ZONTE2NLS
yAxrTpqZZXDHtiMG28ann6yOd6/kK3w1d8BSxp1ClozcVoImsso+PzhWjvgkBmqK/ZlLtDOVYNCP
PEeKX/9GdYGa7tLnu2aRDRyLzblYmg8pbL+2O7B0Qys2+GC/gfxYXcr6xGUTfslhJ6wZLrM5892u
Pbq6NCSgpOOwN/iq/sAveLsaKmYWqyWxI7xQC3RZt8v+1zu/b1a/3Cud8juvu4lm5g2UfJwBF5XR
nu8pfCB3aXaSbZpMq7I3qVWn3R5l3zyRk3ySJdvf+R7+9mMHtfnKBFYvpjomvX6UjiIiLfcDD0VP
7mEScFhkCSWFCA2XMmSQfvr/qEYeSzrI0LtW8LeV/K0b6AC+rP3pzzzQs+zDFV5ecIyj5FZWYRoH
U85JYS/Ckn5jQNb6m1PrW3HGjrb5sJRp/B9PhVZe7ke1pgSXuttOraUfvmWMmEyS1HuZ9LS+hRpX
ipB8iOYmze7Ox/WukUZ4/Nq6wBnJAjYjw7xwyHgo/WkFrUfLRve+iLK6TmiuDS2/2nXrCKH6/d9e
3fU9GjxbPQb//Ov+ojaq+jiV2ZeN/fop31VAoCllTlEU7jRL9zP73cL685+OzOYIdtSSiO/7Ocm+
rnOBG1di5tTiJt0NbxTxW2y9AooYdJwaVBr7DYmF4OHFnoEHFprsPsPlGq5vkfzjGFxWI9nFnifl
JBjcQivqg5DH/PXPUQJ8ECnc4HOlJ2QNTHFeK2j5ON70muHt5A+0pT7nlesvGyE1tfKkteA8Cqnu
OpFfiiRLvZ+tdQHKPga6Be4n5R2RZ1911ZIzidFCZ3r+cdwSWTx4Dquj3Of7QB+dfJfImhFqKyhM
0R73y1GHFq1VlByKo9YAJk5gtvNOQyWBsgogw7dFYvAyevRJvsx0v7EdnAiYnr1FeMtNNqnVL+T3
rAz7+rWwseZbsps07BnF+Elr3JbaV/Ami2uf74vlLut5bgQMR/uJQatsrQxwMCAlejHCOW15Pdrl
F0iLqpOlqtHGrgHnQ2I2nP2YwdGH/gU1OiLDukfse6rTDoWA5rJtF+ouaCL71Gg2f/6SXTeNQD4W
Dt1Nf71Yv77HQz3s7al7u+dSMU7g5CxZERneAeW07hdCZteKUpJBkuNMGCFhccwWzYiar+Ip+6+M
ppLsBZBcCj9Ymc6Tg0ct662gp79AIXeYjiNF35xbq53hcWK+ad6QmEPtSUXoc6jwBktAUrvhUG0e
qzB62nPx23Db7nMtphrsrjUXersgZR+Fjo/LS/wW26svdoPwpoeLtDLnLRq3uteMQt98kdCiJkdE
bCi8i32PUtVSxwhZvQVuGuqpknCqbwdgpJGzuu//qbEW0ACuGQXxsmo0q4x35FtsqHPyXSEfNzWj
x0CZlU3lLkrKKA2D1loLwbmDWa9MY4NlddkivNnrsWuj06r3klPoF/EtWY0VlpJalT+k3XO6jR9e
VdwYMTGQtsNPnB+Z770P/RMQ1LekD6IKHXDtAmVSP6rXeyMEzGCvWMxtVYp7G2dMAzQLLgiPQEuV
UbpbQkzmrHpMcZRIdZFdj6y+uSgyc3pcCzoP1xcybJrI3VexIT9a9ZRlgmAIjxrQQi4fmJ5U46yU
7+68R+Xu+ENowWjqsQ4KUzZR7xulRtHHxVuD3Z61zHVKXmodhuM29AcwMklwStjq8XFLm45GqpVW
UqNTd2ZDvpZZVdHxm+upLyozYv4N44EmR+svP3G5xBRYeiLZEPDulO3tPoFHfwnoKkDhWgdncfga
kQaLP+PLixIjohwaLbtyqHzt+asW5aUgHASDeleJx2iOWm3SlTbxXwnlD/zEauzHLPEvMVVp5E1B
6TBf3Wmbk2zV/ZXu49E7qV7qg1ysUgJYArOBR2QgKnL5no7KKmhJ4QRdEuhqAhq/4sIzjzOzm0ta
x7DVTqyj3yGo8Q0iDs9t1MutDHqzYx2iEAwS0j09NX5TauZbxHQSjW+V3RDaWms9sFxNEe3iimQg
Ohs1Zz4xUaAvaXAhpui6Vq80+5O5Yrkj4Q+4Vy7x761cgM+WFlosJO0jJ0YdXVWqdc1GKhg+8EOX
jI/vQiE5Kzjdvr3/oNPzS+WoSqDooLks0wDsVTDtXB1NuhewAVSmPT7KoIq1N+MIWx7rHMXJ4hIV
QSvO/gciUhrAgvi+sI6Enb5WLZtr8OsZX3zpjra3QZ4G7+ggYAI4zS6C6bja1MjiuSuyPi+NT1ev
MEFvFYQvmcwR9enibdg/Du2DSWwvExsg6j9ED5t2F5i/UAvr4CmZDxlLuviIDfrXTvwZp3zqxt9L
+GzbGncbMH7s/cGGMhGPPQRjgDkxrJ8DoeXw3anzuVw3y0G6RSXpBHvMitwfS9tiWe5sbaX2zE6/
T2JUyXeuXojns2Hf+8+gX6/MKDVcYC2WcJ274LNVolgq+X6+XPPbcGccI/n7xsE29RTYbl6eEW4V
ukXz18uWA+WtBi2+//PdWIqdDTDexAdS7omhbpZUbbTbDgxTpnq3oyRHofgGY/qq1fGoZwPGqoZ/
lXn0tMENiFCnk02Y0YyUeJT1MwDAXiDCHFTrfVrglTWfoZr5Xw+jpq1oBNdAAIdXpTVvfaaPh9tR
htluSB6ExTtyTFXB5wXH8wzExP4Z3CqnA9NDaclJRf8JOiTnzE3+I+St5qb7nMJVjPB8MSyud0SS
TqqU9P2C3TInCpKNnke6iCNVNPMV3AbCWLU4PkvIQQyy+fowwchbwCqJQx3hYo9NKremc1ytH19S
jrPX1umplyYki9E2OngZS4bOqs5PiqUc5MA+W5CPo8X2Ir+E7XwSFW1mxhPMR0Wgz9+Yyy0mh2eE
nE0W2MnHqs6Jv4mF8nhvxpJIb20/2XokfTim4SjJ5kJNI/EH2oOqLPlpJAMGrARXrUKZt+56hGER
7C3y+I+/5L8lkKY3tI0c34FwqKvgdl9N2tzrE2AhrkA+7cQUgNg1W+Pd4R7Z2bHBep3ga2fydlDO
KRPRZvf286aI7s99TYDciyM1O53vTxg7/UFzxbm0zz7o7QOyvuGTx+p7raiVs5lMG17FWaf4ooyo
34fmkkBAt5VCHoaQnjDxkGKsdkhngT7nP7F0DJcn6L37d3jrPYva8y0ynJtrvPWU7h4rtRS19wMA
6Z9NuLVuBI5Mq1RNgsKsZ6E1Gc3IQ8Qom9r9RTenSeQbN2p47K4/CBgNQsrUnRLRCr32Jjx3NWxH
2ysm1aK0631D+mRQtvMeiuE41t35VAIDEgPALQckztCy6lhN9k97cOQTeKPVFPqGysxzncm0coPx
qlfKSMJ5S70KDFtQJEOePjiHlkCcmMs2ep2xoowdYSt7hFgMFTwJk0TrHQevgru3RtGdq2CupXTj
N6FVivUqsl4ZUvT5e1qn4hqTngfBdOg7rIBfn10XKSR485fsxzmSTVKX89dvpTTArJZrp09JCMMW
t9ACX4/wtR+NAH9BayNCrtMPC+6jhkYOYuZFe+oGqgvH0Tg+kj4s8OWht79JplBJuTH2azD6Gaug
19A4J+Pt595UE44lpeo5X/CLB0kXHBczgo4n2OWwVq+54la/HocdJHahBCvdXtu95OAPeQS1aNdJ
K+V262rS3LT2avTxhPf6Ow6FyaGbj/mpPt5iViNGcDD+tPGkM+wcwJBA33VgyybjUyz3SKmqD/sC
DeEBEelHtBlBHzX4MUt6oWoRX3VYqxEb7CV60EvveeAHQbLTaWR1rpMLa82Ui4XVkmQ8bJxDZ2ly
IMSiaDSMmT7W7sy/cFvdLl0Trrfg13MRZgN5pda7rX68OHlMMZupK9CO+faiKOZzVJ4++iIoYg1q
gzwtee1V6h3hfCTSu8dbszpDq83CxEaSq64LzpuSzbFqrg+Z/2nbojidJA+M67oiLf4d0WW4uj0i
LYNcCU2WySO0kkkgK49cyQ3R4SUvLfuZAvOWtzai4EwIfwdj3gGNfpuGAxoOtg10d0JDyDWg0OTv
6b5j/U1ZMLtDKAWJj14/rD6XSKZ34VulBj6/XwiyDKcBroftCLELMyLYkcHgImm/xMsVrZ7SVbaq
cbGjVFL1A0sRKlUpX6xE0nWSvjfzn6tt4lq9BPzpxz2tvknH20+mQNmoRl4IWvnlusfuT7ja7RTa
iBsYCr2cTJdXwtaAaioXgaJV2g1LkIDzkZSXfK50IjXCiAKiCJekwpKbSr9UJcXnzYv2SlBMT2yd
BKuZFJzmDzvcO6onYXQrmqc8c8C8gG65CbaKNBKZ447jJBBK8WzelaAISJsNg1uWPJKP9t4zdlfo
xzdeAmA6aLEKjtazrLosm5usq/Sq+zVYlExy6waCAC2R5/k/iuG1B3YIz8WNt6q6beDedzYQ5UKT
asdZMjd+m9LyGCKwxe6/IF6Bv8I1dttojKuV519iL+vDrRxaukBzEvxkTdTxejHVMYgBRLunIvN/
vFXbrw9B1tKLN7LRAlZ9KBnKu1Ka8evjtsSLcL4cYb0tv2N+90ZfBF21Z4G9C7vEaTZNJY0eFfbL
uVr04aJeZG7Rjd51svg8GF0AQccKVQ/VQwm5mxcfp0zVBPVq23NQEahf67xoWlgEGrqLo8KUhfMV
BVX5rgWTQAjwJm1+1Xlf1ieY2/iYeHiUvUAnNjNB37zm7pw8gcRIz3hgUgGzlLjX3dqi6n0w9ETX
6O5BIbiCVFHQbeZSqT3b8MNcHkLbCEA/E0sWdNjya9BNWlhuPZ4sZ4qwVjhu7hHuXKZAaSWGgvdu
gnHlo0n/ZxoKoUM+aIRUQV9G0p+9hdI8oGfmfQlSsP2K6+PV2a1k9asODQVFbOGTQXEhAGWae8+s
RKPj4dvjrEqCPW/lTagjUbuxdSAFCsSRUhXt7jFTaGlMkauV7mYk4LD9DiBszS0y0GksuoZkcDeW
zBkz/Fa7ASJkKYEKH+3QUu8Bj3IiiSahylj0P31/1uZREXA5Uzbtw9vBZkeaF3SHCaz5RsiQPgaW
SeMhwkKFSO8a6xkPAXrCwaRP5OXvDY6NOmaOE++2GUbHau5ulzvQOjz0QOnAEFKKIfr4CS5Ivrhe
jSdY29gpcG92XuaS9f7hicSnaIoxx9PX1qTJDQauGpvly7bWn0l0bw7afVUTiOvU90k7rJfdVdGF
66DEk/iC6mySCSKfLHign4Cg5GBOcAO2g/Qmj9NduVvFUuyGkBk9E7lIq525U4l4DgTRvZ1RsC5t
KcDHzK2YeRYGF1INjp/vZT8uVDkAUAOCBgOnz+dqe7J4MVeVOiGVyaLHT3LLUWpD1kP+D7gp20fC
MXee8DEQiTGZCQKGhwn6Gv6B19OjJssNd8nCbL0K8r1Xw7p/pKLT4SufjyFgdcRqSjb50kXsukS1
tcP6Ra0zm2NHQZEsbBEcCv/D6+Nt6Wuy/lc5KBNOXkH4bBHzRepoWTD57xtjk+Y/Zrd1ZudbFDui
EFqYeSMFFigegwogEGxYyq30vgeyWeiXZYLkOcoi/dut3/jKazPilm085TQTFprVd5/gHUU7P4l2
6hQ9cGgsH5uG7iUSM3Kj3NUo/LYiG0dhdEcznJv0+7g04h0i1zU8l4hKEQXAB1DcW4xxH1kb+vWt
8AOvQh11zjz4xJInr9J8iXGSKSiWri3JcSbsFtA/7mUfxzUrFzlFvzFG0keLztTDIVLxAPRvoCzQ
dWAfK4cfzN5orkmMra3VDcZFCNVp2hGfXyRXGJWETzm9PS1cZQXYlHJKmBKtf48MXFwx6USn96An
Uhm2lQqNaVYcjIHuIbBxYB/OFgp2sjMbHhDJjmcGOHOWzy5aS4yVvev/leIxdZd3KtPiQopDmr6v
8vndzWfwP1xNWm+WpuqoBLDyWZGQXJUIFEWtSuH5i7zicJQT3JRj3lc/EdrVqGBvb3IsuUiAw04n
9nWdRXiNbgyQsQCHQChB5pGHaqVzn3yc3lKrgjvqW0zPfoiGfbKAqtzt2thyjPawz1xBvXS7AHvW
dZ4EVyJxIATNLmP1gbmcstxS74CJi1rJdHN66b7DxWEbbdg2E1gancc5oWSbxkosX2GzatLaBNkm
vEUA2U9OAKRx7W278trVO4R0b7zd6l/5bOuRXTLc9kaQ6BuVpJpx9A/xn0C2h+Hew9M1nzZsEjuZ
+6LoGDOL3Q0PJVb2N2sWTpkYCJuNKYHxwSpEEG2iFdujw56lgVgosDZhhYgZMbdktH0gxBPBCva5
ybx5le3hu5Cqq+E9y3IeO9ai4Ua+ug/XBToMhUTlEK0RepRljWWDEaw4XIuK4ICc4PAHOJsMPIZl
z1nOQpMntxXCprkRC3KmY526jss4rZlscClehZvzErkk9bccJ7K9AL+hIf2JBUAuZWLtBRUEecKT
2Qh7aZCP5VkPa7TThrSYloOa08WbQJWJqy7K/TomIdiJsfj8F5Y20pGm943J8XMeI4KW28fXMQ1t
HoXjAQKW56Vo59URNhY8MLdFQL1CL4AwR9gQOLnX7VoKdFiMdQGpCwxYaVVH5vM944qi/VfHuNyM
qI4elOunttVx+NhuBYNV4rRYVkYxpyLepWYqJYC9BxoeFmxKjKYjr7A4sUA7Br3fIzI891UJd1Tp
GswbJYfZcnNA35wtU2qc2KXP34V1ALhrUVoXl8cyit1rZ4y6FlHt93bqGFHp9uylfHOpn4nKT1Dl
Aw8giU1sINBVHl6BlKaIFM2PalJWa4IqHsmjezLh0bBYS/75XccK9ozc3cLwhqCVmvkoRILL6JO4
RkPwHTV0a2m0SNT/fuLLzsxHWO0ybqaG8tXfWlQ7pK/TAj5jvcj6KdjcgnU7a0NfGvZVG7zDZ+FR
XkDQ3pBQ198dUU38xYl0BL5rhyWPD+Q6y0XhIzlfSQAXopIloo524/G9BX14TItr2IEEp7MwyxCb
3slQnJKELAJd2Erx9uuWvnc7aour1lqB0bUGq3d4EwQbHTjiqUrn2uDgLrdvt8JrsAl6YxPJwTuI
SJ7hscS8CL+xFfK1rOArMLsnb64m/X1NLaWQP9yIXkF/8MsyR481vX1C5F57wXfeBVRTDdbQjjH5
xLtmAaKMQ1oTxZ3yUTzMIYOPuDO1gFnmVTYryvzDQU7fHEg36E/RjD+asFpOA/rdlKGaJcFlxacq
WEfODJ7hl/iPk2IPrC4GrkxEFNOfAcHVXyM0kwlpbZmwdUpshEcjm+tKYvnI3GLudbiUCOP255pb
rZ0js5cYctRJMfn6URTGh9jP6LvC3Vk//Y0I9Cj3u7EmZZ8xa5D+9Rw+hYy2rT3aEazBvDvN3RN5
bWsmTgV9cPrM17/3gZXrkSrgkxWCpPVHBU7wwungnhhlD6ETXDntFqhGc2v+XNdm5yEJD8kVb2Wx
iPAlVVW/NUHAJGbCler80UnMSeNMfvxpjwXHV/y/IuQrcntnr8p4YjQdtRj1hU6hqK2smhhJF1f2
3AmGcE21GqmZZPuMfGEGxfXg/29HJReWRd7MQDCWww+StL5yPu4zcJzpxRK6q038uX/gXF7CKIAB
szx6eI7FRjdC7DfIaDY7FtE7bYaww8BIVlnRfjIERV7ikH1jBVE5an1AGcArBD/15I+IUc7A3+Az
PPEwibA4owkYjz+clNUPxOJbYSWb5uoOwGsrYG5OMj5seEs2vmBxIWvHIa/BHHImBXI6VK9s4d1v
+cNVuc0I02s5CaKT9rsMfEgDc9uTwjriv6nrudx0fb2ic10Sznfq9fHuLooZH4vmFVkWt0TZw/4v
vrHoIYYOoqIwD8Uer01gzJ9QndlcpiV4pR8/Lflofwx9Pg3OOuevb9ehxW+KPnnf2ZtYd8enJHb3
mFl+5/S5T/Mth1lfidLhATLwLYxvmIUAjtCsxdhFW+pawrrXDx1Z/1u8vYYcTpzO9AW5yjjC4MDU
sqC0oNepLghCcbkbHeMSxzIgretn04Eh4hOTLE3NQ1bBUy6LqFAI2j7PEz2IUlshsKm+75vmJz6g
9AhlYzVJaL8JHkPohozmLQTKrOfNsp+sqYGKSQaY/MmwBKwsMquY7kPjhhl8QhC3WDzIac8LH9LY
A8nub1aSmyNCDlmf0nwAtVyzW1MSXlIwfFcQS4AWJEZ0CvG/J+FxKuJOWQwrEmU4kAYR850CatUy
F6w8+Q/nPIpvavnDI1tgsrskqAHd7rGU9v96Bmy2EPo10eJ5hRrjCC1G8gWf4h2ADxqU0hol1Ah/
7n1nqZtSsny0RXxpTsGEO2hbnfbKQ3cwvaajA/pR0LS2QvfDwfnvGzr5dqWbYDCvj9uJ7IL/+0nS
PzKMBsg92nBQjailo+vIc3ngkl1hVELmHJ08nDi0ZbctBvKD6AtQgrrBhu56KnF4s2BZaPQ+2fDc
TspnJSZ8TtHitBkGF/jQiExuFodraHZ8gWsICbymHC+24D9kG+2qNb0h+m0vwdhPKhvtxeHd1sKx
Z4AIMGUWWnixpXALWBsmgm1GgnkFaQuSxut18smRi9DpZR9YkDjMhR6e+cuVavlpioU6jp2O8Hdq
ZYdcAxr/K4IF9N39+te77Ny86MuNAVFI/ROZW9pzeQaLs/qvZudFwSqWI6e9pHWhqHsbskoMb3Nd
/dmknV5CMtP/TdpOw3XpZ0crV0B6hRTm+uyVRXU7ligQPTb1H0oU3qokNR0bXbFORTQNDWmtHeem
QDHE4evi2UqkXbqUjl3Sl6B3A4Qn4OPyqVg2oU3Eb8xQtQ8n+FKxhsPTUYL5TU15FUzOQR/JM8T5
pvHo7uo1aBL9OivDCX6MPckHWAoVLSkhpYpeYiCByF8s8Xw9jtrx1liRox4CGCkwEYNpqgJoJEQS
S6eQbxkRwLo6BkQTw1C+R05gNqjvbBqW2Yo4mmwCQfXJXCeZQpbcGe2jqYBhRt99ej5wYgqN16qP
kMhJQuPvNQMe77z8664oN92e/m53czPnYqBS1dE6BUH5EJFa+wuBqOXl45j6Ak61Kpy4Qm66IR9G
yBXnQZlx5ROPsP4v54pRklVzVpAjzyGc/WRE/RmYRDRjQ0E1/wHnauHvAhtQZ9ZKnjFbsZXBJMIh
iNm6gF5GhvRCmgUf3yMhGza50FHvOgBid97eFyJzl4C7fivvX9hV3i644x678IjrIGKQ9ATJVPta
SOLnJ0CoUwMIY09zLTQ9cJyr9TWchWUgEpvWycWGPtRxKEaX8w0cS6RzGKI+mBybsNJzSpzgULyw
BDPrk1YKTIiLtnEvUUBFfkEaid26lWKqLaQkVKGuHthyf/srNTM3ayobxA341Iiuy+1Mb0GlB/iq
7LyMu6AQkz82WxLK584J/3hkNSORYDAM8BDeL/tNuFtzmLIrRaVDQC/zMqWZ9gnYd5VeQSx8jINl
EBPxOjIXRlwRJmuTV49H5ZRoGCvRg4lkLSomu9jYA4X4u5vdZ/cnprpso4iE3WrgwWVL6a3h5aLg
pz2vA1e21C6mzAIywE8yiCZG533PIZD/OdjCk7CrsAM50MW7OiWsbmwybPGXli/RoDFIcFMCkkrt
vgcwQx7RA7ur2grndsRELE12HPPPrmEtEKQCboZVzuNrTwOwUj2FwEq/EElo5zRGL0sa9h/OofZo
a6WifplW02zJbj+XzTBzNvrVLdGncfL829ENSCpAekF3OAbaJJRI4njWMM/lcI/UaSF2st8RzQ7u
JOn2Aq3kY6yaGeTqgWS4NcBpWYVWowA2BtCMYryFD0GbUGm2N/GqXuCYq/V1IlHjvUCY18OJ67Ju
3DYHknTEPg8266T3aSTCJUR10dsTKzjVGhI88oeYkZOTkJguhO04H3OTDfor1lBsK/C3SsAFZB2e
rHiMiI3wb7SuQ/lU1yqU92pFEeyNlUr4iTngPHbsFTSKuwFMUs0jhOh3fJLpi4QFxRjarEYX6Wx9
YdgxESkArBkuHdabB8WZzZJUUbTTGjIrH8PglCnWypUiYU6uj5Z9nCFkMhQ4WhCtkoplvglyKxd4
flT53DS7gE2jsofAxgOdgrHwRZNMIz0yoNEPJz9HNqLYW7YBwcYCzIGprP13+H7RDYqUjHCVrpoR
xk/MS9FWPfWyFst4HZjE6BtqJLEVnVBdJBClPSGKvdwq3VS0ICkAccpJVFRb878B7NsLFjYqind1
KLR6BCMXsWcobu6r4NGcPnol4et43BvsKU8xCz1JYLiRXEWLdhvK5ooWBKDcuhBqmF8ow9CbG3RL
3DVWWKKSiaYTaaJX8g6pFfHRkTJYZlH2IvRrg+WxPaAC890XeMqb0zUrl8yaT8Xz8Miv5eBrQxUJ
i0RbKsfM4IyE9R/Q4r3anMtyEeaWPdpZxpuiyLP3TZsQRBx4RTwFgSax5dIjGQCK2jIPRQ6cLkjp
oWO8Lws8n5sidkHQYM4vICsDgT/jNfd7w3ni1Ae+Y6fSz082Uc5HDqQ4+rLq0bqbxV874CDIkufR
Vd6iwtP5N/mRTUVB/c0hPbZy/rCgyIumPO4AojkmVyM//B9/ffvR/5LmKhjvdbsBUeEdNhDuj7wA
KXUpUyBn5IsyuwKPJ/KibPcJqbjsim2ifquhiGjPJvMQ3GkDJMG6pvhG82+7S1Q9aKyyG1vLGego
gnQT2oR6OiByOKqQonNUP811sSuc+FbhLdix7OZp3DrKz1a2VwdMtRTlZzzF0SiYs5r6dpi9P6cO
Q4B9mCQO3NnA6EXcwPAFrilVntd7yRVh8jboawFJFIbtv4yogYxBGTZuaRSp0TUdbhAh2fr6h9Cb
rhVJ9uMjNuS8h6HG51+1U5Ggm8b1UANCJPDDPs8vKDLc6dSEoDKnjOC/K7taUcAg+OlvW17hO8cw
61Risdc+BMJoWp8In7IbpDNpIeQAZ9ApLM2cHkFIPxD81Qv8Mt4mHMx7qcKMqlqM+rvYQPC19sWu
XCFNaOPQaKdScV7DV0wHPKjEuqR09YYCxIWeqJnxHK/zjmoxqMyisddTIDzoElz8m3uHwBwqpdsX
JfOXJV5MQ/V4poAeJUTcL2lAvUTXXBF7AAxrLtqSD0N4cU5HtDOFm8rSLrgwDrLaFTYecwcxBO8f
2YHtkbSkvTFCd4KSsFzQAOG1SjbYiYdqPXpdNFRUzBe59nV9KjlhbqeV7lTvI59mmeiq6Rp/JX3P
W2WLrBoeZFqkKPXOl9Kclo7AL2Q38awE/v4/GMMPnn5Ibagmcq+cIrBFuSFJpFdRoZl+RtLWeVIc
4h93etMxoxjxF8eWyFtc8GAqkaHbV11dZBECLpGPwdajGqD7fa34Gkvn4gVzw96glxjFsDpmyvlR
YOEWYfRzY8KgcX33olVZ8Il//uo6nR0G6Qw5DPQ47GPSmZjttI+vj1b+iQ3Txy9HcGiKP0hQgcWh
GZJwSI7ZkVSS511RtjUgUMjNUpk1n9uLEG4xfRfBEBsdOX8iLs8kzEDbJHDVpD2gK631tSyGJDn+
KjEdaojWStGb4Ep9C1jZuWygNsAew1Hq01p6cmYr3RZhZtgONyV5fJkp5A38xqwa+WspK/GP13MU
o6V1gd+rsnUj+zV7yE2wPlD1EWGkd+SuZTbt89jlOT5/G5VhEkWUbhznLwqEytU59j406kmT7MDA
E8wpk18udlYwklX9sMlPnBtfL6rorSs8f7B1mUXJo6WlHChQYd68ZnbyQpUiTIeSFK2CDiK6xBiX
CxO6zKgnyUKOtX+IGCfe9MxvI+8epty2BEKoT1ViyR9i2elAsXIenwyQyENAdyR0zRNPtxnNNR6e
+n4mFdYXhQnuMfaf0p65P1Sb/lBCdb/zIWtr5c4Dbw4VZww+06fD+y6hp+7DaJYKL7Iz4WI1x9UQ
3oPFR0dDbiVLZhPQgLjXrq/Z139bbtnCYyTmHs7V/SDZSsPIRkEhIbL63DIyZvUqEwSsDYKe8Mpg
Q7l4ksCDtFHZdYtOAoe9937OChU0aXFIH5KTKmbPq7o2Yylmmr8ihWRYssHM2vQICdeRPexgZyps
TJeJTYu4RZXuWZWFH7QIJ9+jB6/JhN95yHdUIjd/YdxsQ54BSjyPmkZOACLCCvOhzzvRzrwzP8LL
0EkVZjVwk2wk3RhL9v1mLWD4LvXbprB0A0wK7oU5h4/BXi2ZY9pYLfJ5KR6TrdOSeaNtcrQ+YF+p
N7aC8LT/ymERu+dY1erOe3bL8RMCG+ycRan8hDj5mzdLggSMopgx1xv6l3goZFtsey90Owtws3Rf
H2xFDPR90HH8KZknmpv5W2yawnplHR5dfhvdaOrZvtdwQy0d+JxLklxDumjvFZzA+jrgHz7G1brc
EIFJ5JrSZnfizrKInVPiv2tCxz5gtaXAxZUz6d0tp9NWjigkvXAph4c0eH8oJ3tFOzTTayb+OQyc
26eI6kNw9dGB7A5RAhBRXa9ex7mN/AKNtVBJ0F1ZpCdA+nNbbpYrunk5OkcDNrUlZowEbuH0XIqg
I0NmnPNEQCSQi+0V945R90dH8h8X/ApkmJnaxgB2rKgjnRmu5hgvQWNfyHHGe1PemLEWh4nRRE1p
Y7S15SCqYXRQ7WgRaeN2ig8uK7giGsDw7J9vfuBkh3mKu2otYEw6fuPCJ996YPSN+CEEGLuu8X44
l13K0XZ38N6rVHbDza8dfPiNc2FkpfZ/9IPFSDywgoUArZmfX4wyJVJ8RMmaQwc6eMPMbx37GSsI
/cZfm/Tty3edZ+pytahRVxa24Tvdp4egQwdDskYsCdHclb6qVoxy5B/ttsnjATdbuXiYa2GT5hn1
+nQZTHZGFuIWC6kc09CYPsFbMGZ2fzBI6fqP7Fm26+2dYcP+1S5wUb27NNiyVTqBJY+B/02XzoV0
co00LMHilktcAboqTsgofcppUFxCh0he16vXM0Bl+G2tF9A5vp74XY6PLGvfXVmhsrvM0rZFyDdR
CQnPh1lyDXYUZcBthV/H+b8B0/y4zSQxkNowoNQjXenP1yMvrMF6WLPm5ZQTsgzxIrFQdMNcpJfJ
qIWKQFFRAOBk+oywesY3A5UuhCR9MXgFQWUcv/Pm7jlnS8zsCzcBo7mqAHrM9OF0h9JA2ZdZf2ZB
5O0sgdrLw7Sx+YeVJ/O/7rcqHMFGgfPV0wTuSptrYTZLjROXzVOoDzX81H4bsLxaf/HzsgaKPxk9
RrVt98Fj5Avrw+4EirSvwsuKBlmL1+NoIjRECq2+gZEjJ9lttyJyynG9IRRytiDHvyiYEVG8s1t8
ZHcbrLmveX/2iQfwRGWFmb6ISbU0SeFTedHks1yDWea8M0IDWsxYsLDUyTU1XAKc/eA/Rhy7NfVF
IXbjc+0YCfwDAQKAlA3IiiLWx7ZkxpGdIS6/AX1mOggfMl7VQpSYKLJ75UUI0TcopeEOWUaIFKPx
Fvye6KmcvIga9BCPNLMvo/D0E+hv2/4ROKsPekdcASFb4yfazjohmmRFfvEqZ0QuvKegoFsZQ/Qd
VDwg7rM2w7YY98aICy8ChdwN6iRQwPKDW0md4wLsjI2+RKEOq/tH16iZ6g0/TX+2afxtC9R7GJ2Y
nr0leloC8xBF42NugJowgqJGw8PNB807olndi7BvjoI/QTZk3pw/rd3tfjCM7p57/X96ntz3mMJc
OFsE5P+Q94nL1z6nTc6SLWvJlR+f6+9/N7dQTC77A15vda3hr8caD3FEThRryNr4J7LqxD6NrqL0
qXCtZjwT8kggr2Z3uszxaQ+54icWHnKeJMfV8CQoXIstDUI5lygf5LOyZ622e/DNqATht/Px9rJA
Nzh4Xy27YFOt6bN56HTofje5R0eFgIsP7yeMJInWZroiXdvaFC98PRnRPB/BPa/PynGwDYYRDd5E
hOnTU9xJo8N5StQiLSmmxYyyQ6SQtHzdcUirL4qmAwDGQbF4W898R5jhhRQZe0SD+A1Y5Ex1XEqV
xG8m7sGTL90GSi+8CMhsi0GGnkOa1KGi4Ui2W/6I/AddVf72Wd+ihuoDX3xKz6JezxcuuJgen1E5
pXVsNhrkim2pFPtsT9NJJE1+xCJqXEyDgEDugmhECHDLPLp3cu5csK41FkdIk3TqfFwKulpouxz/
lfpnrcabz1Oo2CXhkLkUsKIvE/FlybGz2HAfqxprcPd0O4jxNgvA6f3j61AU2DEP4Xeny7BW4OuR
M3LFxZnc1Er++NUUZsoYfR5rwDpP+vRhjJULp/w+GdA5IdDwmYknfItRmfBcXGfpV1ZFslkejQLH
gWtj76hn5Gt718nkt97DeIDVBX7wqOID4JUfTyqvATQkCOh7sNhARrl0Tu7RXf3OKIp/rIibKlOe
07A2sLwwi7s18s2G2jiJrfpUNsHaklPaAJEdgjgDezSsloKaHRw8SR5Uclc4RR92yaYPFF/Z2iAR
TUV9si6QK778QnCKYSqKaJXcZGpSX7+IByq+NUrYoWmBPLX+Apr3IE54bPwCd4ktKDtPQYhc+frQ
szXtMy7EGHyRXD8+0QT9YITdQnJpb6zdM5WvlYLfRg/11Z8S/KTKGx+Hz/T4NId+bHEze8C2lQ0X
nR4xpwoPi9aeqW6uwqGZ0QB+datNK8WzuT/3xUzSUHbQGOKnt/A3xlEt0qhCsQQRzaFhS70Mx1ia
CajULElnXFYSs3541u7ez53tiyf/828bkm008QMUaoz76FXOmh+tijq8Mv/tJ7neBMaxZaU3jH36
dmQq7cQfjh36YOTsVhOj/Y3GNpAEykKUIuQPlty/X5X1RBSeU+I+T8s+9TB7InX76N8kdFE4rvOJ
4vE8dDOggQ8fpLMKhv8WwUmmqJJRkOKOMxXKKJz08yBhlAttsfN+7nplTSkDjYgPjTgLrH4pV45z
vv0dxj0XLDDXz1/TxRRKXPhhoCBPzrfwffQ4UnT7TPpko/8EBXkKZezXDfT9SYUy9EIVnI4d3VAt
SqtAhmI2k4jc8TAgbxlq97sdNRkwL21d/YXTSiIRzDJFOLCIk/kijmAPNQLsrYrwZpopPpddUwaz
LV9uvO2BFrfW8xhcnz0ux45b8xgef7HN8kRHBcpXvfjdbB6exSwGE/yN9QlJw0+vAKp1WpEUrGRP
AC6RYM+1MnJAD4G9jzI6KyWjlp1DTRLBkLi3LEQrwlYp8zIn3d5bm227zzGmAYFIoRbXpT8irzgx
05/MCT2lCU1BGFkmr7EFGBpr2uEXnirBQ3DkPwsHTcJSyTRnK3AuBliqtpLRD60AX5OqtQgK4/VD
q4Iy91nvJtn8omcCOEK1vliurExHvui5sz720ovKYODo5hqYgrpDIkDhvNCFSSKdEufFwyWg4550
UW507N77CdWMdEqanjy3RWlQf8ZsQRXT/hl++tnhuLyxVsYiOwvM6G5RmxX4bs5XdkvalMitpxTe
m6dHNUJ7PF9dbwRcgU68G/rrkDuX7K5IvUZFwu7e4nyvyaMQNGXWwuDEEY42IvbW9/M6Siyyca9p
6RpcwHmi92YgobNXwvp3LF+gsltvfnh/82pgwe774QU8dwg55JTmezYt6GEtvF6d3D31rxNWglFW
OcyNfsmfmqEUFqd4TLPlFD2m2xhGJVy5caPVgZgmVnPoHqQVMvFAsBnPWUZ65EgmAXooJNZAb4al
y88Hn/MY1tZAx41qAWGNt4WIO0AevwMkOXQTpxp9v1/1aTwNaqp2Lw6LpCqtchci3yoQhEdSZydo
7EBpoS8svJBT8u0KfjgyWRH/eWlgNmyAEauw1/sx9oPE06mGf6rQvl/mqcvanyDG6RUZwCVxA01/
E2a1frckO03kn19VWCPNohCBU3tugyIkDELBtSrEJ0b6TkimOvg2aK52kwPOrruiDcHdd63ouBuC
nwKEDzraeG/yXm+0aVEPBiV7EkxADDus39lDm+2w8yz9uKssqH9vNrsT+UA6T7V15OJGjh5ay7cZ
xURBknPbSSHcCD24dPUfEH8SXlT6PRepsn9sSKjYVHVgWX5SFiFAg2zHklX1QyaeouyUw6ftUy0X
UUZxBYHBv4S+tKYcJZAqKp7oor1qPN5rTd68i7jjuv2F0I4i/HDrxXRIJzbvL/Ah56beE8wm3J/t
Gs3FGTtzHtyGpBbZlXpTXCMtlBKvHGaufNoKK92wxgOETlNs5wd2BsgPvgl15hJCAO07PHYWNEnI
dQ+41XLJXQW6gqY0AZ5D/C+czI5rojwgjXV/hG4nnU/ckFs0D9n8bDF3yuJLLpBhGPywNhtZT+FC
mMZs8tKS7ODw8BGMcvPyKzsPUab7ZylHsiWKHUXoe7bqSOX1Qp0wPho2oO2W5LF+5BoDgNgeu0zI
CYczuIbuqD/tf22cAqFE0bXdsFxk6ScMeegrrOjaR5uh/X1EgRhPjgLG9tl83miODBVkS+NaFcyb
SwbHHVfKIjBTYsK3WloN8gD87OqdNVyVmlN2pm6OD/FxL1gWTajL2bLRwms3W0hVP88KIYKlhWbo
wiC8UMztGtdP4lmyDtHcve5M7l7txxJ+toLOqIStZrcpjNBQBBeM9HZ/PcEQ1nzTEuK3whfWEmYQ
+altnSYoKqgs4uctyTP1kVM4WChU4RhIryZ3RQuvGyJWmt61ICI1OiCPIX/OZcUmcatdu821tuAv
0N/keMkYo5yTmUwMcDxjDYijQTnfpyC+kwOCxt8jHISdTePhgTraNoZRWo3M5ijTlchJ9+lZ3vQE
N2PxvcIlsUhlA8u+E04MYydOkrstUkieONpAmxjOcoQ+7Y55p3wNKLxjZla9so69lYz1qnTY1XbK
QgGmUhprLLhpK1WXYoJWU7+OMsf4HJCB3dz/WVQcaetQZxp9T6xPqhMw3oCsrBsOtCFp166H2JA8
S5Z42fb7rzlGRdTpPoCS/0evCkkL7c5OQy2GKKBWcpFrg7WkkHTvHgLbT7OybX7uUG/hbVM6LHw7
qdbn9eenzMjQaXKutMh3/T8Z3SXrUxytUx2Uq+CFVVAYGZkT7tQa7HpVQu83PyRaxozMHXrb6LBi
ByiMfkmsW36MeLZ3xRarm9ZLeiUyWZS1nvUOhyKW6c+2Tc6cYsk1Lic0Te7vlp1T0MY2JLt55Q4e
73UU7rvyCq9xQztaXedaMuS3xPi+kPD0AZDrMfKsqUz5MsnvD9PKCo5nhBgOv39gpOZk6L0jngC4
2oZPVnD+djqNmq2FcnFW71whXH6A+J7gwKdYj4Q5mMFXr+WYbqSokT0sVO7HnuPcDXDlmWEWgT6+
wUG/4mNi57l/3hVKRV1JJukKSUgkyuJJxjLh8gI9sM1CL7rgGaMDEZTGCx1e4JxXVW5PMrtwjscJ
6QtkEl0BOQDDcbdKJMoJMTV/OhX3Nn6Ws8+kBTK9r8/i6UO8TmRK1rilB+zBr4gfdeg4aIIsxDJU
XsKJz/t1dcsFJGoeW+RcvSOvEjSgTZm+ZqlXeClVxbrP+dSMJ7f21rbCxOuINPimKthwblqseaOt
OidNGGDL4tY9FFZEc4M3QxCpEXwcrY/lNCDGUgXJs1hB4yjyPMLBeIgHvwxzEKTaOcnwjq1fTua9
UzWLEWli4LB87aUppoo9u4ZIUXXhyzlYmNQR98DiWv90QXNkCZhJHkac4zD80ldYSWW1D+W+iCea
BbSRXHSKqL7g8bIKbaGSOVSDm/pSKalB3Ui6GIHMgIO1Nu3AiSypE80tJUKf9OdIhhPcTCaXz1SV
mYNa9d6XPTmKyU3Q11i62GpuImLIZCJyj+wvppyEmczAPw52w23PV4lmmFsX3NL9DQRJLULVYbRN
QO3FVBXxD/AVGo/Q+g/zi7WEnpQFurld5QIVnAiTGvakuOwsCwXaSnRNE+drcnppReIdFWaB2QLE
0p4/dKGnBF00/mdpXa5z+JnUz4K5RTqmaarppTBReoe5GRCZ5Ei+Ln0IF6k01dVF5tYFnPAdd28z
Fk2+vbIvzSNUwvx5XBicWvB49/KFyP0iTw5R08v1PrNgw0H1ZiFr3/26TDhFw+vnECApBgfa4JXo
IV3QEnX2yEIjtSulRkoxDKL1yjIn/pb488LnV4Ku9Wcto/VMSHl1VGj5npOm0SuaEBDJ1V6+jsbH
Io18fnWPPfNpLLPT1x/1k0hgvppfjh5oCsXbiSSTqiRGqLiyXjWpAH361Emec8vyPucf6iFI2ZT5
lfkzUEfbRhlUv2B8H/UMx06/H+x5uhZD0HRRKwB1LLa/7kFb3lpLXMBaVWIgbRBMUNrCXyedkO/W
++TZfRWDnhfklkLDs+SxbaN4i/3maDAakdfHG5agbCv4YF8KM1hKYkgw/cKNTiUuBEzagewXap2t
vK51/g31JzgnaeK2i1dSs9UETIo4919gXKz/Kk8+0aVP4JymVzyg900idR63Qlb19JO9TIBDWv4r
ZvfYGvXAfiHtBOLlghIQqINdnCggPD5sZSVawsnXwR+9UZp7L9TOuC1CMxbSTagELTS3r3gkWfN9
bdj+CNhCQZwi0t76Mh9TEEcxWt/Mysl9c88O/CMUuZU/xFSGlB8rDyOJWskUqQOlKDoG0bNG6B9Q
/TQmDxw77KEknZxALKJMxaiFenAbF/vm0+JZnJ4h3oas1D3aH6iyW+sJ6sAT82ZCIjBWkiXvgZpB
OScaMd7wdvKroyOwVW3Z1FOWObv+ENRkuS9SquNB4yp2xlnIJ7H6WxG0ruk+yic4QGDSMZKx3nPC
8gA8IVbHsgzmyaIvx/DDuFm4GYNYn9X3TSWw3echXw6uwUS3OzyhYW67iwxzjKjLF12V8S4idJIR
+bSIgGosjVQZVF8wrLU8mnKcjspJnuVFJuDR9R/B4VUes9mK6x/FcF7NovkWtBTPUhpBi0UdE990
1UaHy6AzZUaGPeN3gx2hMiv/g3dBtP58yVAeEmS44wP8jnUqcMoxwVt2Pv48O0Kt5Vt34mSiLPt+
8EjC2HRSUtGxpc5nrhcQj2MqXXgJWstxIMVBow+qOfIbwij88lmbP2h/jN84eh+WufF6u6b3PxWD
TZisVBSnWCVj5Pgugjvs94CO0n4OEo31yUM72vXWGokZkMzYLn21sO/2XZyCAloT0yp1mWrdICx5
jnhouubGdC9q4VY31C5EzbYCGjbkvhUNxJgf+C2hzanf/G2X+nNPtaBPcHs9Pl7m+fwB6RcDyRot
1O203dBKdR8jVpqQXPeZ03VhqL0frVjyi6Yn5amGIeplEHYDIFw+00QrukuGYLq34oj8X+leVSte
2c57JuaK678i8UAvdP+X8o1kXEdhvQLHmPScRFveszZPtBhl4Yh9krLY+uVhGDbNT4bjw5TR2AAr
mm4jBnZwsV11s4vMbE3vOOONnM5i1+Jj7Xs9Iv0vgO2pBnUXm0QM1Scg2DgesVtXIbi79nYzhcFQ
LuK9dUxY6RY1zVrJARHHNuZ+1lW8IfnhY4ovzsgqaDVat/Cb9b5WwNj5+AxnBtr+Om8hL5Rbx5Ll
auw+fNvd8rPISXp83gagqmYkGj9FG/KwvE1qVw4tfOt49vizFTsyou/20JzJuUrQ8DxeUNe/C9Dg
Hol45fC7sRcCU1lHLo/X+dk/bIJ03C/aHvg/cbZ7eDMdH+ouPmWqvXzGgZluTWiRT7A20B7xjj35
Cq0lmGFSd0c8EFr1x3Mdo+MEKRiF/aqzvPgbVPWYrJpxGr6lCOIbe+FT2w8VqcebqoSqqCIVOc9x
GQnNPCedYXR6FAtHcXM1GPxqNtboc2o6qFr7DiejlIz7UcyvwNox2Q3F7Hwqlgys8dPyvHS2RU+L
CeYDSD+m5sE9AejqFacjuBxsjB+SfqlosQfKu/rGEPTbfB4xzkwUS/sUq76IuFgjJSsYNGXRF6vQ
xdeua/RwNSKoJeQ12QBSkbSZ/g46PdJmgsy9UEeA/3fZupOqKGJ7SObOs4doz+T+GlXhDZ7voZhW
naCqj9tq9gVGMHfxAl78nPBHek7ZadUklyZ3eZHYJ4sxm2mr5TzTwGgOS9PsLmY/GcduYZikjzlu
SkunLbgh13dqTj/Ll7gxcur70cXUerjB+A1bqjHYWtRn3dUq4cqdJ7RM75zekHE7suyJ51ezVCv8
QEA79dwTu4YcewjXR7+AiIS9EwtRtosRVc67p86aKkKFoKnI+9u/Oy9OUWd5JbVdYv5jxJYSYq9E
OGPdFAF22kS/nszVAiPiMf8xnCdjfVP3DnWZmyRRr/agMPlCr9n+FQY/7JrEG8I/uyJSMSLzLipk
nR9WQOnfZCGY6gTDO2EdHUEv5MWdYBBPjzGL0kTvHn0vzGawd/mhq3RitFuuJ/+xroA9EsbBg/Bn
J1Dksyb+sixhPdVVt5BvTnzji1hnRjaOZyMVlW7VDoPX8yow7lDUKCOQilxz4Mc4Dv5m6AIocxuP
tWm9pNgEdWxefyTbTXQOxsZXi++Ipg2Smeihb5+9BUsOc/GQ4wT/kWfk6JQSr1nxlESDAyDBTL+K
Orx2gTwyCxr2sg6FyrUXEYUeo0iNtKGTYjniAUnNclLcdnaAMFIHQDHMSGJ9BBlHQpfa8/brAfvl
vaORprylg2i9hEmd7WqWa/hXTCtocDsyv5hERNA2cJCU/MfR87d/Hkmr7g1+kB4k6vBONI5vcXt5
FoQkvQzXZKZz+F7wXIh3K4JRl6mULvOch7OJg7xWfpY7mM9o02kdU4yvVJHNfXVrzKPqFHiiDzdT
PYvmtKkrUFl3e+lXQVGgDMLsGW0PVBcEO+mwpc1cuub7rwTYCRNakhmnk5BZnFW2SpbA6fIJnGmp
T8GqbAEiJjrMmsVwpZz6dYGYN5bIX4L0iA9qwHHmNd0e3uVnsfpfQKdBtqVxQh0mRpAaiI4GqP/q
0ZFffYj/rzzhMlaEED1h8VTdF08ooFVe4EgE9Bt2pc55yhPLLVrYa66BU0h7Z9RG+3zGJjGVZzat
6VDG8QjJpaZa642pS42UYqKtUcLNY6WTFFyHvBm2L3lu0RWOD48Dt4QBtGt9TjFEnx3TokP1Gz2p
UivElEJCp6iWyhr7rmNVTq26ezTFGfjpuSvLorDLAaJeTUAqIBdcg1ExbxcwUlEuZUumq5flPmUQ
wX3pF8UFg1DMWNqZzyIM/6TlML4dibwNYev6EqzTugktoW4oz40hfPnboTbkLHIkdwbAA8IgKJlQ
QbUHGZKgwVXYCsw/XLxFB9+QSGUBvTTu+1eS5lUeBvXxZSO0QDvNZNUGRRhl/3athrV1+0LKqvQl
XTk3g5fA5t7PhvUD2suGpqaEWQMtjpgGUw1n/9JZwaOk3Uo5vmo7DTGdcuWnygBpf/3A9vqaWfOO
Yxny/HC6IKawZzyJKUVp7N2ayIUicjyAZOAOFrRg3uDDjWdVYj9Myfh+EUzQRu6aPpEC82nQBiui
4unVPe+DBrGULufR5uKi0iqOQWi5f289Wmgu46Z9s8ji8eex2FccqKVe4ydHgSdPJFq3LDFoLuMg
ApeVqsXi1+X+ydRhUMmoj1hncQir2Jm3x2rrrpbZlMB6RfHMGHr+qV/Uzp0QMpCjtCaSpW1RvR+a
BcMpP5stYFv5/GT4T1FiJUvHz9zWx5GEQWCh77416KY9q+ysd3sbKlAXpMFfSk0hBQk9mrk8aO/j
JSQvn5ATr2ellOHBOOIFf97DdP1gdamnKfrfCSbZSsrbsMhBmV6hZHK+UA5KRg+9yQjtxxhbnuct
W6wf8FsEb5cVHlxmOG4JVcowXB9df98uCHOdKMnEBdhH17yHf6cgwKb5T9ELb11vZkqPmiO8Sm9w
xYglUiHFYNyxhlj+upHPSiKX7UgRVZt6AQdd+T/rJQ+kwwqavYCtBae3/sm5bArxH3uItKxnJlQC
uXgLpe+pxYF2n5uX73VG6rDsGuSRqcWUUzRX8r15pSWO7bianfBmTuUOUeI4T/yid0bElV1ypyeB
tz3YlSu4Dj5PAXCOtRE3a/v9ELjM9vT3RQjC2p0Wxyi2Pibi04Oi8SL9LAHyfQNe5NvGgS0aItvM
LKb8/Szd2jQ3vSalwaR2rQgEc42k4lCELEvEsJZPK9uU37mjJbkBwiGcI5lwwJE3fecF6ZOzxj5R
NN2ZGeNbee7Tqa+ttsiI0vgjQIrzuqrE0JXGUIn7ra1tO3y+OuYL3RELg+UlbCq5AZ8taextP6xW
/lKa2jfT77ApJRVLHUXRggjHXTGbE/ZFeF27hzIH+rvYsIRz6NIM5xurSHqGSNTFdtm0fmCbWpU8
fPY7Vj4vTN8C4G6tFrlodS+mboIw7lYXStA+XxENYIETMxHTsk4HrA+jb17XMr6QHYtSGUoBLnj4
JgktxhH5EC69aDvyaFgLJBnHQvxmbP0JvtwtzkJMUiD9KZ6FSUvLKhFeCdghMDs0/X6rIHWsgbAh
J3ThBvkfBOvzlDGL7/Xn11aXDgfQUmwUuqmf7d9LOoTa3Lb8jECUg1q/UkSTEUKDUHsR/IxFPdOw
B0Wd+l2wRrZ5YKUWLGP9Z4HFsTi5RayiNLUK9PR0F93Gt9pdWAFJ6EBU+D3vmASrm8jAvGuU9S8J
VAV45Mbwkd9eg29238MWhafUnfGuFLPC7Wb2zI/sqKQvkyNq8Y10OI/2Xea5vtmdhD6Z/gRMkfN2
dGcn4fF2+2BhvXyh8rA1XWuxnhDAN9Lt2Fyaje044JN+oHAUExBcG1TRcF/6ACvXN/dvsCsakBq+
pkEVhhwAWQZJytgiog5ZQPBP9PbuXZPblJOFukTqitMevG8tpuWX1Ws2GoHfefvcfYh0dgJm2tVu
ZQxNkYgbyQlG8WPM3Oh6LXiYkm8VeP4zASVQDWXJrmrrzl07kFc40CYqAebdkz8N9t1o4SncY4Md
OcbG8k7htU60muikQ7QHBw6QYwqx9h3ucLaX2xs0KnG9A/m2B9H+zwX0+vUJqcGVc0voUuzK0Pf9
IzyMP2VJp28TmF7TB4lNSvCChw4P1I9eqOtsssBcQTSkYSiX8CWXHGxesv1jn6rmNbJCQEqpLRTX
fatRuLkLL3B0Zne+ZUuJsbpO04DJuC+HosV3h2OuGcwnHS+EJqdwfi8PanIyO412uvUkWephtCx1
6T+9bzs2jeBat3VuFecIfmMcHKVdQRMJGiPmpX9/UxsNyFOUNtddOCujGkWi4ld30EO9YRpCYGja
nPpFrCIs4qdtmuly6Qs6QVqtviLw1ihne7kGXcYsJkqF2ksfwfh6OJylQ/f1OvQ1cIuMaUGXLWCO
FcqI2+cAVDfwe9m7tBgDNuXeCQx6V5+kNfc20rx3hD1J8TII1PdvZQCUBA9JlpsrkXSjYhD195dc
8y6SBLopPMbor+Pd7qHekmrvbjc8onRako8ZIAPqwkeMyNMRR54Nzw5U/9zxsd6kEWxv6o+mWzNq
gw1TLShi803pN+jvncgNTBO4QVyiNxhuhlnrR/bNPaR5gxHooPfWBxTI9yFJyM8m9/38HOf8RmTT
OcSkgZoglZ0nSysdxm9fK+rQBzOXlXJXVJFetFeJjX+y7s7j3VH1XpOQiToGP1k+ZO+JNnz/JoV5
PhmTMDIdS/Zlkc0Onhom7louif+xH3RRNirdlU4DkAgqZrzxjNtXGzTswueINwd1LENjrcButOGm
nCqmsty6TPCO53n1YmS+ZTdtaAvdBubfZmR02b6rl2jfzMCNCO5j9s/xkgNbEzmFKlp2NQFc59uE
4QILAWneSsFFNCH7nrwkq3vrNb2dkhEIu6DHKyysJaWZA4ppU2S8/pn0uZJlmmG6x6tJ4uaX7YzT
ese33NlI1EowGCjrLpze0Qt8CWh5fpAxzUfV5E9JREfTZSJFjzLmhIAXujoURKvJiEsXrOC3o6D/
ax5Ojol7Be1QGhJ2vYcW4JfS+FJzUYjgr5M1sAFWtlhFE4Ihh7GJXAEggajeJWdDz87qSfnKbIBE
oMBZzA9gWtNnYYtQNuOTLr/BUBvCqN3tYUjNYZYTWgl8yqzOeU2IoqoahDtrTULEjiVOWZbKHyml
aQPULTJeJd8Jw/hrn9D0sISAVX57gajoib1mq46PpG56rpZvYNnz9Kj9devCiEF2Of5iLiPpY7Qw
ogteXwVMGI0jeDvL/fYnJCXrkZ1d4zk7OKJfRmBqHgPn2DlpQCw5ubfoy1jqAEtxyDXoqbitGIaa
sqS9vqiJNiyS90QunCUvf9INp/1iPfaKJuUeNsqUL0EWdJmB1iPnHeea/LHTWqVTvwCJ9Orh3yiS
dOQyurR1JDJ+QMwLO9T4Qh8WWEz3DrC1xLu8G/pHcRLlRq4p7xXByzBvnN17UIhhDqqEQIPYBH3L
6q0aWsgTOseXY534tCdHY5876WYbSeaHSkJqV3WMlr+3pWB2geIMWibmSyfc7lfExSaZinSlZQbP
Z7z+/xQBpsDBCBbsB8c24ey6vuEdppYU+AwGCjo8CuoGShZNChgaWf2Z/P597vdD6xLZ/B2ovEyd
T8sa9RQPmXIQYddqjdE6uTo2XPpCtHrx5hXxA7L2NfTe9Nf7lxj7ij9JC+KI1+Sl4zb4C3dH8RH0
n5E0/V7njoSXCtnX1IsPcHC4iQ9f/9vdhsu3qao/MZ/THRgh31YeICX70vpRUmV50WjoF22ZeBdz
24Acd8laqxekqFzctxKxZj7tuFyVtcNrVivbXL813v+JJ36UOhTRyXYncrQZNrhEUJYt4cJ6CJG2
cwyjrnGQfzTdphOqxnDL5ALfbS2B5no+GW2ckgGOuEbgYxEEuMluDJsoTK0QmKk8mhkOojjRXXhy
GIwdEYBn7w6iQuLcJI5TD+vKRSjyUrhTZPsBDWjlgtMK5ATJt9cfN52rWqtHzT+Wlk6oNmJmiPAI
SAtfZgMAiC5NJDixIIqJ1PzWCHsErDQMjxFXjoGAThaUzE7vVOJk11AaggfsK0d+wnbOnSfJ0GFg
N4Do5eqaR8GvnATuZlcj0xMwy602l5wWdWwmW5I0pQmTD/CiYswE4FokGPpSu98uNmSxN+Hq9IPm
yv69T3atT4OmFPDKBV5r7z5gU4l/NiVoBhqHimK8NbuK1BGWD0mVQugUML9Y2bIcxU1QLeDZLqwG
g5TgekOBuob+3H5x0XpePV0M427epm4MqLCpKS8mPWNvdWctL8LAu/QrhpVhYnvzP7qyHcOgInVM
RXeVYRX0d2oX5B3a57lNpoDZSZwiL+e5tNcYDB+GQ70GnjTO/Ms4y58yERNQ8vgdPNqtK4vzZlWj
r5hJK5+byGQiDzEUJW3vsVlvmlRM0l0u63heBqZihoEeBY4hC+sEVxUAhBGLblzsv1dLCKeRQNlk
+erWMlzAqzxnDfImrLV+Ymr5sNK+PSdVpHu5z0dRI9Ysbw7r/GlM9txouMsrirH4hq4HeVi/uJEt
hxY8x0VX3EtHS4WWmHcudBiBWx62aVXVJYmX9vNfoxUqcNmRdE/2uzvwqkx5zZsEvV8GH3MYW0ZD
q6kGT9IGalZe5ijTZSWzicj7OYUfmS7qNuRHnmY9a5BgXCdgLimm0RiKFqQNE9f7qkqy2uCAzMig
mBLhoVsWt8eDbRabXryr0SxX6gsaWEinZHVX7HsjibWOhpM6p5rj1U+kF0vCVg/4nszMQ02/mx+Y
VaTzq1kCDq3Vu5cjQord/znS4pbJeGh7fJqeL0cMIeLlJKSwx7DQEEbNaVyXxRSdCnQB76kEqQvF
9k6nerQ9XxRImkCJDXmb8xQaVbOoitcohbaVeWRkjIJ5aQceEUK8YbgWGNXxRdJkpagJozNBT+rT
hMA+mSBy1ZT7xmTyUig1y6tmr+vKNT7jFU3jhEJu1fINxCKLBrcvmolzsrJPqK2aF/2gkNUdl7N3
VMLfVYmtYqYwrCEyplsFtJwHbNNPtzT8WVc7gpLe11jrfLd11bdb7s3TOhYLeJddHD0lXH481JDc
oe5b++BzkFjzENGlCgK+mO1LxrZyAwEFU3yaRl/J1Ln5W61y5O0J0IHdm64xgADhH0xxQKFnS/Gz
PkXf+rwle0mJsI63gg5OjvRyPGUwqzOHkmxmtAgibAb1mdTSB9dmO9ZrYyUuCrnZPJJZCOVMYYn3
szLBTsgVDoWcheUom5HEkGWd4N6LlO1ba2ySeKCj2/Qxvid/sXDsoOFfJvCoS6ooq/ykWSugKPdA
hawmweZCXe3UKsT3g0Yvd6A0wIlufEES8G60kO5TyQSe4uBFWkiofE6rwj8VaFgDUb1cqC9liLVP
V51HuqNDLygpdPvuOEhTugNLIa5xuch3nFuLxfMAW2ijyVuTkn2XBmHK3AnX0o3vP34YDVFSHLg9
Uu/Cfp899SoX6w8DdmZemJAuVw6fZm4W58x6BFM0Zf1lEuk8FKdqaOieWQIMxrGznamuq9gBQNrJ
FVZE0waTUUCRgVwRpGDuYrcAKXCHGtIpho0anGcOkbbqAmOlFIx4xc76MwhzNI2iTV4pJQh/+an4
p4N184XckJRaJlIvEquIjw+dbga0vg8Jz5gIWc6KX7pnkTXQMT+Q9K90UTJPSFD/5eHTG7Zd42of
RIbn5NmY+n0x5UuxXjYEBG84gKrUJbH9EiGbHCzchxRM0e7piWPtHEEZgc0mUCTvBCgmcKn8LEow
XLc2VQV5nJNXZDo69fe3FkRmMNQ2stplQxQPj2MQSHBWsWLxofqPk1alxUVISfTKJWw5r6/XsGLx
ZPG7YsfOrgagZqXThlWf3iKA9e2fjnisNONsXIjKn6XEfB9o8l5FwfI8H6RUPTayGStY3zc2bZWB
SaBLH/OoAhF5u9Ad+ujEE1hwjnp5lh24QN+gZyA0cgBQWajAsJSnzIMJ9rIM4novmQIuLQkzfA1/
qfI8uAxr2ujt1sE8ajflRJmELfTvSyhoVgI1Rbe6QzMpR24wdPSGxaf9Zqm564tMZOp5L4ixkTj+
D6/d4eU05b2WRTu6O4Pc7e45zjaVHC6d8C+e1mU+f9x8NNDBvOJYWeIHbhRlUAvpKCApT+STggdm
pNqqwVS0SjC7QtTW5GUjgL7zCvcU1rWkw6nim79xugUg+cYQGghjX2E8AR8xBkI1czDP2zRVp/1W
UhPW9viAVeiLJ2T/SHGG/44s4p/cjZq7KpuENbBvAvZEhBrAUYiruA+kAjvx4TfZekXoyaZ8VseW
HLXIn7qwBQnV0FBdumMOgGM6HFZVWGnRB+Jv5s+xbyIlYGoSOBEDupBGsa2uyDMmPt0yOomCb8eC
2FQ12fXFKwzP45Jij2qL3pKeiJVGDmD8Bf6KJrOgNWmhs9UIIrtQ+0ebMppeDKzp3pIwDS5kG4o7
ngmj8OjQW6TgVeAKsQmRbU/d7XDRedkYFZ6KmVvxeclfTKwckaiYQelsSo7aFqmfLe5CDhAUhBrP
YOV6S2j3HwzpWK6D1Zz82L5hYJiMWtx6hrv7oBPUqm5VsnEtDRhkY2GiBZCf9Cv/DNUo9uQohVxa
e8O8wkVBN+egLHCGt1xhsCAS0Qi12EjskV1thEcfC8zuy3yWrmytemzybwu5lbqcY67dsKCBy3fJ
EdqeKVr20T0Omz3TXIjyGjePEhd9W9J3Ai/uEn0BKXtPaj0x5ahQ0Zh/v2rtivMZ/ovpo+S2NT82
yg3ZFULSnBRHo0himbC6fcARWriBYDXw8PW1KxiRKjUdo1zgXGBnATs5WrvWSTSkCErAbU3cent3
tWHZRlr9vEaxMdOE1oISrZV+NTfOY6fHhOxjv/F5sS3Fkhi3lZ86fNhoGu5mWQol+q2RzEokSBP+
5o/23DgK3y+Szf907Hi71ajB9iwzK+9IimLhiBAv09LiyYBYseRTT2iDEawDGH5FX+ZfkteHAVxV
sYrpWWQeLP83+aWi0lypEr2jxSlkL03xHFhVj7EXtJni7IA6WwxALHqmWxyWhM2O9XyrvOMFpUWL
PPauqmu3p8RHFxXC2o4NhQuNm4bY8Gy2KiFB/Rbjqpr60y04xLahNi9xgCg0u8gj+OHCO5AfLi44
wr+PavqnHsG/7cMWy6+y6efqYmReafZHFSTlzzAimaaGMD4Ghx//ppoVM+NweAX8xD8h1FHhfPEc
vy1OcxUXtQYqeytrWNjqK5X54KSb80O+hQbc8Qy+ngyCKEhZIHQXTBE/ruWuh/pqzasENA6MXJZd
Au3GCyGi0gdJFnvmwRjqXK8hUmMUJYZfatAF7alEPxCKo+zZG/Dbh8xmfnw4U7J8a9zFc2ld79DO
+qJQBQ0Fx7IGYLvtlRe3akFAy+p1bHkkstBIbpnx+ke0S9ieETo/s3kEePs5xxoxSQNVpwnIzHet
4zwZupQwW+BhFV/06SKCLVeci0FO3xIHIyLqJ/bHRaQ/5EyCnzqvCvP+Zq2tKGC7Ur81hBxxw4cP
+cvNDBD/tjaQwrXLGOykgaDGx3Ja0DbtPvj5Tja0QBxkmWQ3CHryY+swXSfEbH7n6d90I0rP4SDu
A3d95pdHrTv+OnY2dFDSj/Lv/qHegNgiJ4kcygdcsb9NgyMFDumlvJ4Tz1Tqtf0zPm6fehCm4v9c
y/4J/3ZwgJCl8f6B5DY9hghSOrP0EFfQl8njs/pytLIpxhjIqoctB2k7SehsO/Z8gnLn+7HSXLYV
6NnjSa1QSW94kLhBwAzriwJkOJofhuxW0l3zuGqdRqnMMLecPmKpIcB5MKwkcUybuR/H6xL5s3xT
I58W0/xz1YisJJrqScU4rn2x+uDRpX8aRP9L4dktUFZr02j3pgFaYMAx99aaP5EqcLDfgktkZSqd
x0QFooJtjObcJkE50GjRpu1ZJcFdwpfzuNTX3/Nmaf2xTZIDW4aEL9yu0gnc92n3GqBPqXR5EmGH
DY77crzicvqS86Z3zzK5mxSyLmoAj6ErAFk+56XQme+fWiUsHjS7cjcJ4gxLo2rjEkEQsG4k7D5A
/XYdFetWOiuH1Eo0RttwgkgU7HL2hORSroc4ro/l+UaxE4RvXFtPRsWTI7nmSYMGCcOEac1YWjHY
NbpnTpq3WzMU3PFKuvT/0R+MMI0J2Hm15EMljHp2+HSghsIhMgjtbBNyKHA9MciuxvE8dOL3unfD
Vypi4sPGmujmKIMWf905SWg0yUDB6PKEW+SZhbCd7APDhUogOrstczMdf3Mr61iiCnDOTNaUrDiI
/uiPYyM+vDgci4mfbhuCXuRvGc5y4jF/+d1qIdUyDSCFUpobPw6rRBc21tPBmwb+pcQbLqBUG5iL
1cwlNSXxSGTwe0US4ZHAAJcuK07g1jJbbAgeYk5j8FJU4U+6gqDZHi8PwC3qh3l6X/FYpjnrhKIQ
rygPwMxkor68jZrsiZ+BLfFTejFRD2jLZZ5qNX7H0JQ/efX7LLN/xMw8wdsZV16z5DO0CKwbjdhz
AZNGLZCbFcpPwg7b1thJXYu6PQ7TI99GFh9oetpNcL4W6pi7mwPXNxtGHVqOT50bspSoKMjRA9Sp
f7gpKUExGwc78dARvuSusgQhsSOUOG3+ib6OGu846ov1HzVmnUl8fHuo4IP7zh+8BDpGX7hHnxv7
uUEAFUAqYbSEP+Q6okYysuiIxk22FfwWSirBEsyCnqb9Nz9VQBVXXGkqjMSyeu8PZdg3x6J90GXm
SuPk5rvZH39S+M6LImult3ucrONe56VgtbJHpQzKE6vwpOrWnDWUv6J5Nz7PyMJV34VcHVmRS3kf
gjH0ESxELqF1ouyoNJpXEvT7sW1AF7PNcaAMZ3TePce6pyzIlkkJdo77s1zT6k+Ew8A7Pn1/gcHk
OR6lDcX6BFO0mEIV+xua/pf5IEz+n8q4y7CetkV4ai+wZ4Wwk1apEhtC2lBz0aWFnC5F7hNXzsVA
JqDHMPmJqT9nRwr1kysfAAiz38+Lia+AI/Dxstklj9N1ewUVGgJx3C304FMPhEl0dJq5e0jpFu2r
QEjNLKAdEZ5umC9MvQUY7LU4OkSsTc6N+2tdoeh7RKnRwrs85cSs3jkQju6f16XTmAyYWaAWdpcN
OD0GB4AtoIVVNJ9WPAIN6My8UD20MumIs/Cse6yNv8hRbjqmyV6X7dv0+PCegdkFT89vRR6R0lV/
r0XG6SArYL3PgZbkxXi4zA1Z6AYxLKeyvGVGSS09nR1VNT5sVtbFp8JNJAfUC8HLkQC/u+X0Epjv
HHtz9SzK+wMXWLQVCIqHaGZZePeB1Bt4upozYKEjxMBvVF6FnkyE+Zx9UYvwSKrfTzGW88fk3qvf
w2zLqNy3dYTkogU4FehGcCJtWuZ+lqafiPQgBQX9ZcIyrnPdlhLKJ1+XuO4QjdFoY/PKQYlBRaLK
aZSjK0nC16/xfBLSZ1WJeUw5h9v39GnfKksrHXEN2Ip36Q0mvL6lzEZp3FexJNXlpdQnrYE+4XT3
xpU+yaDjr5ppkPypZszfroxjXcdCvB1QaagUQLQDdEtO17n01LWHsCqhxEQYi+Xd0JPy5txSATxc
ttgbHsk3+enhS5b07qdRyp8CdxbIdRh0NYZ0OjtlW3NB1K4U5xmI+ZO2eos7rh5klzZbGMUz2Esv
cDB8qtJpvH436lZzzR3O17DxLKr1BVTvhgo12WRKtQjFZN17Gl57CZ+uSyifhJ+DTAaNBxM4FjKn
DSLTxjEkYMKECJbQsXLhToQqzTgiKp4yaAEKL0mjFB0kOcldv8oVMeQgp1CnzMjvoV47j06A/UgQ
WzQiQLnRUNBmD05QgssSc5jbXdEu9JjokgmN7o7okiFd4DfDvwGHuTPcRmw5pWZcop7lrmjZpMm1
PanxLzXNiq7EFdaiqBsP4cHWHaQk2Y1GncQ3kbWZLsumP8eZkwFhcNllLADZp6N5NK2eZ0IgJqhz
YPt49qgQZsgLSPWcuO9ywNJ+40l8o+ngsndqaoCvEC8lpAwpGwWp4qkhXoppPzlzuUfj7Me8tVgq
GO4I8x4XgqZc83dIxx70TX2fTcuA/k2q5JE0Y3/7tZBJV2IraTz6Fh+a41I9F/8Wgp2/uvHeQulS
prQg65no3KnlxGW9BJXiM0nXyuNkqVaAXk0kNRxPpfniafdSvHgMhQf5XOyrU4xE7tzLac7nm2jV
Ezc8WnCliIFDny5HAUckvUemzhfwnTxjJ8BBkxFmaLyM2jT4D2JjrRrF5IzWibiAE6W0lu+D3o79
oQrSI9eDK3ypofP2HUeAUt6qbJVUDnQNWnNIjKJM5ZlNNbSg6aVB+f2U4vHHNZw42RYeddVv4m95
zh3xIpSFipJ1x9ABVdn9NypRi1rcnQjBVWisdhtoxyb2IUuGxSHn6rL4ekPa3PY92Fhm/UImkt3Q
5LV9HuVVUC90xSCiXQnyT1YyYwlxXN35upSWwnvVK6OhQvc62iKFtUbyPjMf8XK0w1bnNyHcSvzH
K1QKyJm8BgSCKA/cPeSFz4bKsdG4C87l0vCfLG6PW5zTWty1Q9dTz5t/CmUdCZRriWjGTnj0cSeU
syqE7Kpqqf69gPP3xFzNoxa618EPuRPuOTm3Z0wfll52DJHoPF4qHP/Dr/e4M/lBUnp9BKokgnLZ
5qSia4wD7fVqiZTVYpkEkZl19CmB5AMSkyXk4alqVhU+SBThH0IvX4bCbHqW7ojoiAe72IXAlssX
NzH9N3uUat13w2QYTKZ8c/dZqfj/kv4FYAgqAz9HTofvbqyHiD65eUMvwwD5stkb/D0vs9oSg3ss
rZ1+SgbSM5SZwrF8c0KNCEPWbZ8iISnSaNjBwDubLGINvyZJ5zW4SvfsZXsIGvuu5YCK9dlOBg/0
4d+jpqi943Y2vVoM7//iFGVbB+SjFdGelYU2qDIlqm8BatM3aTHTCPMCQsBRBjL38fzwVT+9fpOl
Hc4BkGfzWRDgWiVwrZ+zjvjaxACzgLzvhy5+JjDPU3h53kTzVDED2IS6DM7CV7acWyTDe8RP1G/i
cVTHRhN+zzX9cPsnNumoXIL316AsDAIzHJgrmcaUPo06/MG1SN/A4RXAy7wjFwMyqK/DcscWG8DO
Tz3EQwMYTrDrQsms8NzUy7aMy7Z59gJGyiUoIoONAheJpMKKkxE/g2XSUo8TbbsTuya96I5y5yaY
oyfMR+lFsAR5PKa1anuabV0b7F2vY08FtBlxEBDQq/KGW27Yar4qXTiBSSEOZc1KagJ4tSa6+a4M
dkaNb7uOXK+0AWl0HAShzaQrA1UCR3PDIs/vVRJbKrshlcaBrxI+AuudE3IYClWmrYBpEPTFM7Ps
Q2LlKCPIidII2MDbV0z8CB8B/2R/e75oNR9I2LlLUZLELl/HC81PeJRUtUmZc0DpRnna9E5YhGz9
bqjmKhmLAX7/1spxJmSVFUW4o8X0ffaQUjznNZ044MHtCyTu5W6yj2vLV55dJGG2+ss4J95WeGHg
6DcDYIiPljRXyTMspd3YnCoRtkq66xeNBzYmE+hDAUc3oMukkRMaEnj8IPx9ngOuPl+xpIoNFukY
bkLBOnfuPKk7l2iojzRJmv89lq2hechKcxHsp4U3abJHRCpWAeRQvKhGXU+2TCVNwdhSahdV8CyB
DhvWwrirFpwjdU/UfhruhK495DWL/AlkpErOpJpPJ2t0KSwo9X7RxwkpV2WYYBXk1sF5Fx4tlAfa
npiwef1OrxJkfXGYw/GCUj2c7zxaDYFs56Se++zawdncbAJGXYqf3czXoMa5pLQxf81V4tX1LCLL
R1D2RkIdTD5y7qKa728jOlWjw3GG1j63dLapkDL4+v0r1dbN4DGEjB/RSGeR3kjY9YA0DI3vLANE
ZSxL39Ew8+38pJQ++4VaUnhAlKJUgRBEOKouYRUAFN9imFqti6mDTy3qUIvcXUDaPzIwvzV36Hi4
Pxsxy3M6laK+QXhjA2LTlrzNr39Z3lVIvz5JSf/upVZVt9l3OTGDfY4OnAEByRx8FzFYI8YynAIq
4powJPP6DWiHU4+9la76kAwYlkNRIwMHEBE2VBl36nVpqShvvI94NXdQ4TkXdlMWisEu8/lrrjvt
OTPfpsL5uY5y6XRortLXgQnEjXVYnhcOxEQkt6QD9ywiC1PniJl3RAw1AVCgzSMYTAcz6yNHrNIR
HEkHouX+/1sNj3ODM9eY4JzYW2AJdyphOR7qxbOa7MIOr3LAOkaPn4BPQaSUOB3h+RPEjW256QUU
Nma+0v/VzxvWRjtCBG92f2WlbIxbkDes5A2Y2wpJaCjl/aZ/s0UkmUwMuw74udPLnEv7hsJyJCQZ
n8OHfzmF6wHGYprocbgqLlL95VgrYckg2UVxXpEe7BVveXcJ3KgWRM3npENg3L8b4LmCFIGmb0y2
vS6edsR+kLVh/inN+y2mCvXkj8uTeG6GVyX1pqmIzl3LK/NeGDl8Av2gzD1utzT0Kb2fhifvX8J3
acrVChKkoNtZ5U1g7M0+6Sq5a+8H0F3Uqs7cyvKGhI5xZKD/KQpI8EBRSb2B1RBDaHCSqQJ/G/Av
41tGXnHmFsjd+oBaEyxOj7MBKDPajBEcqBii3OYPRhfRGB7EpzWpeD1wTrdrzuUy5PaghWQe9+Qu
lOGFWd0MVj1WJ5Tm1/LpZfmjbxPyq4c3GZginngSu5k1wHPHvecpY6/apb/k6Tp56AoYMSD48cKG
D3SaE5rirECwE+r+bNGicGMUPefev8cx3+4JAg2+q2Gc9xTFrWHIaDyFxrq++w6pkCvqITzTywmB
g2K3cX7ZbXHXwdPL9X0ApZdVqFJzcUo48QiRF1NIJaCgyYqnAGi06O2z0o/DP2PgnFaS9KvFUdXc
X4gq2nyNm84phdVntQsjVQ9PJM02q7//mSchWW7LSEf+FxAhWXYENYoKXixrdZerg8T8IrKQK7bm
3LFMq/JbJ4wzJAIaJf7hh07EFZOAeDKAKm5CX9aiLvkqzx+7MpcvckjCuPzPvC0v5wEcsO9LY3Ym
+dEB17XKg4y53AEXVR5nl4sOt4zleYai2ZvBpm1wTjS5rsfS6/dYy/DQciRJZgWSmQWo/4o5/yee
BoXeIYyHMjchfRtoVDQBQm6UnAlBz2L8ZIVni/uX5u58CMKeroWw1ZkoDR8VRVq/AAypPfN7KTzE
kef/4ehMZIqlTNmgwYvi+KshwWWCH6aRUvp5gQFEvKTg1jYp29OAuslPFaf8jvURq2NSw7QVi8D/
5LZ8EeUMfVpDANVOZrvQ1no1rbbW6XCUgeNjeQXziIDDyRvK73EKVwMP5yWUisw6hcgj4F8HX5Se
fgUZp+Je+4dGgvx4DcRJX8LJ6FWbFQJwIAPYMlufKvFyzzhzgKEjIIHuqwKXKz34NEcKo8tzJIl+
KhE1xqrPP4xfa6rmFZQWnplbHhLYP4m6fPqAJr/AqKD1qjmcFdsKc8h7JpSXggaUcWqCQV47kCUR
I3DS9JnpLKHHZKEz49GwLXl0R1PjXAtK3ZZNHrg+NMX01wCDfsahPVBlujLnx4ZCIrmeimUyhvxn
ygIGdTkaou6jGhJUmCzQ2/4EoVx4qXI+kbd7sa4xZDAYx/I6SOzIHIImNjQrMl2yoCMhHvjHLBz9
ozfeNFW8DF8/hlEoY1y8Da+B3K9lJtcu5zU7Rp8CXSWUeNS+THoeWLFywLIQDSNslgkg8w23e0UJ
dUrgCJioPGXmBzjfI0xA6uYFeJ+9DRcCAzPOfyO8paQulGpOms9iGAYxps8XTd5/VDMziuFAn4N2
a8KAbwTZiShQ5jtq+baxhGGztr3ndZLDCqIQuhTgA3xLQ6hcEbkois4ddG8G4YV7CYcZ9quIiCfv
Og95O//geazsOm7KtoQX4nsUTjBjlZgJrw/3y31PmzkCVTVD3Zth+rmWrxapH9xq0nV4A8WX9SW3
/uCWOKW9hPBZ7m58wzmi+HiH2aeWlaY2/Fml2sfdTVfhZ6PgZmzbLKHhGEG2sEjW0LmrZyr1FSS3
CX6IzbUplnWcHecLWgSA/XKF0hu08AUHNwepBiYsOhdoNE0mOtJLFyhqHtJiTxB68Wfu7+KK3OGw
rwmiK7khrobhUVXwsrPulQeEeo5udPawX/eyhICWTq3D00am0b7cM9GpJgmkgcoWoe3JEAak7x0T
/AuRSndVz0rRPdZ1d5nmU/71hrxNRBfdIeBJrikNAhqdM/hUzjELNfGdYjH9xNRuqbRL8TNGfyZy
IH3q5bQBumYCWFYhld4RpMpn37YKQAJEc3mBjjJgMpUupO08i2BAj/3TFXUwyC+XpJYHl3aGESW7
g+RLGDn9FweOASbG/2QMI8DqpeONt4pdtjkNXxTBRR8QA89dKITaT4n5R+QHkPSFhQO923oGTQWg
yGPnLIE2yInZwnAvsFKA8w7np9NUJBYnrjG1t1Y/rmysp6LNjBpE8UyzrnAJYI83rSDDJ/9Tsx55
wWbmAqJ+qMxBRMLDzJv5Zvoxghj7sRgY71YbZ6a5p2isA/XOlHtZjgL4ldQnIPu/Mc+/pJsWGEq4
nRnIGr1+/SLgNEk/Y7SlPD+KEG3KbBcSd1wS9Kn5oZqajJdmz3/cEI4UAqknqhfhkgutf8BMHr6y
vDqkzuPy+xaM9NQALkIduhhJHwSbjGl3qVTDJEMAJY2mUJ9yTaKavH7oxgqESusIKMjOZXyG/Rnq
xyxgALLseyFc2DC0j78xV/97q4M7EcMW94AnlecLMoVYbUS5r24RSp8ir/FTA5nXmKtJwFNS6TVb
yoL6AyKFbX4gMwII/LRcZtTXLKNV1169ci5NrKTbVqqcJjAvPuS7KiYRetWbbNFlD9n/3xxlQ+Z7
+Rt9UChuJNre3OVYu//9On8viCL8Jl8PN8j+MNhyx9h8pPXzCiWRTlP+/3VV0ZIqkzwy13Fzmy8N
wh/JRbZ7/yD0X0MwuUw683x2D2mdGIZxuKHv3U2FLfmI8+rmaUyyMbhd9VlicbhmnayTtaaAGL+9
MDS6kaqOFJuHEF80SjQLAya/JfSJc3FarLnK//6VJBFGhvOgEIqYI7Bi78VbthSKv11yYBSt4ecr
J81hgUn/nskkrM3EAVjvBkxajzIHT8RYa08oXuG3KxfqP1YZkmknwHxBH9NXyzWVzhS2upYjIDCP
RCf9PTJhwAlpHGrZ/KQ3vcryOx+KMFI0j/Ne5m3hrV/augv2B91OjK92m1uK6VAngiV8ohU5JzES
TU9kI8F07H5c81DZq3EHO2kLUKXctbTVNKEdPzjncMJE3Y58w0qfDrheriZzbnToRvoXWlV/FPxT
1IcmVnLTTRvZc83embvF3a9dOOBLfPqPsPxx9JJ+A0eCGsHYngzI1xvytaOzzA0zozYCQ1EF4Nm1
3jjnQexD6rYoteud9wPKEnShOmDDDl/qfJZrScUzyQ8Lms0+ai2HZXE66ssYJ6XGPWw7GofWywBH
iEfu4+6Rk2J3g1oZOi3YTdZSNahI6kopDtVtaxCcNt/5GOsg7ZsREKdnznChQMWbxenR1GhLvwGO
essbu+RLB716vP6DWnko+P3cWPudFeoytZ0f+UerTW+h1WFD26kU+NwI7uQiMbYo5FGyc1mK3jCZ
p2gobvKJubylnr81jMovQgurwrtwK9FHEiEHIsrGnreIYCPfjiIAoZiUbS46LMNN2gWqHduYgyer
eSN8FiLS1Ds3MciGTJSlahK0hNm/jCmAD6Ch28Fne9Zw2k8qsc0HzpwDHoW6mFhtQRDrNyogWdW0
df4PUyK+Fjxn1VH5zXED4L0ETtWcNaOi+MzE2v65D17A8ws4EF8Jcmoegjesll75Y6+YGvk+Rw+P
6wAuZX+NqTVHABQbR2twQCrX36o6MQfzoH2gW7pnN6NhN44cSJHgw7qpAax7QGeP0E/SGxH4VqCp
CLG1sVRKdiYaz1OurUz3z29l0L26H55Yw2XXJuQy8KrpRvTz/dp2kQVxcMCyJebJdad1QUXdIt0j
T/36uNbRNZsNN3paLOSCbX1BsrYa6PfIdvyDA3BI1iy4ocTvvgZeR+xx7o+vm9IbuvFvHLY0RyxJ
9MJcLiGUq6zX7Fsa7Zk0Jiz4BXN2Ly1m87hsNiCzU2H4mj5Cj+bNARJz1OJ9ZA0HPIdX1FotkS/L
TaiFCjSSZMQSrJw9/VZoV+GBd0c/mv/iTicYXWFpzBKx9WfmcnnnbcUJsmPzR3nRgGP5H0wa+PdT
goztgWPYJZOMsgX2jZhpTtrhMZMb4KI/bVa3OSNmXfqoXIQrjpO6LDCnEUfRJDKqOAL1lzU/elWe
JtYzGsMA4JLiI0Qorx+tO7a4P37FKZCg1VKnz32evGBx0OHhmoPVEvDQgzWZ+Sey6V1AURBq4LJb
UEeggCnrFrBpp4pL7nrhbLfCuDOTx7VKlX/1iCodmByu2AIpK3Ozz9VytvORCHPl5Uzn3Hwl26mC
DM6BPhSEn1n7PuyjrMSMhAwbJfFSjyIMVD3l9WK7y5j6ZpAWEI6HoqGWNBGjyjpu8voqPp6xPCz7
Aud8TW4+Vv9FJQLGF8ghGQXqLWJvqRTyAvR2ZvAg6MAm8pzcL5POUU9VfSOyhIpc+SpAK7zUn55g
ymG44LixT8M31r10+q8yBUktUuhQVIfPD9+JBgQucMU7RUJQzZ+GVWgA0L8C/xOQLapnson+WHy0
sLMJpKTDiddKP5emKFE6VXEyS9Fz1/Ny1qn1gRVdLIM8aj5L0CnFRwSyPcMRetg9sJ9mJvNsG5hD
xNsAa0Qh3h3VxBNl6enmuaajWYq6+/m+AJFPTx6g+J0qsZANkWu5R7isFmFq9ZYqKe90q09yMPJs
xMgx3W2I/cB0DXe8ejoHuZF3tDb+WsodLo4JCYTceXAeEFJxQr+JruP5hEMEbvIS4cVmf2VN8yni
5Wm1MLjRoIXI4C4IiWgYv18H5uRIAsu2wXqk223MoXDP0q3ddNH0zg/SfF+A1PHDg1FPJU716unv
deXO18qEBxM2NMRq2yFGfg7MlJS6IKKxhVutfATrtkOItigfl5NzhWDBH0wy8HHzrRcwyIc7K71u
z39BT58sXt9xwZsHxXa+qkFdIuoCIxw17n5ADEcA44BdWc3SN8ayD30+ovur5mr0rTs6/+YsoAJe
NlzArGeyiIDvnCELpC7TOeSDDjH7pv4WxnWtumgq9UYrB4Ac6RFtDfGfiDdxa6HqDjO2A+fY59qP
2B7rB8WaSsrJkOOJJIqllYqTgHQgxGDHn2nwT0ov4Vxpax/AaNH+xPRHL6cMqVW7sQqjEpUyqLCF
gDuDs6laoapuslL5Adlcpkrec9rElsv9EZ+wV/1KWi7YvL4mDYh+AIH4QPZ45AWtsdxoWAYTveSZ
iV5BUIfyYuAraCTRUUKZK30gkZXrTSOGHdWofyn93EEVYbKDzP6e8o6SdhBNrwlVVfZR5evLgj1r
RZZehiyIbIemNXY3arLd3kXVSElnPeFS15aCIAd1j/lHeJ95KmGvNw8uus6P8h6Jt34qWYu14isd
6gzdKc8pByLffyDYSksaFq2gjOvtm56rSCiWtNi8j6/N4EBuI/ap/225fYQpDFP0Gdf3a2wOXXzP
CHsG6pYAiKbvVe1geEaEvcFO71X8cT34moep+Zvvh8EB3B4MIeuNxxvCWDqYg36vCHQm/cT0xXVL
rRBSbyOV8+VtIOpcHy+h/e+X5RcvOMjd2V2Of8CBnxfi3vtEMEapGVuKMW+MVf1IWCTrsVdPO2nc
o7We0/5zbCnM1TNmy/IeI4ZJuO2T4KdMzsjsQxWaqrOjkVZbYQn53Zhe9hJRhy42oXZYDKlc6B4d
JjQ+Us4A3e9Zj4GNw7z1BaEfeCsvg/uhVHmQ3CxNZfjIbV7bKMsZrsPm2BvTWuShZ7iCL5IKCmsq
FUso1lGyzZnBVv2131u/tzDUW+sTVl5p1lKlHb+6vr6hGLUasxes5hu+S+l6XZaOqEYKGfLIzzxq
z5kCNBOSzt9f2/aWqUzhrpaNS5wBLbsB+/oRIFNQrwkeTMfxFS4580P46ElupAe2eARtgeeU6DPi
pEVN/MD5bdctdo+aBSzjOUdrFd/tFBbNayssseDQLCjwio0xQ1NVt6iv+xnLTqzV47K+9swC19xW
gLAkybNq6JZn0d29GZDxZpgpXQBaCkqouekUkILrqP6VX75zpwStJFX3TrwSvwuNuMRLHIf21vMP
EBvGsTjQ01bQPqjIgB2wvsqxzgGVCspdXGyGpguKlRzhD/n6+sfvvk+gs++3jjEdextrnyXe5tZx
aYKNbPXylNW1JZC7cnEK/XA5H8DvNPrZJndjgW/BJyLyM0j52f8c4xoPvBqkpLch80EmESUolXh2
8MxIC2He09XxiWpM31toxujsuGbli2tktQjTE1qJfO4FR3i8WrL5q5jCwv4S4RWXareSdzcDqnLT
UkARR1CyeVjFKw5xq8G3gJSCVMDMa3LGavrTR1f29Bqdtu5/uc6hZFcMFNmP1tMKqf86fHOjkFT5
a9jmwm+fy1cSPRd9vqda51avq/CERmptNUGIuT7VSomKd08RJJKRsMZgjioHaPuDMwEl1KLz9CTZ
X0I9EOX3fDIyIZjWlOd72kutTPmlA2vTyzbKI4nxwYs8O7JT5lyl2zsHwvhjn1T0/bo6Yv0b/7Nz
HgTr1pqx9PxKzj020lMr469Ix/NnD7grwitBwKzs346/FotGEicBfcPNlvWXXD4Z9hJC5BUiZZZx
lLGo/bcpA4QXq2loPh/+X1Zmxp5tp+M2AZkgWu7dkQdcmAE6UR/bufy6Zjp4zplSutlzLUxQspl4
Kmf188qxRIf9co1JF81RdwvqLhirxLxibc0RAYKNH3EJ+1n0YS/d6g7U19IBN1VMqcl7ZmUevPMF
3p0jozcxUVd98uO9xP1U+ddbF5BOtUmQsUtwuKUfY1vfzmcYHnFAev1GSZUYfWnAwJZBio3VlDxE
2r/4N87sZRdJvgE8r42SjBTYWCqFL+ITy5w0k1Wr4Ko62LqUs+0Y7cQfcMZ4FraanRMlmCIsi3UW
kl4AYVR13X4I9aqpX+3aJ/Lg7xSzCHIqtuC+eJ0ToZ09eNehAD3FzUhLykyX6Jgm8LfD1r+T2GBf
l1kEWDVYCJSeImOKHuIw7p4x8egYPIae3E59+aDwhIgKgBtbFu4AwBnIED/acsn841mEKcQqHYn+
yGfXzZ6PZy04b2W+1EYCSAQIB3YmKCSNJDMDx4FyU19Ci9uXzfD/gwjwFqByLeBhpdRn+zjLqAFE
qcGXBXSvizyPCS/pYnUYVALrTCaPh2givs9unMNidUSiF1ts8hD75xjfKIqb2OFtwH3H8K7uAXL5
F8mOshYe722LebazKMaK65uUO6NRMuPG017YgAgis0jxDBZ9DlYiF//f1whY6T34LCqmtxBRbcJE
rtq0v1h8Ah/j1Wn4i+1vjehGZ529mtrCa/upym3sG/4UpSJ2XesK4j2xNOQrbzzaTHG3nDNjdHl5
28e4Q33WZQR7ZQwx1r6HQwSBoVfTPa+Ec5XxhiiSe9i4sKH28re0tXbmemN0ZPDfXMb8Y/aOhzDI
fwWPeCV/Z4rMBm+zHtlRcH+1DWAsmzUXpxtsDcSa54dCx/gfp103S2Lsq59cpe9NMn8hbCbuhm4U
SAISf0yC8j6b8fc0b0AVlNWnof4O0/L5qNdSNwwT55S0fiEae+OJW/2rLv7PrjuDe/dxa5NZWeOy
ts/0eUZydYbuIP7POz1VmF0LK71zqbolOZIS0ZI4mZMngPEpwxhewFQxwpPPV0CBsmYw85KsYC3i
9L0W6W5AGKCzCr2kSQ==
`protect end_protected

